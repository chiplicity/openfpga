magic
tech sky130A
magscale 1 2
timestamp 1605121091
<< locali >>
rect 9229 33439 9263 33609
rect 8585 32283 8619 32521
rect 9229 25687 9263 25993
rect 8769 7259 8803 7429
rect 6469 3995 6503 4233
<< viali >>
rect 7297 36329 7331 36363
rect 7113 36193 7147 36227
rect 5365 35785 5399 35819
rect 7297 35785 7331 35819
rect 5181 35581 5215 35615
rect 7113 35581 7147 35615
rect 5825 35445 5859 35479
rect 7757 35445 7791 35479
rect 3065 35241 3099 35275
rect 4261 35241 4295 35275
rect 5365 35241 5399 35275
rect 6561 35241 6595 35275
rect 7665 35241 7699 35275
rect 2881 35105 2915 35139
rect 4077 35105 4111 35139
rect 5181 35105 5215 35139
rect 6377 35105 6411 35139
rect 7481 35105 7515 35139
rect 11325 35105 11359 35139
rect 11069 35037 11103 35071
rect 7205 34901 7239 34935
rect 8125 34901 8159 34935
rect 10057 34901 10091 34935
rect 12449 34901 12483 34935
rect 1593 34697 1627 34731
rect 3801 34697 3835 34731
rect 4261 34697 4295 34731
rect 5733 34697 5767 34731
rect 7481 34697 7515 34731
rect 13645 34697 13679 34731
rect 2697 34629 2731 34663
rect 9229 34629 9263 34663
rect 9873 34629 9907 34663
rect 11437 34629 11471 34663
rect 2421 34561 2455 34595
rect 3157 34561 3191 34595
rect 1409 34493 1443 34527
rect 2053 34493 2087 34527
rect 2513 34493 2547 34527
rect 3433 34493 3467 34527
rect 3617 34493 3651 34527
rect 5181 34493 5215 34527
rect 5549 34493 5583 34527
rect 6101 34493 6135 34527
rect 6561 34493 6595 34527
rect 7205 34493 7239 34527
rect 7849 34493 7883 34527
rect 8116 34493 8150 34527
rect 10057 34493 10091 34527
rect 10313 34493 10347 34527
rect 13461 34493 13495 34527
rect 14013 34493 14047 34527
rect 11805 34357 11839 34391
rect 1593 34153 1627 34187
rect 2697 34153 2731 34187
rect 4353 34153 4387 34187
rect 6009 34153 6043 34187
rect 7757 34153 7791 34187
rect 11161 34153 11195 34187
rect 12449 34153 12483 34187
rect 1409 34017 1443 34051
rect 2513 34017 2547 34051
rect 4169 34017 4203 34051
rect 5825 34017 5859 34051
rect 7573 34017 7607 34051
rect 9781 34017 9815 34051
rect 10048 34017 10082 34051
rect 12357 34017 12391 34051
rect 11437 33949 11471 33983
rect 12541 33949 12575 33983
rect 11989 33881 12023 33915
rect 1593 33609 1627 33643
rect 2697 33609 2731 33643
rect 7389 33609 7423 33643
rect 8125 33609 8159 33643
rect 8953 33609 8987 33643
rect 9229 33609 9263 33643
rect 9321 33609 9355 33643
rect 10609 33609 10643 33643
rect 11161 33609 11195 33643
rect 13461 33609 13495 33643
rect 8677 33473 8711 33507
rect 10149 33473 10183 33507
rect 13001 33473 13035 33507
rect 1409 33405 1443 33439
rect 2513 33405 2547 33439
rect 7205 33405 7239 33439
rect 7757 33405 7791 33439
rect 9229 33405 9263 33439
rect 9873 33405 9907 33439
rect 3157 33337 3191 33371
rect 9965 33337 9999 33371
rect 12173 33337 12207 33371
rect 12909 33337 12943 33371
rect 2053 33269 2087 33303
rect 2421 33269 2455 33303
rect 4261 33269 4295 33303
rect 5181 33269 5215 33303
rect 5917 33269 5951 33303
rect 9505 33269 9539 33303
rect 11437 33269 11471 33303
rect 11897 33269 11931 33303
rect 12449 33269 12483 33303
rect 12817 33269 12851 33303
rect 5457 33065 5491 33099
rect 10425 33065 10459 33099
rect 11897 33065 11931 33099
rect 12633 33065 12667 33099
rect 1685 32997 1719 33031
rect 1409 32929 1443 32963
rect 6920 32929 6954 32963
rect 9505 32929 9539 32963
rect 10333 32929 10367 32963
rect 5549 32861 5583 32895
rect 5733 32861 5767 32895
rect 6653 32861 6687 32895
rect 10609 32861 10643 32895
rect 11989 32861 12023 32895
rect 12081 32861 12115 32895
rect 4997 32793 5031 32827
rect 9965 32793 9999 32827
rect 2605 32725 2639 32759
rect 5089 32725 5123 32759
rect 8033 32725 8067 32759
rect 8953 32725 8987 32759
rect 11529 32725 11563 32759
rect 4997 32521 5031 32555
rect 5181 32521 5215 32555
rect 6561 32521 6595 32555
rect 8585 32521 8619 32555
rect 8677 32521 8711 32555
rect 10057 32521 10091 32555
rect 10333 32521 10367 32555
rect 10517 32521 10551 32555
rect 11621 32521 11655 32555
rect 11989 32521 12023 32555
rect 6837 32453 6871 32487
rect 5641 32385 5675 32419
rect 5733 32385 5767 32419
rect 7389 32385 7423 32419
rect 8401 32385 8435 32419
rect 4353 32317 4387 32351
rect 6193 32317 6227 32351
rect 7205 32317 7239 32351
rect 9413 32385 9447 32419
rect 11069 32385 11103 32419
rect 12449 32385 12483 32419
rect 9321 32317 9355 32351
rect 10885 32317 10919 32351
rect 7297 32249 7331 32283
rect 8585 32249 8619 32283
rect 9229 32249 9263 32283
rect 1685 32181 1719 32215
rect 4721 32181 4755 32215
rect 5549 32181 5583 32215
rect 7849 32181 7883 32215
rect 8861 32181 8895 32215
rect 10977 32181 11011 32215
rect 4813 31977 4847 32011
rect 6285 31977 6319 32011
rect 6929 31977 6963 32011
rect 8769 31977 8803 32011
rect 9505 31977 9539 32011
rect 10241 31977 10275 32011
rect 10885 31977 10919 32011
rect 11529 31977 11563 32011
rect 1685 31909 1719 31943
rect 7205 31909 7239 31943
rect 7656 31909 7690 31943
rect 10517 31909 10551 31943
rect 12081 31909 12115 31943
rect 1409 31841 1443 31875
rect 4905 31841 4939 31875
rect 5172 31841 5206 31875
rect 7389 31841 7423 31875
rect 11437 31841 11471 31875
rect 9689 31773 9723 31807
rect 11621 31773 11655 31807
rect 3709 31637 3743 31671
rect 11069 31637 11103 31671
rect 5825 31433 5859 31467
rect 6561 31433 6595 31467
rect 7205 31433 7239 31467
rect 11529 31433 11563 31467
rect 11989 31433 12023 31467
rect 7573 31297 7607 31331
rect 8217 31297 8251 31331
rect 10057 31297 10091 31331
rect 10701 31297 10735 31331
rect 1685 31229 1719 31263
rect 3709 31229 3743 31263
rect 9689 31229 9723 31263
rect 10517 31229 10551 31263
rect 10609 31229 10643 31263
rect 3617 31161 3651 31195
rect 3976 31161 4010 31195
rect 8033 31161 8067 31195
rect 8677 31161 8711 31195
rect 5089 31093 5123 31127
rect 5365 31093 5399 31127
rect 7665 31093 7699 31127
rect 8125 31093 8159 31127
rect 10149 31093 10183 31127
rect 11253 31093 11287 31127
rect 7021 30889 7055 30923
rect 8125 30889 8159 30923
rect 10241 30889 10275 30923
rect 11805 30889 11839 30923
rect 10692 30821 10726 30855
rect 3893 30753 3927 30787
rect 4445 30753 4479 30787
rect 4537 30753 4571 30787
rect 7113 30753 7147 30787
rect 10425 30753 10459 30787
rect 4629 30685 4663 30719
rect 5641 30685 5675 30719
rect 7205 30685 7239 30719
rect 2973 30549 3007 30583
rect 4077 30549 4111 30583
rect 5181 30549 5215 30583
rect 5549 30549 5583 30583
rect 6653 30549 6687 30583
rect 7757 30549 7791 30583
rect 9045 30549 9079 30583
rect 7389 30345 7423 30379
rect 11897 30345 11931 30379
rect 2237 30277 2271 30311
rect 6285 30277 6319 30311
rect 8493 30277 8527 30311
rect 9965 30277 9999 30311
rect 1593 30209 1627 30243
rect 4629 30209 4663 30243
rect 5641 30209 5675 30243
rect 6653 30209 6687 30243
rect 8033 30209 8067 30243
rect 8769 30209 8803 30243
rect 9505 30209 9539 30243
rect 11069 30209 11103 30243
rect 11529 30209 11563 30243
rect 1409 30141 1443 30175
rect 2881 30141 2915 30175
rect 9413 30141 9447 30175
rect 10885 30141 10919 30175
rect 2789 30073 2823 30107
rect 3148 30073 3182 30107
rect 5457 30073 5491 30107
rect 7757 30073 7791 30107
rect 10425 30073 10459 30107
rect 4261 30005 4295 30039
rect 4905 30005 4939 30039
rect 5089 30005 5123 30039
rect 5549 30005 5583 30039
rect 7113 30005 7147 30039
rect 7849 30005 7883 30039
rect 8953 30005 8987 30039
rect 9321 30005 9355 30039
rect 10517 30005 10551 30039
rect 10977 30005 11011 30039
rect 2789 29801 2823 29835
rect 4721 29801 4755 29835
rect 6285 29801 6319 29835
rect 6745 29801 6779 29835
rect 7757 29801 7791 29835
rect 8033 29801 8067 29835
rect 8493 29801 8527 29835
rect 10241 29801 10275 29835
rect 10425 29801 10459 29835
rect 3893 29733 3927 29767
rect 5089 29733 5123 29767
rect 8401 29733 8435 29767
rect 11152 29733 11186 29767
rect 2881 29665 2915 29699
rect 6101 29665 6135 29699
rect 6653 29665 6687 29699
rect 10609 29665 10643 29699
rect 10885 29665 10919 29699
rect 2973 29597 3007 29631
rect 5181 29597 5215 29631
rect 5365 29597 5399 29631
rect 6929 29597 6963 29631
rect 7481 29597 7515 29631
rect 8585 29597 8619 29631
rect 2421 29461 2455 29495
rect 3525 29461 3559 29495
rect 4353 29461 4387 29495
rect 5825 29461 5859 29495
rect 9229 29461 9263 29495
rect 12265 29461 12299 29495
rect 1593 29257 1627 29291
rect 2513 29257 2547 29291
rect 4813 29257 4847 29291
rect 7021 29257 7055 29291
rect 8125 29257 8159 29291
rect 10977 29257 11011 29291
rect 11253 29257 11287 29291
rect 3433 29189 3467 29223
rect 5181 29189 5215 29223
rect 9137 29189 9171 29223
rect 2053 29121 2087 29155
rect 4077 29121 4111 29155
rect 5641 29121 5675 29155
rect 5825 29121 5859 29155
rect 9689 29121 9723 29155
rect 1409 29053 1443 29087
rect 5549 29053 5583 29087
rect 8493 29053 8527 29087
rect 10149 29053 10183 29087
rect 3341 28985 3375 29019
rect 3801 28985 3835 29019
rect 6285 28985 6319 29019
rect 8953 28985 8987 29019
rect 9597 28985 9631 29019
rect 10517 28985 10551 29019
rect 2881 28917 2915 28951
rect 3893 28917 3927 28951
rect 7297 28917 7331 28951
rect 8309 28917 8343 28951
rect 9505 28917 9539 28951
rect 2513 28713 2547 28747
rect 4077 28713 4111 28747
rect 4445 28713 4479 28747
rect 5181 28713 5215 28747
rect 6377 28713 6411 28747
rect 7021 28713 7055 28747
rect 8217 28713 8251 28747
rect 8585 28713 8619 28747
rect 9965 28713 9999 28747
rect 3525 28645 3559 28679
rect 7481 28645 7515 28679
rect 4537 28577 4571 28611
rect 5549 28577 5583 28611
rect 5917 28577 5951 28611
rect 7573 28577 7607 28611
rect 10701 28577 10735 28611
rect 4629 28509 4663 28543
rect 7665 28509 7699 28543
rect 9137 28509 9171 28543
rect 10793 28509 10827 28543
rect 10977 28509 11011 28543
rect 7113 28441 7147 28475
rect 3893 28373 3927 28407
rect 5733 28373 5767 28407
rect 10333 28373 10367 28407
rect 2053 28169 2087 28203
rect 3433 28169 3467 28203
rect 4629 28169 4663 28203
rect 6653 28169 6687 28203
rect 8033 28169 8067 28203
rect 10425 28169 10459 28203
rect 10793 28169 10827 28203
rect 11069 28169 11103 28203
rect 11529 28169 11563 28203
rect 1593 28101 1627 28135
rect 7021 28101 7055 28135
rect 4261 28033 4295 28067
rect 5641 28033 5675 28067
rect 5825 28033 5859 28067
rect 7481 28033 7515 28067
rect 7665 28033 7699 28067
rect 8493 28033 8527 28067
rect 1409 27965 1443 27999
rect 3985 27965 4019 27999
rect 5549 27965 5583 27999
rect 7389 27965 7423 27999
rect 8953 27965 8987 27999
rect 9045 27965 9079 27999
rect 3157 27897 3191 27931
rect 4077 27897 4111 27931
rect 5089 27897 5123 27931
rect 6285 27897 6319 27931
rect 9312 27897 9346 27931
rect 3617 27829 3651 27863
rect 5181 27829 5215 27863
rect 8769 27829 8803 27863
rect 3709 27625 3743 27659
rect 4353 27625 4387 27659
rect 7113 27625 7147 27659
rect 8769 27625 8803 27659
rect 9137 27625 9171 27659
rect 10977 27625 11011 27659
rect 4629 27557 4663 27591
rect 5089 27557 5123 27591
rect 11774 27557 11808 27591
rect 5181 27489 5215 27523
rect 5448 27489 5482 27523
rect 7645 27489 7679 27523
rect 10333 27489 10367 27523
rect 7389 27421 7423 27455
rect 10425 27421 10459 27455
rect 10609 27421 10643 27455
rect 11529 27421 11563 27455
rect 6561 27285 6595 27319
rect 9413 27285 9447 27319
rect 9965 27285 9999 27319
rect 12909 27285 12943 27319
rect 3433 27081 3467 27115
rect 5641 27081 5675 27115
rect 6469 27081 6503 27115
rect 9321 27081 9355 27115
rect 11529 27081 11563 27115
rect 6009 27013 6043 27047
rect 3801 26945 3835 26979
rect 4261 26945 4295 26979
rect 10885 26945 10919 26979
rect 10977 26945 11011 26979
rect 6377 26877 6411 26911
rect 6653 26877 6687 26911
rect 7481 26877 7515 26911
rect 4169 26809 4203 26843
rect 4528 26809 4562 26843
rect 7726 26809 7760 26843
rect 10793 26809 10827 26843
rect 7297 26741 7331 26775
rect 8861 26741 8895 26775
rect 9689 26741 9723 26775
rect 10057 26741 10091 26775
rect 10425 26741 10459 26775
rect 11897 26741 11931 26775
rect 4077 26537 4111 26571
rect 5549 26537 5583 26571
rect 10149 26537 10183 26571
rect 11069 26537 11103 26571
rect 1685 26469 1719 26503
rect 4445 26469 4479 26503
rect 6184 26469 6218 26503
rect 10793 26469 10827 26503
rect 1409 26401 1443 26435
rect 7941 26401 7975 26435
rect 10057 26401 10091 26435
rect 4537 26333 4571 26367
rect 4721 26333 4755 26367
rect 5273 26333 5307 26367
rect 5917 26333 5951 26367
rect 10333 26333 10367 26367
rect 7297 26265 7331 26299
rect 9689 26265 9723 26299
rect 7573 26197 7607 26231
rect 4169 25993 4203 26027
rect 6285 25993 6319 26027
rect 6653 25993 6687 26027
rect 7481 25993 7515 26027
rect 9229 25993 9263 26027
rect 11253 25993 11287 26027
rect 2237 25925 2271 25959
rect 5181 25925 5215 25959
rect 9045 25925 9079 25959
rect 1593 25857 1627 25891
rect 5733 25857 5767 25891
rect 1409 25789 1443 25823
rect 5641 25789 5675 25823
rect 4537 25721 4571 25755
rect 5549 25721 5583 25755
rect 10793 25857 10827 25891
rect 10057 25789 10091 25823
rect 11529 25789 11563 25823
rect 2513 25653 2547 25687
rect 4905 25653 4939 25687
rect 9229 25653 9263 25687
rect 9321 25653 9355 25687
rect 9689 25653 9723 25687
rect 9873 25653 9907 25687
rect 10149 25653 10183 25687
rect 10517 25653 10551 25687
rect 10609 25653 10643 25687
rect 5457 25449 5491 25483
rect 5733 25449 5767 25483
rect 9505 25449 9539 25483
rect 12633 25449 12667 25483
rect 13185 25449 13219 25483
rect 10149 25381 10183 25415
rect 1409 25313 1443 25347
rect 4333 25313 4367 25347
rect 6469 25313 6503 25347
rect 10977 25313 11011 25347
rect 11621 25313 11655 25347
rect 12541 25313 12575 25347
rect 1593 25245 1627 25279
rect 4077 25245 4111 25279
rect 11069 25245 11103 25279
rect 11161 25245 11195 25279
rect 12817 25245 12851 25279
rect 10609 25177 10643 25211
rect 6193 25109 6227 25143
rect 6285 25109 6319 25143
rect 7205 25109 7239 25143
rect 7481 25109 7515 25143
rect 9137 25109 9171 25143
rect 12173 25109 12207 25143
rect 1593 24905 1627 24939
rect 6285 24905 6319 24939
rect 10609 24905 10643 24939
rect 13461 24905 13495 24939
rect 4629 24769 4663 24803
rect 5733 24769 5767 24803
rect 7757 24769 7791 24803
rect 9505 24769 9539 24803
rect 9597 24769 9631 24803
rect 11069 24769 11103 24803
rect 11161 24769 11195 24803
rect 13001 24769 13035 24803
rect 4997 24701 5031 24735
rect 5549 24701 5583 24735
rect 7481 24701 7515 24735
rect 8953 24701 8987 24735
rect 10425 24701 10459 24735
rect 12909 24701 12943 24735
rect 6653 24633 6687 24667
rect 7573 24633 7607 24667
rect 12173 24633 12207 24667
rect 3709 24565 3743 24599
rect 4169 24565 4203 24599
rect 5089 24565 5123 24599
rect 5457 24565 5491 24599
rect 7113 24565 7147 24599
rect 9045 24565 9079 24599
rect 9413 24565 9447 24599
rect 10057 24565 10091 24599
rect 10977 24565 11011 24599
rect 11897 24565 11931 24599
rect 12449 24565 12483 24599
rect 12817 24565 12851 24599
rect 5181 24361 5215 24395
rect 5733 24361 5767 24395
rect 8309 24361 8343 24395
rect 9137 24361 9171 24395
rect 9965 24361 9999 24395
rect 10241 24361 10275 24395
rect 10701 24361 10735 24395
rect 12725 24361 12759 24395
rect 13001 24361 13035 24395
rect 13185 24361 13219 24395
rect 11222 24293 11256 24327
rect 5825 24225 5859 24259
rect 7196 24225 7230 24259
rect 10977 24225 11011 24259
rect 5917 24157 5951 24191
rect 6929 24157 6963 24191
rect 3157 24021 3191 24055
rect 5365 24021 5399 24055
rect 6469 24021 6503 24055
rect 6837 24021 6871 24055
rect 8677 24021 8711 24055
rect 12357 24021 12391 24055
rect 5181 23817 5215 23851
rect 7021 23817 7055 23851
rect 9965 23817 9999 23851
rect 11529 23817 11563 23851
rect 5825 23749 5859 23783
rect 8585 23749 8619 23783
rect 11897 23749 11931 23783
rect 5273 23681 5307 23715
rect 7481 23681 7515 23715
rect 7573 23681 7607 23715
rect 9045 23681 9079 23715
rect 9229 23681 9263 23715
rect 13093 23681 13127 23715
rect 3065 23613 3099 23647
rect 6285 23613 6319 23647
rect 6653 23613 6687 23647
rect 8493 23613 8527 23647
rect 10149 23613 10183 23647
rect 10405 23613 10439 23647
rect 12173 23613 12207 23647
rect 12909 23613 12943 23647
rect 13461 23613 13495 23647
rect 2973 23545 3007 23579
rect 3310 23545 3344 23579
rect 4813 23545 4847 23579
rect 7389 23545 7423 23579
rect 8125 23545 8159 23579
rect 8953 23545 8987 23579
rect 9689 23545 9723 23579
rect 12817 23545 12851 23579
rect 13829 23545 13863 23579
rect 4445 23477 4479 23511
rect 12449 23477 12483 23511
rect 6469 23273 6503 23307
rect 7573 23273 7607 23307
rect 8033 23273 8067 23307
rect 11069 23273 11103 23307
rect 2329 23205 2363 23239
rect 2789 23205 2823 23239
rect 4436 23205 4470 23239
rect 7941 23205 7975 23239
rect 11345 23205 11379 23239
rect 12602 23205 12636 23239
rect 2881 23137 2915 23171
rect 3893 23137 3927 23171
rect 6837 23137 6871 23171
rect 8401 23137 8435 23171
rect 9945 23137 9979 23171
rect 12357 23137 12391 23171
rect 2973 23069 3007 23103
rect 4169 23069 4203 23103
rect 6929 23069 6963 23103
rect 7021 23069 7055 23103
rect 8493 23069 8527 23103
rect 8677 23069 8711 23103
rect 9689 23069 9723 23103
rect 2421 22933 2455 22967
rect 5549 22933 5583 22967
rect 13737 22933 13771 22967
rect 4353 22729 4387 22763
rect 5365 22729 5399 22763
rect 6193 22729 6227 22763
rect 6561 22729 6595 22763
rect 9597 22729 9631 22763
rect 11437 22729 11471 22763
rect 13001 22729 13035 22763
rect 2789 22661 2823 22695
rect 7205 22661 7239 22695
rect 8769 22661 8803 22695
rect 12633 22661 12667 22695
rect 1593 22593 1627 22627
rect 2329 22593 2363 22627
rect 3433 22593 3467 22627
rect 3801 22593 3835 22627
rect 4261 22593 4295 22627
rect 4813 22593 4847 22627
rect 4997 22593 5031 22627
rect 10241 22593 10275 22627
rect 10609 22593 10643 22627
rect 10977 22593 11011 22627
rect 1409 22525 1443 22559
rect 2697 22525 2731 22559
rect 3157 22525 3191 22559
rect 5825 22525 5859 22559
rect 7389 22525 7423 22559
rect 9413 22525 9447 22559
rect 10057 22525 10091 22559
rect 7634 22457 7668 22491
rect 9045 22457 9079 22491
rect 9965 22457 9999 22491
rect 3249 22389 3283 22423
rect 4721 22389 4755 22423
rect 1685 22185 1719 22219
rect 2789 22185 2823 22219
rect 3249 22185 3283 22219
rect 4721 22185 4755 22219
rect 7573 22117 7607 22151
rect 2513 22049 2547 22083
rect 6173 22049 6207 22083
rect 8033 22049 8067 22083
rect 10057 22049 10091 22083
rect 13461 22049 13495 22083
rect 4813 21981 4847 22015
rect 4997 21981 5031 22015
rect 5917 21981 5951 22015
rect 8125 21981 8159 22015
rect 10149 21981 10183 22015
rect 10241 21981 10275 22015
rect 4353 21913 4387 21947
rect 13645 21913 13679 21947
rect 3893 21845 3927 21879
rect 7297 21845 7331 21879
rect 8585 21845 8619 21879
rect 9689 21845 9723 21879
rect 3893 21641 3927 21675
rect 4813 21641 4847 21675
rect 7297 21641 7331 21675
rect 8861 21641 8895 21675
rect 10241 21641 10275 21675
rect 3617 21573 3651 21607
rect 4353 21505 4387 21539
rect 5457 21505 5491 21539
rect 6653 21505 6687 21539
rect 7849 21505 7883 21539
rect 8401 21505 8435 21539
rect 9321 21505 9355 21539
rect 9505 21505 9539 21539
rect 7665 21437 7699 21471
rect 4721 21369 4755 21403
rect 5181 21369 5215 21403
rect 5273 21301 5307 21335
rect 5917 21301 5951 21335
rect 7205 21301 7239 21335
rect 7757 21301 7791 21335
rect 8677 21301 8711 21335
rect 9229 21301 9263 21335
rect 9873 21301 9907 21335
rect 13461 21301 13495 21335
rect 4445 21097 4479 21131
rect 6101 21097 6135 21131
rect 7389 21097 7423 21131
rect 8217 21097 8251 21131
rect 9965 21097 9999 21131
rect 8861 21029 8895 21063
rect 6469 20961 6503 20995
rect 10508 20961 10542 20995
rect 6561 20893 6595 20927
rect 6745 20893 6779 20927
rect 8309 20893 8343 20927
rect 8401 20893 8435 20927
rect 10241 20893 10275 20927
rect 5917 20825 5951 20859
rect 7849 20825 7883 20859
rect 4813 20757 4847 20791
rect 11621 20757 11655 20791
rect 12541 20757 12575 20791
rect 5825 20553 5859 20587
rect 8217 20553 8251 20587
rect 8493 20553 8527 20587
rect 6837 20417 6871 20451
rect 9321 20417 9355 20451
rect 9781 20417 9815 20451
rect 12909 20417 12943 20451
rect 13001 20417 13035 20451
rect 9689 20349 9723 20383
rect 10048 20349 10082 20383
rect 11437 20349 11471 20383
rect 6469 20281 6503 20315
rect 7082 20281 7116 20315
rect 11897 20281 11931 20315
rect 12817 20281 12851 20315
rect 6101 20213 6135 20247
rect 11161 20213 11195 20247
rect 12265 20213 12299 20247
rect 12449 20213 12483 20247
rect 7205 20009 7239 20043
rect 8309 20009 8343 20043
rect 10333 20009 10367 20043
rect 12541 20009 12575 20043
rect 9965 19873 9999 19907
rect 11417 19873 11451 19907
rect 11161 19805 11195 19839
rect 2789 19669 2823 19703
rect 5089 19669 5123 19703
rect 6929 19669 6963 19703
rect 7941 19669 7975 19703
rect 10609 19669 10643 19703
rect 12909 19669 12943 19703
rect 9965 19465 9999 19499
rect 12449 19465 12483 19499
rect 2789 19329 2823 19363
rect 5549 19329 5583 19363
rect 10517 19329 10551 19363
rect 10609 19329 10643 19363
rect 13001 19329 13035 19363
rect 10425 19261 10459 19295
rect 12173 19261 12207 19295
rect 12817 19261 12851 19295
rect 2697 19193 2731 19227
rect 3056 19193 3090 19227
rect 4905 19193 4939 19227
rect 5457 19193 5491 19227
rect 7481 19193 7515 19227
rect 7573 19193 7607 19227
rect 11805 19193 11839 19227
rect 12909 19193 12943 19227
rect 4169 19125 4203 19159
rect 4537 19125 4571 19159
rect 4997 19125 5031 19159
rect 5365 19125 5399 19159
rect 7021 19125 7055 19159
rect 8861 19125 8895 19159
rect 10057 19125 10091 19159
rect 11253 19125 11287 19159
rect 5917 18921 5951 18955
rect 6745 18921 6779 18955
rect 10701 18921 10735 18955
rect 11437 18921 11471 18955
rect 11989 18921 12023 18955
rect 1685 18853 1719 18887
rect 4506 18853 4540 18887
rect 10149 18853 10183 18887
rect 12449 18853 12483 18887
rect 1409 18785 1443 18819
rect 6653 18785 6687 18819
rect 7113 18785 7147 18819
rect 10057 18785 10091 18819
rect 12357 18785 12391 18819
rect 4261 18717 4295 18751
rect 7205 18717 7239 18751
rect 7389 18717 7423 18751
rect 10333 18717 10367 18751
rect 12541 18717 12575 18751
rect 9137 18649 9171 18683
rect 2973 18581 3007 18615
rect 5641 18581 5675 18615
rect 9689 18581 9723 18615
rect 11069 18581 11103 18615
rect 6653 18377 6687 18411
rect 8493 18377 8527 18411
rect 10149 18377 10183 18411
rect 10609 18377 10643 18411
rect 5089 18309 5123 18343
rect 8217 18309 8251 18343
rect 1593 18241 1627 18275
rect 5641 18241 5675 18275
rect 9597 18241 9631 18275
rect 11161 18241 11195 18275
rect 11713 18241 11747 18275
rect 12449 18241 12483 18275
rect 1409 18173 1443 18207
rect 2881 18173 2915 18207
rect 5457 18173 5491 18207
rect 6837 18173 6871 18207
rect 9505 18173 9539 18207
rect 2237 18105 2271 18139
rect 2789 18105 2823 18139
rect 3126 18105 3160 18139
rect 4905 18105 4939 18139
rect 6285 18105 6319 18139
rect 7082 18105 7116 18139
rect 8861 18105 8895 18139
rect 11069 18105 11103 18139
rect 4261 18037 4295 18071
rect 4537 18037 4571 18071
rect 5549 18037 5583 18071
rect 9045 18037 9079 18071
rect 9413 18037 9447 18071
rect 10517 18037 10551 18071
rect 10977 18037 11011 18071
rect 11989 18037 12023 18071
rect 1593 17833 1627 17867
rect 2789 17833 2823 17867
rect 4353 17833 4387 17867
rect 7573 17833 7607 17867
rect 11069 17833 11103 17867
rect 5610 17765 5644 17799
rect 9505 17765 9539 17799
rect 9956 17765 9990 17799
rect 5273 17697 5307 17731
rect 7941 17697 7975 17731
rect 8033 17697 8067 17731
rect 9689 17697 9723 17731
rect 2881 17629 2915 17663
rect 2973 17629 3007 17663
rect 5365 17629 5399 17663
rect 8125 17629 8159 17663
rect 2421 17493 2455 17527
rect 3893 17493 3927 17527
rect 4905 17493 4939 17527
rect 6745 17493 6779 17527
rect 7205 17493 7239 17527
rect 9045 17493 9079 17527
rect 11345 17493 11379 17527
rect 11989 17493 12023 17527
rect 1777 17289 1811 17323
rect 2881 17289 2915 17323
rect 4445 17289 4479 17323
rect 8493 17289 8527 17323
rect 8861 17289 8895 17323
rect 9873 17289 9907 17323
rect 10609 17289 10643 17323
rect 10793 17289 10827 17323
rect 2513 17221 2547 17255
rect 11805 17221 11839 17255
rect 3433 17153 3467 17187
rect 4997 17153 5031 17187
rect 11345 17153 11379 17187
rect 4353 17085 4387 17119
rect 4813 17085 4847 17119
rect 4905 17085 4939 17119
rect 6653 17085 6687 17119
rect 7113 17085 7147 17119
rect 9321 17085 9355 17119
rect 11161 17085 11195 17119
rect 2145 17017 2179 17051
rect 3341 17017 3375 17051
rect 3985 17017 4019 17051
rect 5825 17017 5859 17051
rect 7380 17017 7414 17051
rect 9137 17017 9171 17051
rect 3249 16949 3283 16983
rect 5549 16949 5583 16983
rect 10333 16949 10367 16983
rect 11253 16949 11287 16983
rect 2513 16745 2547 16779
rect 2973 16745 3007 16779
rect 3249 16745 3283 16779
rect 4077 16745 4111 16779
rect 4445 16745 4479 16779
rect 5273 16745 5307 16779
rect 7849 16745 7883 16779
rect 8953 16745 8987 16779
rect 10241 16745 10275 16779
rect 11253 16745 11287 16779
rect 13185 16745 13219 16779
rect 4537 16677 4571 16711
rect 6377 16677 6411 16711
rect 7665 16677 7699 16711
rect 10149 16677 10183 16711
rect 6285 16609 6319 16643
rect 8217 16609 8251 16643
rect 8309 16609 8343 16643
rect 9229 16609 9263 16643
rect 10609 16609 10643 16643
rect 10701 16609 10735 16643
rect 11805 16609 11839 16643
rect 12061 16609 12095 16643
rect 4629 16541 4663 16575
rect 6561 16541 6595 16575
rect 8401 16541 8435 16575
rect 10793 16541 10827 16575
rect 7205 16473 7239 16507
rect 5641 16405 5675 16439
rect 5917 16405 5951 16439
rect 3801 16201 3835 16235
rect 4169 16201 4203 16235
rect 6193 16201 6227 16235
rect 10793 16201 10827 16235
rect 12173 16201 12207 16235
rect 5733 16065 5767 16099
rect 7665 16065 7699 16099
rect 8217 16065 8251 16099
rect 9321 16065 9355 16099
rect 9965 16065 9999 16099
rect 11345 16065 11379 16099
rect 11805 16065 11839 16099
rect 5549 15997 5583 16031
rect 7481 15997 7515 16031
rect 7573 15997 7607 16031
rect 9137 15997 9171 16031
rect 5089 15929 5123 15963
rect 6653 15929 6687 15963
rect 8585 15929 8619 15963
rect 9045 15929 9079 15963
rect 10333 15929 10367 15963
rect 11161 15929 11195 15963
rect 4445 15861 4479 15895
rect 5181 15861 5215 15895
rect 5641 15861 5675 15895
rect 7113 15861 7147 15895
rect 8677 15861 8711 15895
rect 10701 15861 10735 15895
rect 11253 15861 11287 15895
rect 4077 15657 4111 15691
rect 5181 15657 5215 15691
rect 6009 15657 6043 15691
rect 6837 15657 6871 15691
rect 7573 15657 7607 15691
rect 7849 15657 7883 15691
rect 8217 15657 8251 15691
rect 8953 15657 8987 15691
rect 9965 15657 9999 15691
rect 10517 15657 10551 15691
rect 4445 15589 4479 15623
rect 6101 15589 6135 15623
rect 9229 15589 9263 15623
rect 10333 15589 10367 15623
rect 10885 15589 10919 15623
rect 4537 15521 4571 15555
rect 7205 15521 7239 15555
rect 8309 15521 8343 15555
rect 4629 15453 4663 15487
rect 6285 15453 6319 15487
rect 8493 15453 8527 15487
rect 10977 15453 11011 15487
rect 11161 15453 11195 15487
rect 5549 15385 5583 15419
rect 3249 15317 3283 15351
rect 5641 15317 5675 15351
rect 3157 15113 3191 15147
rect 6837 15113 6871 15147
rect 8309 15113 8343 15147
rect 8677 15113 8711 15147
rect 10057 15113 10091 15147
rect 10517 15113 10551 15147
rect 11897 15113 11931 15147
rect 6193 15045 6227 15079
rect 7941 15045 7975 15079
rect 1593 14977 1627 15011
rect 3065 14977 3099 15011
rect 3801 14977 3835 15011
rect 4997 14977 5031 15011
rect 5733 14977 5767 15011
rect 7389 14977 7423 15011
rect 9137 14977 9171 15011
rect 9321 14977 9355 15011
rect 11161 14977 11195 15011
rect 13553 14977 13587 15011
rect 1409 14909 1443 14943
rect 5549 14909 5583 14943
rect 7205 14909 7239 14943
rect 11529 14909 11563 14943
rect 13277 14909 13311 14943
rect 2237 14841 2271 14875
rect 6653 14841 6687 14875
rect 7297 14841 7331 14875
rect 10977 14841 11011 14875
rect 14013 14841 14047 14875
rect 3525 14773 3559 14807
rect 3617 14773 3651 14807
rect 4261 14773 4295 14807
rect 4629 14773 4663 14807
rect 5181 14773 5215 14807
rect 5641 14773 5675 14807
rect 9045 14773 9079 14807
rect 10333 14773 10367 14807
rect 10885 14773 10919 14807
rect 3249 14569 3283 14603
rect 4077 14569 4111 14603
rect 6009 14569 6043 14603
rect 7297 14569 7331 14603
rect 8493 14569 8527 14603
rect 9689 14569 9723 14603
rect 10057 14569 10091 14603
rect 11161 14569 11195 14603
rect 12909 14569 12943 14603
rect 6101 14501 6135 14535
rect 6929 14501 6963 14535
rect 4445 14433 4479 14467
rect 4537 14433 4571 14467
rect 5181 14433 5215 14467
rect 7941 14433 7975 14467
rect 8861 14433 8895 14467
rect 11529 14433 11563 14467
rect 11796 14433 11830 14467
rect 4629 14365 4663 14399
rect 5549 14365 5583 14399
rect 6193 14365 6227 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 2421 14297 2455 14331
rect 3893 14297 3927 14331
rect 5641 14229 5675 14263
rect 9505 14229 9539 14263
rect 10701 14229 10735 14263
rect 2329 14025 2363 14059
rect 5273 14025 5307 14059
rect 6009 14025 6043 14059
rect 6377 14025 6411 14059
rect 7021 14025 7055 14059
rect 8309 14025 8343 14059
rect 9689 14025 9723 14059
rect 10057 14025 10091 14059
rect 11069 14025 11103 14059
rect 12173 14025 12207 14059
rect 2973 13889 3007 13923
rect 3433 13889 3467 13923
rect 8033 13889 8067 13923
rect 9137 13889 9171 13923
rect 10517 13889 10551 13923
rect 10701 13889 10735 13923
rect 2697 13821 2731 13855
rect 3893 13821 3927 13855
rect 4160 13821 4194 13855
rect 8861 13821 8895 13855
rect 8953 13821 8987 13855
rect 11529 13821 11563 13855
rect 11897 13821 11931 13855
rect 2237 13753 2271 13787
rect 3801 13753 3835 13787
rect 2789 13685 2823 13719
rect 5733 13685 5767 13719
rect 8493 13685 8527 13719
rect 10425 13685 10459 13719
rect 2421 13481 2455 13515
rect 4629 13481 4663 13515
rect 8861 13481 8895 13515
rect 9505 13481 9539 13515
rect 1685 13413 1719 13447
rect 4353 13413 4387 13447
rect 5172 13413 5206 13447
rect 9934 13413 9968 13447
rect 1409 13345 1443 13379
rect 7113 13345 7147 13379
rect 7380 13345 7414 13379
rect 4905 13277 4939 13311
rect 9689 13277 9723 13311
rect 6929 13209 6963 13243
rect 3801 13141 3835 13175
rect 6285 13141 6319 13175
rect 6653 13141 6687 13175
rect 8493 13141 8527 13175
rect 11069 13141 11103 13175
rect 3893 12937 3927 12971
rect 4997 12937 5031 12971
rect 5917 12937 5951 12971
rect 8217 12937 8251 12971
rect 8493 12937 8527 12971
rect 10701 12937 10735 12971
rect 11161 12937 11195 12971
rect 5273 12869 5307 12903
rect 2513 12733 2547 12767
rect 6837 12733 6871 12767
rect 9045 12733 9079 12767
rect 2421 12665 2455 12699
rect 2758 12665 2792 12699
rect 6285 12665 6319 12699
rect 7104 12665 7138 12699
rect 9290 12665 9324 12699
rect 1685 12597 1719 12631
rect 6561 12597 6595 12631
rect 8861 12597 8895 12631
rect 10425 12597 10459 12631
rect 4905 12393 4939 12427
rect 6469 12393 6503 12427
rect 8493 12393 8527 12427
rect 10149 12393 10183 12427
rect 12449 12393 12483 12427
rect 5089 12257 5123 12291
rect 6837 12257 6871 12291
rect 8401 12257 8435 12291
rect 10885 12257 10919 12291
rect 11325 12257 11359 12291
rect 6929 12189 6963 12223
rect 7021 12189 7055 12223
rect 7941 12189 7975 12223
rect 8585 12189 8619 12223
rect 9689 12189 9723 12223
rect 11069 12189 11103 12223
rect 9137 12121 9171 12155
rect 2513 12053 2547 12087
rect 5457 12053 5491 12087
rect 6009 12053 6043 12087
rect 6377 12053 6411 12087
rect 7573 12053 7607 12087
rect 8033 12053 8067 12087
rect 10517 12053 10551 12087
rect 10701 12053 10735 12087
rect 4353 11849 4387 11883
rect 6561 11849 6595 11883
rect 6929 11849 6963 11883
rect 8033 11849 8067 11883
rect 10057 11849 10091 11883
rect 11437 11849 11471 11883
rect 11805 11849 11839 11883
rect 4721 11781 4755 11815
rect 8493 11781 8527 11815
rect 1593 11713 1627 11747
rect 5733 11713 5767 11747
rect 7389 11713 7423 11747
rect 7573 11713 7607 11747
rect 9045 11713 9079 11747
rect 10701 11713 10735 11747
rect 1409 11645 1443 11679
rect 5549 11645 5583 11679
rect 5641 11645 5675 11679
rect 7297 11645 7331 11679
rect 10425 11645 10459 11679
rect 9965 11577 9999 11611
rect 2237 11509 2271 11543
rect 4997 11509 5031 11543
rect 5181 11509 5215 11543
rect 8401 11509 8435 11543
rect 8861 11509 8895 11543
rect 8953 11509 8987 11543
rect 9597 11509 9631 11543
rect 10517 11509 10551 11543
rect 11161 11509 11195 11543
rect 4813 11305 4847 11339
rect 5181 11305 5215 11339
rect 6377 11305 6411 11339
rect 6837 11305 6871 11339
rect 7849 11305 7883 11339
rect 8033 11305 8067 11339
rect 8493 11305 8527 11339
rect 9045 11305 9079 11339
rect 10057 11305 10091 11339
rect 10793 11305 10827 11339
rect 4721 11237 4755 11271
rect 5273 11237 5307 11271
rect 5917 11237 5951 11271
rect 8401 11237 8435 11271
rect 10701 11237 10735 11271
rect 1409 11169 1443 11203
rect 6745 11169 6779 11203
rect 11161 11169 11195 11203
rect 1593 11101 1627 11135
rect 5365 11101 5399 11135
rect 6929 11101 6963 11135
rect 8585 11101 8619 11135
rect 11253 11101 11287 11135
rect 11437 11101 11471 11135
rect 12357 11101 12391 11135
rect 6193 11033 6227 11067
rect 2237 10965 2271 10999
rect 7481 10965 7515 10999
rect 3985 10761 4019 10795
rect 4721 10761 4755 10795
rect 5181 10761 5215 10795
rect 7021 10761 7055 10795
rect 8585 10761 8619 10795
rect 9689 10761 9723 10795
rect 10609 10761 10643 10795
rect 10793 10761 10827 10795
rect 12449 10761 12483 10795
rect 8125 10693 8159 10727
rect 12265 10693 12299 10727
rect 2053 10625 2087 10659
rect 2697 10625 2731 10659
rect 4353 10625 4387 10659
rect 5733 10625 5767 10659
rect 7481 10625 7515 10659
rect 7573 10625 7607 10659
rect 9137 10625 9171 10659
rect 11253 10625 11287 10659
rect 11345 10625 11379 10659
rect 11805 10625 11839 10659
rect 13001 10625 13035 10659
rect 5089 10557 5123 10591
rect 5641 10557 5675 10591
rect 9045 10557 9079 10591
rect 10333 10557 10367 10591
rect 11161 10557 11195 10591
rect 12817 10557 12851 10591
rect 1685 10489 1719 10523
rect 2605 10489 2639 10523
rect 12909 10489 12943 10523
rect 2145 10421 2179 10455
rect 2513 10421 2547 10455
rect 5549 10421 5583 10455
rect 6377 10421 6411 10455
rect 7389 10421 7423 10455
rect 8493 10421 8527 10455
rect 8953 10421 8987 10455
rect 1685 10217 1719 10251
rect 3157 10217 3191 10251
rect 4077 10217 4111 10251
rect 5273 10217 5307 10251
rect 5917 10217 5951 10251
rect 6469 10217 6503 10251
rect 7113 10217 7147 10251
rect 7481 10217 7515 10251
rect 8125 10217 8159 10251
rect 8953 10217 8987 10251
rect 10241 10217 10275 10251
rect 11713 10217 11747 10251
rect 6929 10149 6963 10183
rect 8677 10149 8711 10183
rect 10600 10149 10634 10183
rect 12817 10149 12851 10183
rect 2044 10081 2078 10115
rect 3525 10081 3559 10115
rect 4445 10081 4479 10115
rect 5825 10081 5859 10115
rect 10333 10081 10367 10115
rect 1777 10013 1811 10047
rect 3893 10013 3927 10047
rect 4537 10013 4571 10047
rect 4629 10013 4663 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 5641 9945 5675 9979
rect 9321 9877 9355 9911
rect 12449 9877 12483 9911
rect 4997 9673 5031 9707
rect 7205 9673 7239 9707
rect 7757 9673 7791 9707
rect 1869 9605 1903 9639
rect 4169 9605 4203 9639
rect 6653 9605 6687 9639
rect 8861 9605 8895 9639
rect 10885 9605 10919 9639
rect 11161 9605 11195 9639
rect 5549 9537 5583 9571
rect 6009 9537 6043 9571
rect 8217 9537 8251 9571
rect 8401 9537 8435 9571
rect 10425 9537 10459 9571
rect 2329 9469 2363 9503
rect 2789 9469 2823 9503
rect 9505 9469 9539 9503
rect 9781 9469 9815 9503
rect 3056 9401 3090 9435
rect 5457 9401 5491 9435
rect 9137 9401 9171 9435
rect 2697 9333 2731 9367
rect 4537 9333 4571 9367
rect 4905 9333 4939 9367
rect 5365 9333 5399 9367
rect 7665 9333 7699 9367
rect 8125 9333 8159 9367
rect 9321 9333 9355 9367
rect 1777 9129 1811 9163
rect 2329 9129 2363 9163
rect 2881 9129 2915 9163
rect 4077 9129 4111 9163
rect 5641 9129 5675 9163
rect 6101 9129 6135 9163
rect 6929 9129 6963 9163
rect 7297 9129 7331 9163
rect 9689 9129 9723 9163
rect 10057 9129 10091 9163
rect 10149 9129 10183 9163
rect 2789 9061 2823 9095
rect 3893 8993 3927 9027
rect 4445 8993 4479 9027
rect 6009 8993 6043 9027
rect 7656 8993 7690 9027
rect 3065 8925 3099 8959
rect 3433 8925 3467 8959
rect 4537 8925 4571 8959
rect 4721 8925 4755 8959
rect 5089 8925 5123 8959
rect 6193 8925 6227 8959
rect 7389 8925 7423 8959
rect 10241 8925 10275 8959
rect 5457 8857 5491 8891
rect 8769 8857 8803 8891
rect 2421 8789 2455 8823
rect 9229 8789 9263 8823
rect 2513 8585 2547 8619
rect 4169 8585 4203 8619
rect 5641 8585 5675 8619
rect 6469 8585 6503 8619
rect 6009 8517 6043 8551
rect 1593 8449 1627 8483
rect 3249 8449 3283 8483
rect 1409 8381 1443 8415
rect 4261 8381 4295 8415
rect 6653 8381 6687 8415
rect 6837 8381 6871 8415
rect 7104 8381 7138 8415
rect 9137 8381 9171 8415
rect 9393 8381 9427 8415
rect 3065 8313 3099 8347
rect 3801 8313 3835 8347
rect 4528 8313 4562 8347
rect 6285 8313 6319 8347
rect 9045 8313 9079 8347
rect 2697 8245 2731 8279
rect 3157 8245 3191 8279
rect 8217 8245 8251 8279
rect 8677 8245 8711 8279
rect 10517 8245 10551 8279
rect 1685 8041 1719 8075
rect 2421 8041 2455 8075
rect 2881 8041 2915 8075
rect 3893 8041 3927 8075
rect 4353 8041 4387 8075
rect 6745 8041 6779 8075
rect 7481 8041 7515 8075
rect 10241 8041 10275 8075
rect 2329 7973 2363 8007
rect 4905 7973 4939 8007
rect 7113 7973 7147 8007
rect 7941 7973 7975 8007
rect 9413 7973 9447 8007
rect 9965 7973 9999 8007
rect 2789 7905 2823 7939
rect 5621 7905 5655 7939
rect 8401 7905 8435 7939
rect 10609 7905 10643 7939
rect 11233 7905 11267 7939
rect 3065 7837 3099 7871
rect 5365 7837 5399 7871
rect 8493 7837 8527 7871
rect 8677 7837 8711 7871
rect 10977 7837 11011 7871
rect 3525 7701 3559 7735
rect 8033 7701 8067 7735
rect 9137 7701 9171 7735
rect 10425 7701 10459 7735
rect 12357 7701 12391 7735
rect 2789 7497 2823 7531
rect 3157 7497 3191 7531
rect 4721 7497 4755 7531
rect 5457 7497 5491 7531
rect 6193 7497 6227 7531
rect 6653 7497 6687 7531
rect 7849 7497 7883 7531
rect 10517 7497 10551 7531
rect 11069 7497 11103 7531
rect 2513 7429 2547 7463
rect 8769 7429 8803 7463
rect 8953 7429 8987 7463
rect 8493 7361 8527 7395
rect 4997 7293 5031 7327
rect 5641 7293 5675 7327
rect 7389 7293 7423 7327
rect 10057 7361 10091 7395
rect 8217 7225 8251 7259
rect 8769 7225 8803 7259
rect 9873 7225 9907 7259
rect 4353 7157 4387 7191
rect 4813 7157 4847 7191
rect 5825 7157 5859 7191
rect 7757 7157 7791 7191
rect 8309 7157 8343 7191
rect 9229 7157 9263 7191
rect 9413 7157 9447 7191
rect 9781 7157 9815 7191
rect 11345 7157 11379 7191
rect 2145 6953 2179 6987
rect 7205 6953 7239 6987
rect 8493 6953 8527 6987
rect 10241 6953 10275 6987
rect 7941 6885 7975 6919
rect 1409 6817 1443 6851
rect 2513 6817 2547 6851
rect 5089 6817 5123 6851
rect 6193 6817 6227 6851
rect 7573 6817 7607 6851
rect 8401 6817 8435 6851
rect 9689 6817 9723 6851
rect 11069 6817 11103 6851
rect 11325 6817 11359 6851
rect 8677 6749 8711 6783
rect 2697 6681 2731 6715
rect 6377 6681 6411 6715
rect 9413 6681 9447 6715
rect 1593 6613 1627 6647
rect 5273 6613 5307 6647
rect 5733 6613 5767 6647
rect 8033 6613 8067 6647
rect 9873 6613 9907 6647
rect 12449 6613 12483 6647
rect 1593 6409 1627 6443
rect 2605 6409 2639 6443
rect 5089 6409 5123 6443
rect 5549 6409 5583 6443
rect 6193 6409 6227 6443
rect 6653 6409 6687 6443
rect 7573 6409 7607 6443
rect 9597 6409 9631 6443
rect 11069 6409 11103 6443
rect 2237 6341 2271 6375
rect 4721 6341 4755 6375
rect 7941 6341 7975 6375
rect 9137 6341 9171 6375
rect 8677 6273 8711 6307
rect 10241 6273 10275 6307
rect 2053 6205 2087 6239
rect 4445 6205 4479 6239
rect 4537 6205 4571 6239
rect 5641 6205 5675 6239
rect 6929 6205 6963 6239
rect 8401 6205 8435 6239
rect 9965 6205 9999 6239
rect 10609 6205 10643 6239
rect 11161 6205 11195 6239
rect 11713 6205 11747 6239
rect 5825 6069 5859 6103
rect 7113 6069 7147 6103
rect 8033 6069 8067 6103
rect 8493 6069 8527 6103
rect 9505 6069 9539 6103
rect 10057 6069 10091 6103
rect 11345 6069 11379 6103
rect 6285 5865 6319 5899
rect 7849 5865 7883 5899
rect 9689 5865 9723 5899
rect 10793 5865 10827 5899
rect 11069 5865 11103 5899
rect 11345 5865 11379 5899
rect 7389 5797 7423 5831
rect 8861 5797 8895 5831
rect 10149 5797 10183 5831
rect 2145 5729 2179 5763
rect 5089 5729 5123 5763
rect 6377 5729 6411 5763
rect 10057 5729 10091 5763
rect 11713 5729 11747 5763
rect 4629 5661 4663 5695
rect 5181 5661 5215 5695
rect 5273 5661 5307 5695
rect 7941 5661 7975 5695
rect 8125 5661 8159 5695
rect 10241 5661 10275 5695
rect 11805 5661 11839 5695
rect 11989 5661 12023 5695
rect 6561 5593 6595 5627
rect 7481 5593 7515 5627
rect 9413 5593 9447 5627
rect 2329 5525 2363 5559
rect 3433 5525 3467 5559
rect 4721 5525 4755 5559
rect 5917 5525 5951 5559
rect 7021 5525 7055 5559
rect 8585 5525 8619 5559
rect 4813 5321 4847 5355
rect 5181 5321 5215 5355
rect 5549 5321 5583 5355
rect 6469 5321 6503 5355
rect 8585 5321 8619 5355
rect 10425 5321 10459 5355
rect 12173 5321 12207 5355
rect 2973 5253 3007 5287
rect 11437 5253 11471 5287
rect 2329 5185 2363 5219
rect 2053 5117 2087 5151
rect 2145 5117 2179 5151
rect 3433 5117 3467 5151
rect 5641 5117 5675 5151
rect 6837 5117 6871 5151
rect 7104 5117 7138 5151
rect 9045 5117 9079 5151
rect 11253 5117 11287 5151
rect 11805 5117 11839 5151
rect 3341 5049 3375 5083
rect 3700 5049 3734 5083
rect 9290 5049 9324 5083
rect 10793 5049 10827 5083
rect 5825 4981 5859 5015
rect 8217 4981 8251 5015
rect 8861 4981 8895 5015
rect 11161 4981 11195 5015
rect 12449 4981 12483 5015
rect 2421 4777 2455 4811
rect 2789 4777 2823 4811
rect 6009 4777 6043 4811
rect 6377 4777 6411 4811
rect 8585 4777 8619 4811
rect 9965 4777 9999 4811
rect 11805 4777 11839 4811
rect 1961 4709 1995 4743
rect 2881 4709 2915 4743
rect 6745 4709 6779 4743
rect 7104 4709 7138 4743
rect 11713 4709 11747 4743
rect 12265 4709 12299 4743
rect 4537 4641 4571 4675
rect 4885 4641 4919 4675
rect 10609 4641 10643 4675
rect 11345 4641 11379 4675
rect 12173 4641 12207 4675
rect 12817 4641 12851 4675
rect 2329 4573 2363 4607
rect 3065 4573 3099 4607
rect 4629 4573 4663 4607
rect 6837 4573 6871 4607
rect 10701 4573 10735 4607
rect 10885 4573 10919 4607
rect 12449 4573 12483 4607
rect 13369 4573 13403 4607
rect 3893 4505 3927 4539
rect 9413 4505 9447 4539
rect 10241 4505 10275 4539
rect 3525 4437 3559 4471
rect 8217 4437 8251 4471
rect 9045 4437 9079 4471
rect 2513 4233 2547 4267
rect 4353 4233 4387 4267
rect 5181 4233 5215 4267
rect 6193 4233 6227 4267
rect 6469 4233 6503 4267
rect 6837 4233 6871 4267
rect 8401 4233 8435 4267
rect 10977 4233 11011 4267
rect 12449 4233 12483 4267
rect 1593 4097 1627 4131
rect 2973 4097 3007 4131
rect 4721 4097 4755 4131
rect 5825 4097 5859 4131
rect 1409 4029 1443 4063
rect 3240 4029 3274 4063
rect 5089 4029 5123 4063
rect 5549 4029 5583 4063
rect 11805 4165 11839 4199
rect 12173 4165 12207 4199
rect 7481 4097 7515 4131
rect 8953 4097 8987 4131
rect 9873 4097 9907 4131
rect 10425 4097 10459 4131
rect 10517 4097 10551 4131
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 6653 4029 6687 4063
rect 8309 4029 8343 4063
rect 8861 4029 8895 4063
rect 2881 3961 2915 3995
rect 6469 3961 6503 3995
rect 7941 3961 7975 3995
rect 8769 3961 8803 3995
rect 12817 3961 12851 3995
rect 13461 3961 13495 3995
rect 5641 3893 5675 3927
rect 7205 3893 7239 3927
rect 7297 3893 7331 3927
rect 9413 3893 9447 3927
rect 9965 3893 9999 3927
rect 10333 3893 10367 3927
rect 11345 3893 11379 3927
rect 1593 3689 1627 3723
rect 2421 3689 2455 3723
rect 3433 3689 3467 3723
rect 3893 3689 3927 3723
rect 5181 3689 5215 3723
rect 6653 3689 6687 3723
rect 7573 3689 7607 3723
rect 8033 3689 8067 3723
rect 8401 3689 8435 3723
rect 9045 3689 9079 3723
rect 9873 3689 9907 3723
rect 10885 3689 10919 3723
rect 11253 3689 11287 3723
rect 12817 3689 12851 3723
rect 2789 3621 2823 3655
rect 6285 3621 6319 3655
rect 10333 3621 10367 3655
rect 11682 3621 11716 3655
rect 4077 3553 4111 3587
rect 4629 3553 4663 3587
rect 5549 3553 5583 3587
rect 6745 3553 6779 3587
rect 10241 3553 10275 3587
rect 2329 3485 2363 3519
rect 2881 3485 2915 3519
rect 3065 3485 3099 3519
rect 5641 3485 5675 3519
rect 5825 3485 5859 3519
rect 8493 3485 8527 3519
rect 8585 3485 8619 3519
rect 10425 3485 10459 3519
rect 11437 3485 11471 3519
rect 4261 3349 4295 3383
rect 4997 3349 5031 3383
rect 6929 3349 6963 3383
rect 7849 3349 7883 3383
rect 9505 3349 9539 3383
rect 13093 3349 13127 3383
rect 1961 3145 1995 3179
rect 4905 3145 4939 3179
rect 6285 3145 6319 3179
rect 7021 3145 7055 3179
rect 8953 3145 8987 3179
rect 9689 3145 9723 3179
rect 11161 3145 11195 3179
rect 12449 3145 12483 3179
rect 4445 3077 4479 3111
rect 4721 3077 4755 3111
rect 6009 3077 6043 3111
rect 1409 3009 1443 3043
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
rect 9229 3009 9263 3043
rect 13093 3009 13127 3043
rect 13461 3009 13495 3043
rect 2421 2941 2455 2975
rect 5273 2941 5307 2975
rect 7573 2941 7607 2975
rect 7829 2941 7863 2975
rect 9781 2941 9815 2975
rect 11897 2941 11931 2975
rect 12909 2941 12943 2975
rect 2237 2873 2271 2907
rect 2666 2873 2700 2907
rect 7389 2873 7423 2907
rect 10026 2873 10060 2907
rect 11437 2873 11471 2907
rect 12817 2873 12851 2907
rect 3801 2805 3835 2839
rect 12265 2805 12299 2839
rect 1685 2601 1719 2635
rect 2421 2601 2455 2635
rect 4353 2601 4387 2635
rect 4629 2601 4663 2635
rect 5181 2601 5215 2635
rect 5825 2601 5859 2635
rect 7573 2601 7607 2635
rect 8125 2601 8159 2635
rect 8493 2601 8527 2635
rect 9597 2601 9631 2635
rect 10057 2601 10091 2635
rect 10701 2601 10735 2635
rect 11161 2601 11195 2635
rect 12081 2601 12115 2635
rect 13001 2601 13035 2635
rect 13093 2601 13127 2635
rect 3893 2533 3927 2567
rect 5273 2533 5307 2567
rect 8033 2533 8067 2567
rect 14013 2533 14047 2567
rect 1777 2465 1811 2499
rect 2881 2465 2915 2499
rect 3433 2465 3467 2499
rect 6745 2465 6779 2499
rect 6929 2465 6963 2499
rect 8585 2465 8619 2499
rect 10609 2465 10643 2499
rect 11069 2465 11103 2499
rect 12449 2465 12483 2499
rect 2789 2397 2823 2431
rect 5457 2397 5491 2431
rect 6377 2397 6411 2431
rect 8677 2397 8711 2431
rect 9229 2397 9263 2431
rect 11253 2397 11287 2431
rect 13185 2397 13219 2431
rect 13645 2397 13679 2431
rect 1961 2329 1995 2363
rect 4813 2329 4847 2363
rect 12633 2329 12667 2363
rect 3065 2261 3099 2295
rect 7113 2261 7147 2295
<< metal1 >>
rect 11330 37816 11336 37868
rect 11388 37856 11394 37868
rect 12250 37856 12256 37868
rect 11388 37828 12256 37856
rect 11388 37816 11394 37828
rect 12250 37816 12256 37828
rect 12308 37816 12314 37868
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 13906 37136 13912 37188
rect 13964 37176 13970 37188
rect 14550 37176 14556 37188
rect 13964 37148 14556 37176
rect 13964 37136 13970 37148
rect 14550 37136 14556 37148
rect 14608 37136 14614 37188
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 7282 36360 7288 36372
rect 7243 36332 7288 36360
rect 7282 36320 7288 36332
rect 7340 36320 7346 36372
rect 7101 36227 7159 36233
rect 7101 36193 7113 36227
rect 7147 36224 7159 36227
rect 7190 36224 7196 36236
rect 7147 36196 7196 36224
rect 7147 36193 7159 36196
rect 7101 36187 7159 36193
rect 7190 36184 7196 36196
rect 7248 36184 7254 36236
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 4982 35776 4988 35828
rect 5040 35816 5046 35828
rect 5353 35819 5411 35825
rect 5353 35816 5365 35819
rect 5040 35788 5365 35816
rect 5040 35776 5046 35788
rect 5353 35785 5365 35788
rect 5399 35785 5411 35819
rect 5353 35779 5411 35785
rect 6914 35776 6920 35828
rect 6972 35816 6978 35828
rect 7285 35819 7343 35825
rect 7285 35816 7297 35819
rect 6972 35788 7297 35816
rect 6972 35776 6978 35788
rect 7285 35785 7297 35788
rect 7331 35785 7343 35819
rect 7285 35779 7343 35785
rect 5169 35615 5227 35621
rect 5169 35581 5181 35615
rect 5215 35612 5227 35615
rect 7101 35615 7159 35621
rect 5215 35584 5856 35612
rect 5215 35581 5227 35584
rect 5169 35575 5227 35581
rect 5828 35485 5856 35584
rect 7101 35581 7113 35615
rect 7147 35612 7159 35615
rect 7282 35612 7288 35624
rect 7147 35584 7288 35612
rect 7147 35581 7159 35584
rect 7101 35575 7159 35581
rect 7282 35572 7288 35584
rect 7340 35572 7346 35624
rect 5813 35479 5871 35485
rect 5813 35445 5825 35479
rect 5859 35476 5871 35479
rect 5994 35476 6000 35488
rect 5859 35448 6000 35476
rect 5859 35445 5871 35448
rect 5813 35439 5871 35445
rect 5994 35436 6000 35448
rect 6052 35436 6058 35488
rect 7190 35436 7196 35488
rect 7248 35476 7254 35488
rect 7745 35479 7803 35485
rect 7745 35476 7757 35479
rect 7248 35448 7757 35476
rect 7248 35436 7254 35448
rect 7745 35445 7757 35448
rect 7791 35476 7803 35479
rect 8202 35476 8208 35488
rect 7791 35448 8208 35476
rect 7791 35445 7803 35448
rect 7745 35439 7803 35445
rect 8202 35436 8208 35448
rect 8260 35436 8266 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 3053 35275 3111 35281
rect 3053 35241 3065 35275
rect 3099 35272 3111 35275
rect 3326 35272 3332 35284
rect 3099 35244 3332 35272
rect 3099 35241 3111 35244
rect 3053 35235 3111 35241
rect 3326 35232 3332 35244
rect 3384 35232 3390 35284
rect 4246 35272 4252 35284
rect 4207 35244 4252 35272
rect 4246 35232 4252 35244
rect 4304 35232 4310 35284
rect 5353 35275 5411 35281
rect 5353 35241 5365 35275
rect 5399 35272 5411 35275
rect 5442 35272 5448 35284
rect 5399 35244 5448 35272
rect 5399 35241 5411 35244
rect 5353 35235 5411 35241
rect 5442 35232 5448 35244
rect 5500 35232 5506 35284
rect 6549 35275 6607 35281
rect 6549 35241 6561 35275
rect 6595 35272 6607 35275
rect 6638 35272 6644 35284
rect 6595 35244 6644 35272
rect 6595 35241 6607 35244
rect 6549 35235 6607 35241
rect 6638 35232 6644 35244
rect 6696 35232 6702 35284
rect 7374 35232 7380 35284
rect 7432 35272 7438 35284
rect 7653 35275 7711 35281
rect 7653 35272 7665 35275
rect 7432 35244 7665 35272
rect 7432 35232 7438 35244
rect 7653 35241 7665 35244
rect 7699 35241 7711 35275
rect 7653 35235 7711 35241
rect 2869 35139 2927 35145
rect 2869 35105 2881 35139
rect 2915 35136 2927 35139
rect 3050 35136 3056 35148
rect 2915 35108 3056 35136
rect 2915 35105 2927 35108
rect 2869 35099 2927 35105
rect 3050 35096 3056 35108
rect 3108 35096 3114 35148
rect 4065 35139 4123 35145
rect 4065 35105 4077 35139
rect 4111 35136 4123 35139
rect 4246 35136 4252 35148
rect 4111 35108 4252 35136
rect 4111 35105 4123 35108
rect 4065 35099 4123 35105
rect 4246 35096 4252 35108
rect 4304 35096 4310 35148
rect 5166 35136 5172 35148
rect 5127 35108 5172 35136
rect 5166 35096 5172 35108
rect 5224 35096 5230 35148
rect 6365 35139 6423 35145
rect 6365 35105 6377 35139
rect 6411 35136 6423 35139
rect 6822 35136 6828 35148
rect 6411 35108 6828 35136
rect 6411 35105 6423 35108
rect 6365 35099 6423 35105
rect 6822 35096 6828 35108
rect 6880 35096 6886 35148
rect 7466 35136 7472 35148
rect 7427 35108 7472 35136
rect 7466 35096 7472 35108
rect 7524 35096 7530 35148
rect 11146 35096 11152 35148
rect 11204 35136 11210 35148
rect 11313 35139 11371 35145
rect 11313 35136 11325 35139
rect 11204 35108 11325 35136
rect 11204 35096 11210 35108
rect 11313 35105 11325 35108
rect 11359 35105 11371 35139
rect 11313 35099 11371 35105
rect 11057 35071 11115 35077
rect 11057 35068 11069 35071
rect 10060 35040 11069 35068
rect 10060 34944 10088 35040
rect 11057 35037 11069 35040
rect 11103 35037 11115 35071
rect 11057 35031 11115 35037
rect 7193 34935 7251 34941
rect 7193 34901 7205 34935
rect 7239 34932 7251 34935
rect 7282 34932 7288 34944
rect 7239 34904 7288 34932
rect 7239 34901 7251 34904
rect 7193 34895 7251 34901
rect 7282 34892 7288 34904
rect 7340 34892 7346 34944
rect 8110 34932 8116 34944
rect 8071 34904 8116 34932
rect 8110 34892 8116 34904
rect 8168 34892 8174 34944
rect 10042 34932 10048 34944
rect 10003 34904 10048 34932
rect 10042 34892 10048 34904
rect 10100 34892 10106 34944
rect 12437 34935 12495 34941
rect 12437 34901 12449 34935
rect 12483 34932 12495 34935
rect 12526 34932 12532 34944
rect 12483 34904 12532 34932
rect 12483 34901 12495 34904
rect 12437 34895 12495 34901
rect 12526 34892 12532 34904
rect 12584 34892 12590 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 566 34688 572 34740
rect 624 34728 630 34740
rect 1581 34731 1639 34737
rect 1581 34728 1593 34731
rect 624 34700 1593 34728
rect 624 34688 630 34700
rect 1581 34697 1593 34700
rect 1627 34697 1639 34731
rect 1581 34691 1639 34697
rect 2958 34688 2964 34740
rect 3016 34728 3022 34740
rect 3789 34731 3847 34737
rect 3789 34728 3801 34731
rect 3016 34700 3801 34728
rect 3016 34688 3022 34700
rect 3789 34697 3801 34700
rect 3835 34697 3847 34731
rect 4246 34728 4252 34740
rect 4207 34700 4252 34728
rect 3789 34691 3847 34697
rect 4246 34688 4252 34700
rect 4304 34688 4310 34740
rect 5721 34731 5779 34737
rect 5721 34697 5733 34731
rect 5767 34728 5779 34731
rect 6178 34728 6184 34740
rect 5767 34700 6184 34728
rect 5767 34697 5779 34700
rect 5721 34691 5779 34697
rect 6178 34688 6184 34700
rect 6236 34688 6242 34740
rect 7466 34728 7472 34740
rect 7427 34700 7472 34728
rect 7466 34688 7472 34700
rect 7524 34728 7530 34740
rect 8202 34728 8208 34740
rect 7524 34700 8208 34728
rect 7524 34688 7530 34700
rect 8202 34688 8208 34700
rect 8260 34688 8266 34740
rect 13630 34728 13636 34740
rect 13591 34700 13636 34728
rect 13630 34688 13636 34700
rect 13688 34688 13694 34740
rect 198 34620 204 34672
rect 256 34660 262 34672
rect 1302 34660 1308 34672
rect 256 34632 1308 34660
rect 256 34620 262 34632
rect 1302 34620 1308 34632
rect 1360 34620 1366 34672
rect 1394 34620 1400 34672
rect 1452 34660 1458 34672
rect 2685 34663 2743 34669
rect 2685 34660 2697 34663
rect 1452 34632 2697 34660
rect 1452 34620 1458 34632
rect 2685 34629 2697 34632
rect 2731 34629 2743 34663
rect 9217 34663 9275 34669
rect 9217 34660 9229 34663
rect 2685 34623 2743 34629
rect 9140 34632 9229 34660
rect 2409 34595 2467 34601
rect 2409 34561 2421 34595
rect 2455 34592 2467 34595
rect 3050 34592 3056 34604
rect 2455 34564 3056 34592
rect 2455 34561 2467 34564
rect 2409 34555 2467 34561
rect 3050 34552 3056 34564
rect 3108 34552 3114 34604
rect 3145 34595 3203 34601
rect 3145 34561 3157 34595
rect 3191 34592 3203 34595
rect 3326 34592 3332 34604
rect 3191 34564 3332 34592
rect 3191 34561 3203 34564
rect 3145 34555 3203 34561
rect 1397 34527 1455 34533
rect 1397 34493 1409 34527
rect 1443 34524 1455 34527
rect 2038 34524 2044 34536
rect 1443 34496 2044 34524
rect 1443 34493 1455 34496
rect 1397 34487 1455 34493
rect 2038 34484 2044 34496
rect 2096 34484 2102 34536
rect 2501 34527 2559 34533
rect 2501 34493 2513 34527
rect 2547 34524 2559 34527
rect 3160 34524 3188 34555
rect 3326 34552 3332 34564
rect 3384 34552 3390 34604
rect 2547 34496 3188 34524
rect 2547 34493 2559 34496
rect 2501 34487 2559 34493
rect 3234 34484 3240 34536
rect 3292 34524 3298 34536
rect 3421 34527 3479 34533
rect 3421 34524 3433 34527
rect 3292 34496 3433 34524
rect 3292 34484 3298 34496
rect 3421 34493 3433 34496
rect 3467 34524 3479 34527
rect 3605 34527 3663 34533
rect 3605 34524 3617 34527
rect 3467 34496 3617 34524
rect 3467 34493 3479 34496
rect 3421 34487 3479 34493
rect 3605 34493 3617 34496
rect 3651 34493 3663 34527
rect 3605 34487 3663 34493
rect 4798 34484 4804 34536
rect 4856 34524 4862 34536
rect 5166 34524 5172 34536
rect 4856 34496 5172 34524
rect 4856 34484 4862 34496
rect 5166 34484 5172 34496
rect 5224 34484 5230 34536
rect 5537 34527 5595 34533
rect 5537 34493 5549 34527
rect 5583 34524 5595 34527
rect 5718 34524 5724 34536
rect 5583 34496 5724 34524
rect 5583 34493 5595 34496
rect 5537 34487 5595 34493
rect 5718 34484 5724 34496
rect 5776 34524 5782 34536
rect 6089 34527 6147 34533
rect 6089 34524 6101 34527
rect 5776 34496 6101 34524
rect 5776 34484 5782 34496
rect 6089 34493 6101 34496
rect 6135 34493 6147 34527
rect 6089 34487 6147 34493
rect 6549 34527 6607 34533
rect 6549 34493 6561 34527
rect 6595 34524 6607 34527
rect 6822 34524 6828 34536
rect 6595 34496 6828 34524
rect 6595 34493 6607 34496
rect 6549 34487 6607 34493
rect 6822 34484 6828 34496
rect 6880 34484 6886 34536
rect 7193 34527 7251 34533
rect 7193 34493 7205 34527
rect 7239 34524 7251 34527
rect 7834 34524 7840 34536
rect 7239 34496 7840 34524
rect 7239 34493 7251 34496
rect 7193 34487 7251 34493
rect 7834 34484 7840 34496
rect 7892 34484 7898 34536
rect 8110 34533 8116 34536
rect 8104 34524 8116 34533
rect 8071 34496 8116 34524
rect 8104 34487 8116 34496
rect 8110 34484 8116 34487
rect 8168 34484 8174 34536
rect 9140 34524 9168 34632
rect 9217 34629 9229 34632
rect 9263 34660 9275 34663
rect 9861 34663 9919 34669
rect 9861 34660 9873 34663
rect 9263 34632 9873 34660
rect 9263 34629 9275 34632
rect 9217 34623 9275 34629
rect 9861 34629 9873 34632
rect 9907 34629 9919 34663
rect 9861 34623 9919 34629
rect 9876 34592 9904 34623
rect 11054 34620 11060 34672
rect 11112 34660 11118 34672
rect 11425 34663 11483 34669
rect 11425 34660 11437 34663
rect 11112 34632 11437 34660
rect 11112 34620 11118 34632
rect 11425 34629 11437 34632
rect 11471 34629 11483 34663
rect 11425 34623 11483 34629
rect 9876 34564 10180 34592
rect 10042 34524 10048 34536
rect 8220 34496 9168 34524
rect 10003 34496 10048 34524
rect 8018 34416 8024 34468
rect 8076 34456 8082 34468
rect 8220 34456 8248 34496
rect 10042 34484 10048 34496
rect 10100 34484 10106 34536
rect 10152 34524 10180 34564
rect 10301 34527 10359 34533
rect 10301 34524 10313 34527
rect 10152 34496 10313 34524
rect 10301 34493 10313 34496
rect 10347 34493 10359 34527
rect 13446 34524 13452 34536
rect 13407 34496 13452 34524
rect 10301 34487 10359 34493
rect 13446 34484 13452 34496
rect 13504 34524 13510 34536
rect 14001 34527 14059 34533
rect 14001 34524 14013 34527
rect 13504 34496 14013 34524
rect 13504 34484 13510 34496
rect 14001 34493 14013 34496
rect 14047 34493 14059 34527
rect 14001 34487 14059 34493
rect 8076 34428 8248 34456
rect 8076 34416 8082 34428
rect 11793 34391 11851 34397
rect 11793 34357 11805 34391
rect 11839 34388 11851 34391
rect 12066 34388 12072 34400
rect 11839 34360 12072 34388
rect 11839 34357 11851 34360
rect 11793 34351 11851 34357
rect 12066 34348 12072 34360
rect 12124 34348 12130 34400
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 934 34144 940 34196
rect 992 34184 998 34196
rect 1581 34187 1639 34193
rect 1581 34184 1593 34187
rect 992 34156 1593 34184
rect 992 34144 998 34156
rect 1581 34153 1593 34156
rect 1627 34153 1639 34187
rect 1581 34147 1639 34153
rect 1762 34144 1768 34196
rect 1820 34184 1826 34196
rect 2685 34187 2743 34193
rect 2685 34184 2697 34187
rect 1820 34156 2697 34184
rect 1820 34144 1826 34156
rect 2685 34153 2697 34156
rect 2731 34153 2743 34187
rect 2685 34147 2743 34153
rect 4154 34144 4160 34196
rect 4212 34184 4218 34196
rect 4341 34187 4399 34193
rect 4341 34184 4353 34187
rect 4212 34156 4353 34184
rect 4212 34144 4218 34156
rect 4341 34153 4353 34156
rect 4387 34153 4399 34187
rect 4341 34147 4399 34153
rect 5534 34144 5540 34196
rect 5592 34184 5598 34196
rect 5997 34187 6055 34193
rect 5997 34184 6009 34187
rect 5592 34156 6009 34184
rect 5592 34144 5598 34156
rect 5997 34153 6009 34156
rect 6043 34153 6055 34187
rect 7742 34184 7748 34196
rect 7703 34156 7748 34184
rect 5997 34147 6055 34153
rect 7742 34144 7748 34156
rect 7800 34144 7806 34196
rect 10042 34184 10048 34196
rect 9784 34156 10048 34184
rect 1397 34051 1455 34057
rect 1397 34017 1409 34051
rect 1443 34048 1455 34051
rect 2406 34048 2412 34060
rect 1443 34020 2412 34048
rect 1443 34017 1455 34020
rect 1397 34011 1455 34017
rect 2406 34008 2412 34020
rect 2464 34008 2470 34060
rect 2501 34051 2559 34057
rect 2501 34017 2513 34051
rect 2547 34048 2559 34051
rect 3142 34048 3148 34060
rect 2547 34020 3148 34048
rect 2547 34017 2559 34020
rect 2501 34011 2559 34017
rect 3142 34008 3148 34020
rect 3200 34008 3206 34060
rect 4157 34051 4215 34057
rect 4157 34017 4169 34051
rect 4203 34048 4215 34051
rect 4246 34048 4252 34060
rect 4203 34020 4252 34048
rect 4203 34017 4215 34020
rect 4157 34011 4215 34017
rect 4246 34008 4252 34020
rect 4304 34008 4310 34060
rect 5813 34051 5871 34057
rect 5813 34017 5825 34051
rect 5859 34048 5871 34051
rect 6086 34048 6092 34060
rect 5859 34020 6092 34048
rect 5859 34017 5871 34020
rect 5813 34011 5871 34017
rect 6086 34008 6092 34020
rect 6144 34008 6150 34060
rect 7561 34051 7619 34057
rect 7561 34017 7573 34051
rect 7607 34048 7619 34051
rect 7834 34048 7840 34060
rect 7607 34020 7840 34048
rect 7607 34017 7619 34020
rect 7561 34011 7619 34017
rect 7834 34008 7840 34020
rect 7892 34008 7898 34060
rect 9674 34008 9680 34060
rect 9732 34048 9738 34060
rect 9784 34057 9812 34156
rect 10042 34144 10048 34156
rect 10100 34144 10106 34196
rect 11146 34184 11152 34196
rect 11059 34156 11152 34184
rect 11146 34144 11152 34156
rect 11204 34144 11210 34196
rect 11238 34144 11244 34196
rect 11296 34184 11302 34196
rect 12437 34187 12495 34193
rect 12437 34184 12449 34187
rect 11296 34156 12449 34184
rect 11296 34144 11302 34156
rect 12437 34153 12449 34156
rect 12483 34153 12495 34187
rect 12437 34147 12495 34153
rect 10060 34116 10088 34144
rect 11164 34116 11192 34144
rect 12066 34116 12072 34128
rect 10060 34088 10180 34116
rect 11164 34088 12072 34116
rect 10042 34057 10048 34060
rect 9769 34051 9827 34057
rect 9769 34048 9781 34051
rect 9732 34020 9781 34048
rect 9732 34008 9738 34020
rect 9769 34017 9781 34020
rect 9815 34017 9827 34051
rect 10036 34048 10048 34057
rect 10003 34020 10048 34048
rect 9769 34011 9827 34017
rect 10036 34011 10048 34020
rect 10042 34008 10048 34011
rect 10100 34008 10106 34060
rect 10152 34048 10180 34088
rect 12066 34076 12072 34088
rect 12124 34076 12130 34128
rect 10152 34020 10824 34048
rect 10796 33980 10824 34020
rect 11146 34008 11152 34060
rect 11204 34048 11210 34060
rect 12345 34051 12403 34057
rect 12345 34048 12357 34051
rect 11204 34020 12357 34048
rect 11204 34008 11210 34020
rect 12345 34017 12357 34020
rect 12391 34048 12403 34051
rect 13446 34048 13452 34060
rect 12391 34020 13452 34048
rect 12391 34017 12403 34020
rect 12345 34011 12403 34017
rect 13446 34008 13452 34020
rect 13504 34008 13510 34060
rect 11425 33983 11483 33989
rect 11425 33980 11437 33983
rect 10796 33952 11437 33980
rect 11425 33949 11437 33952
rect 11471 33949 11483 33983
rect 12526 33980 12532 33992
rect 12487 33952 12532 33980
rect 11425 33943 11483 33949
rect 12526 33940 12532 33952
rect 12584 33940 12590 33992
rect 10778 33872 10784 33924
rect 10836 33912 10842 33924
rect 11977 33915 12035 33921
rect 11977 33912 11989 33915
rect 10836 33884 11989 33912
rect 10836 33872 10842 33884
rect 11977 33881 11989 33884
rect 12023 33881 12035 33915
rect 11977 33875 12035 33881
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 1394 33600 1400 33652
rect 1452 33640 1458 33652
rect 1581 33643 1639 33649
rect 1581 33640 1593 33643
rect 1452 33612 1593 33640
rect 1452 33600 1458 33612
rect 1581 33609 1593 33612
rect 1627 33609 1639 33643
rect 1581 33603 1639 33609
rect 2130 33600 2136 33652
rect 2188 33640 2194 33652
rect 2685 33643 2743 33649
rect 2685 33640 2697 33643
rect 2188 33612 2697 33640
rect 2188 33600 2194 33612
rect 2685 33609 2697 33612
rect 2731 33609 2743 33643
rect 7374 33640 7380 33652
rect 7335 33612 7380 33640
rect 2685 33603 2743 33609
rect 7374 33600 7380 33612
rect 7432 33600 7438 33652
rect 7834 33600 7840 33652
rect 7892 33640 7898 33652
rect 8113 33643 8171 33649
rect 8113 33640 8125 33643
rect 7892 33612 8125 33640
rect 7892 33600 7898 33612
rect 8113 33609 8125 33612
rect 8159 33609 8171 33643
rect 8113 33603 8171 33609
rect 8570 33600 8576 33652
rect 8628 33640 8634 33652
rect 8941 33643 8999 33649
rect 8941 33640 8953 33643
rect 8628 33612 8953 33640
rect 8628 33600 8634 33612
rect 8941 33609 8953 33612
rect 8987 33640 8999 33643
rect 9217 33643 9275 33649
rect 9217 33640 9229 33643
rect 8987 33612 9229 33640
rect 8987 33609 8999 33612
rect 8941 33603 8999 33609
rect 9217 33609 9229 33612
rect 9263 33609 9275 33643
rect 9217 33603 9275 33609
rect 9306 33600 9312 33652
rect 9364 33640 9370 33652
rect 10597 33643 10655 33649
rect 9364 33612 9409 33640
rect 9364 33600 9370 33612
rect 10597 33609 10609 33643
rect 10643 33640 10655 33643
rect 10962 33640 10968 33652
rect 10643 33612 10968 33640
rect 10643 33609 10655 33612
rect 10597 33603 10655 33609
rect 8665 33507 8723 33513
rect 8665 33473 8677 33507
rect 8711 33504 8723 33507
rect 10042 33504 10048 33516
rect 8711 33476 10048 33504
rect 8711 33473 8723 33476
rect 8665 33467 8723 33473
rect 10042 33464 10048 33476
rect 10100 33504 10106 33516
rect 10137 33507 10195 33513
rect 10137 33504 10149 33507
rect 10100 33476 10149 33504
rect 10100 33464 10106 33476
rect 10137 33473 10149 33476
rect 10183 33504 10195 33507
rect 10612 33504 10640 33603
rect 10962 33600 10968 33612
rect 11020 33600 11026 33652
rect 11149 33643 11207 33649
rect 11149 33609 11161 33643
rect 11195 33640 11207 33643
rect 11238 33640 11244 33652
rect 11195 33612 11244 33640
rect 11195 33609 11207 33612
rect 11149 33603 11207 33609
rect 11238 33600 11244 33612
rect 11296 33600 11302 33652
rect 13446 33640 13452 33652
rect 13407 33612 13452 33640
rect 13446 33600 13452 33612
rect 13504 33600 13510 33652
rect 10183 33476 10640 33504
rect 10183 33473 10195 33476
rect 10137 33467 10195 33473
rect 12066 33464 12072 33516
rect 12124 33504 12130 33516
rect 12989 33507 13047 33513
rect 12989 33504 13001 33507
rect 12124 33476 13001 33504
rect 12124 33464 12130 33476
rect 12989 33473 13001 33476
rect 13035 33473 13047 33507
rect 12989 33467 13047 33473
rect 1397 33439 1455 33445
rect 1397 33405 1409 33439
rect 1443 33436 1455 33439
rect 2501 33439 2559 33445
rect 1443 33408 2084 33436
rect 1443 33405 1455 33408
rect 1397 33399 1455 33405
rect 2056 33312 2084 33408
rect 2501 33405 2513 33439
rect 2547 33436 2559 33439
rect 2682 33436 2688 33448
rect 2547 33408 2688 33436
rect 2547 33405 2559 33408
rect 2501 33399 2559 33405
rect 2682 33396 2688 33408
rect 2740 33396 2746 33448
rect 7193 33439 7251 33445
rect 7193 33405 7205 33439
rect 7239 33436 7251 33439
rect 7742 33436 7748 33448
rect 7239 33408 7748 33436
rect 7239 33405 7251 33408
rect 7193 33399 7251 33405
rect 7742 33396 7748 33408
rect 7800 33396 7806 33448
rect 9217 33439 9275 33445
rect 9217 33405 9229 33439
rect 9263 33436 9275 33439
rect 9861 33439 9919 33445
rect 9861 33436 9873 33439
rect 9263 33408 9873 33436
rect 9263 33405 9275 33408
rect 9217 33399 9275 33405
rect 9861 33405 9873 33408
rect 9907 33405 9919 33439
rect 12342 33436 12348 33448
rect 9861 33399 9919 33405
rect 11440 33408 12348 33436
rect 3142 33368 3148 33380
rect 3055 33340 3148 33368
rect 3142 33328 3148 33340
rect 3200 33368 3206 33380
rect 4706 33368 4712 33380
rect 3200 33340 4712 33368
rect 3200 33328 3206 33340
rect 4706 33328 4712 33340
rect 4764 33328 4770 33380
rect 9306 33328 9312 33380
rect 9364 33368 9370 33380
rect 9953 33371 10011 33377
rect 9953 33368 9965 33371
rect 9364 33340 9965 33368
rect 9364 33328 9370 33340
rect 9953 33337 9965 33340
rect 9999 33337 10011 33371
rect 9953 33331 10011 33337
rect 11440 33312 11468 33408
rect 12342 33396 12348 33408
rect 12400 33396 12406 33448
rect 12158 33368 12164 33380
rect 12119 33340 12164 33368
rect 12158 33328 12164 33340
rect 12216 33368 12222 33380
rect 12894 33368 12900 33380
rect 12216 33340 12900 33368
rect 12216 33328 12222 33340
rect 12894 33328 12900 33340
rect 12952 33328 12958 33380
rect 2038 33300 2044 33312
rect 1999 33272 2044 33300
rect 2038 33260 2044 33272
rect 2096 33260 2102 33312
rect 2406 33300 2412 33312
rect 2367 33272 2412 33300
rect 2406 33260 2412 33272
rect 2464 33260 2470 33312
rect 4246 33300 4252 33312
rect 4207 33272 4252 33300
rect 4246 33260 4252 33272
rect 4304 33260 4310 33312
rect 5166 33300 5172 33312
rect 5127 33272 5172 33300
rect 5166 33260 5172 33272
rect 5224 33260 5230 33312
rect 5905 33303 5963 33309
rect 5905 33269 5917 33303
rect 5951 33300 5963 33303
rect 6086 33300 6092 33312
rect 5951 33272 6092 33300
rect 5951 33269 5963 33272
rect 5905 33263 5963 33269
rect 6086 33260 6092 33272
rect 6144 33260 6150 33312
rect 9490 33300 9496 33312
rect 9451 33272 9496 33300
rect 9490 33260 9496 33272
rect 9548 33260 9554 33312
rect 11422 33300 11428 33312
rect 11383 33272 11428 33300
rect 11422 33260 11428 33272
rect 11480 33260 11486 33312
rect 11885 33303 11943 33309
rect 11885 33269 11897 33303
rect 11931 33300 11943 33303
rect 12066 33300 12072 33312
rect 11931 33272 12072 33300
rect 11931 33269 11943 33272
rect 11885 33263 11943 33269
rect 12066 33260 12072 33272
rect 12124 33260 12130 33312
rect 12434 33260 12440 33312
rect 12492 33300 12498 33312
rect 12802 33300 12808 33312
rect 12492 33272 12537 33300
rect 12763 33272 12808 33300
rect 12492 33260 12498 33272
rect 12802 33260 12808 33272
rect 12860 33260 12866 33312
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 5166 33056 5172 33108
rect 5224 33096 5230 33108
rect 5445 33099 5503 33105
rect 5445 33096 5457 33099
rect 5224 33068 5457 33096
rect 5224 33056 5230 33068
rect 5445 33065 5457 33068
rect 5491 33065 5503 33099
rect 5445 33059 5503 33065
rect 9490 33056 9496 33108
rect 9548 33096 9554 33108
rect 10413 33099 10471 33105
rect 10413 33096 10425 33099
rect 9548 33068 10425 33096
rect 9548 33056 9554 33068
rect 10413 33065 10425 33068
rect 10459 33065 10471 33099
rect 10413 33059 10471 33065
rect 10870 33056 10876 33108
rect 10928 33096 10934 33108
rect 11885 33099 11943 33105
rect 11885 33096 11897 33099
rect 10928 33068 11897 33096
rect 10928 33056 10934 33068
rect 11624 33040 11652 33068
rect 11885 33065 11897 33068
rect 11931 33065 11943 33099
rect 11885 33059 11943 33065
rect 12621 33099 12679 33105
rect 12621 33065 12633 33099
rect 12667 33096 12679 33099
rect 12802 33096 12808 33108
rect 12667 33068 12808 33096
rect 12667 33065 12679 33068
rect 12621 33059 12679 33065
rect 12802 33056 12808 33068
rect 12860 33056 12866 33108
rect 1486 32988 1492 33040
rect 1544 33028 1550 33040
rect 1673 33031 1731 33037
rect 1673 33028 1685 33031
rect 1544 33000 1685 33028
rect 1544 32988 1550 33000
rect 1673 32997 1685 33000
rect 1719 32997 1731 33031
rect 1673 32991 1731 32997
rect 11606 32988 11612 33040
rect 11664 32988 11670 33040
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32960 1455 32963
rect 1762 32960 1768 32972
rect 1443 32932 1768 32960
rect 1443 32929 1455 32932
rect 1397 32923 1455 32929
rect 1762 32920 1768 32932
rect 1820 32920 1826 32972
rect 6914 32969 6920 32972
rect 6908 32960 6920 32969
rect 6875 32932 6920 32960
rect 6908 32923 6920 32932
rect 6914 32920 6920 32923
rect 6972 32920 6978 32972
rect 9493 32963 9551 32969
rect 9493 32929 9505 32963
rect 9539 32960 9551 32963
rect 9674 32960 9680 32972
rect 9539 32932 9680 32960
rect 9539 32929 9551 32932
rect 9493 32923 9551 32929
rect 9674 32920 9680 32932
rect 9732 32920 9738 32972
rect 10042 32920 10048 32972
rect 10100 32960 10106 32972
rect 10321 32963 10379 32969
rect 10321 32960 10333 32963
rect 10100 32932 10333 32960
rect 10100 32920 10106 32932
rect 10321 32929 10333 32932
rect 10367 32929 10379 32963
rect 10321 32923 10379 32929
rect 5534 32892 5540 32904
rect 5495 32864 5540 32892
rect 5534 32852 5540 32864
rect 5592 32852 5598 32904
rect 5721 32895 5779 32901
rect 5721 32861 5733 32895
rect 5767 32892 5779 32895
rect 6638 32892 6644 32904
rect 5767 32864 6408 32892
rect 6599 32864 6644 32892
rect 5767 32861 5779 32864
rect 5721 32855 5779 32861
rect 4985 32827 5043 32833
rect 4985 32793 4997 32827
rect 5031 32824 5043 32827
rect 5736 32824 5764 32855
rect 5031 32796 5764 32824
rect 5031 32793 5043 32796
rect 4985 32787 5043 32793
rect 2593 32759 2651 32765
rect 2593 32725 2605 32759
rect 2639 32756 2651 32759
rect 2682 32756 2688 32768
rect 2639 32728 2688 32756
rect 2639 32725 2651 32728
rect 2593 32719 2651 32725
rect 2682 32716 2688 32728
rect 2740 32716 2746 32768
rect 5077 32759 5135 32765
rect 5077 32725 5089 32759
rect 5123 32756 5135 32759
rect 5442 32756 5448 32768
rect 5123 32728 5448 32756
rect 5123 32725 5135 32728
rect 5077 32719 5135 32725
rect 5442 32716 5448 32728
rect 5500 32716 5506 32768
rect 6380 32756 6408 32864
rect 6638 32852 6644 32864
rect 6696 32852 6702 32904
rect 10597 32895 10655 32901
rect 10597 32861 10609 32895
rect 10643 32892 10655 32895
rect 11054 32892 11060 32904
rect 10643 32864 11060 32892
rect 10643 32861 10655 32864
rect 10597 32855 10655 32861
rect 11054 32852 11060 32864
rect 11112 32892 11118 32904
rect 11974 32892 11980 32904
rect 11112 32864 11836 32892
rect 11935 32864 11980 32892
rect 11112 32852 11118 32864
rect 9953 32827 10011 32833
rect 9953 32793 9965 32827
rect 9999 32824 10011 32827
rect 11238 32824 11244 32836
rect 9999 32796 11244 32824
rect 9999 32793 10011 32796
rect 9953 32787 10011 32793
rect 11238 32784 11244 32796
rect 11296 32784 11302 32836
rect 11808 32824 11836 32864
rect 11974 32852 11980 32864
rect 12032 32852 12038 32904
rect 12066 32852 12072 32904
rect 12124 32892 12130 32904
rect 12124 32864 12217 32892
rect 12124 32852 12130 32864
rect 12084 32824 12112 32852
rect 11808 32796 12112 32824
rect 7006 32756 7012 32768
rect 6380 32728 7012 32756
rect 7006 32716 7012 32728
rect 7064 32756 7070 32768
rect 8021 32759 8079 32765
rect 8021 32756 8033 32759
rect 7064 32728 8033 32756
rect 7064 32716 7070 32728
rect 8021 32725 8033 32728
rect 8067 32725 8079 32759
rect 8021 32719 8079 32725
rect 8941 32759 8999 32765
rect 8941 32725 8953 32759
rect 8987 32756 8999 32759
rect 9306 32756 9312 32768
rect 8987 32728 9312 32756
rect 8987 32725 8999 32728
rect 8941 32719 8999 32725
rect 9306 32716 9312 32728
rect 9364 32716 9370 32768
rect 11514 32756 11520 32768
rect 11475 32728 11520 32756
rect 11514 32716 11520 32728
rect 11572 32716 11578 32768
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 4982 32552 4988 32564
rect 4943 32524 4988 32552
rect 4982 32512 4988 32524
rect 5040 32512 5046 32564
rect 5166 32552 5172 32564
rect 5127 32524 5172 32552
rect 5166 32512 5172 32524
rect 5224 32512 5230 32564
rect 6178 32552 6184 32564
rect 5460 32524 6184 32552
rect 5000 32416 5028 32512
rect 5460 32416 5488 32524
rect 6178 32512 6184 32524
rect 6236 32512 6242 32564
rect 6546 32552 6552 32564
rect 6507 32524 6552 32552
rect 6546 32512 6552 32524
rect 6604 32512 6610 32564
rect 8294 32512 8300 32564
rect 8352 32552 8358 32564
rect 8573 32555 8631 32561
rect 8573 32552 8585 32555
rect 8352 32524 8585 32552
rect 8352 32512 8358 32524
rect 8573 32521 8585 32524
rect 8619 32552 8631 32555
rect 8665 32555 8723 32561
rect 8665 32552 8677 32555
rect 8619 32524 8677 32552
rect 8619 32521 8631 32524
rect 8573 32515 8631 32521
rect 8665 32521 8677 32524
rect 8711 32521 8723 32555
rect 10042 32552 10048 32564
rect 10003 32524 10048 32552
rect 8665 32515 8723 32521
rect 10042 32512 10048 32524
rect 10100 32512 10106 32564
rect 10318 32552 10324 32564
rect 10279 32524 10324 32552
rect 10318 32512 10324 32524
rect 10376 32512 10382 32564
rect 10505 32555 10563 32561
rect 10505 32521 10517 32555
rect 10551 32552 10563 32555
rect 10962 32552 10968 32564
rect 10551 32524 10968 32552
rect 10551 32521 10563 32524
rect 10505 32515 10563 32521
rect 10962 32512 10968 32524
rect 11020 32512 11026 32564
rect 11606 32552 11612 32564
rect 11567 32524 11612 32552
rect 11606 32512 11612 32524
rect 11664 32512 11670 32564
rect 11974 32552 11980 32564
rect 11935 32524 11980 32552
rect 11974 32512 11980 32524
rect 12032 32512 12038 32564
rect 5534 32444 5540 32496
rect 5592 32484 5598 32496
rect 6825 32487 6883 32493
rect 6825 32484 6837 32487
rect 5592 32456 6837 32484
rect 5592 32444 5598 32456
rect 6825 32453 6837 32456
rect 6871 32453 6883 32487
rect 6825 32447 6883 32453
rect 6914 32444 6920 32496
rect 6972 32444 6978 32496
rect 5629 32419 5687 32425
rect 5629 32416 5641 32419
rect 5000 32388 5641 32416
rect 5629 32385 5641 32388
rect 5675 32385 5687 32419
rect 5629 32379 5687 32385
rect 5721 32419 5779 32425
rect 5721 32385 5733 32419
rect 5767 32385 5779 32419
rect 6932 32416 6960 32444
rect 7377 32419 7435 32425
rect 7377 32416 7389 32419
rect 5721 32379 5779 32385
rect 6196 32388 7389 32416
rect 4341 32351 4399 32357
rect 4341 32317 4353 32351
rect 4387 32348 4399 32351
rect 5736 32348 5764 32379
rect 5902 32348 5908 32360
rect 4387 32320 5908 32348
rect 4387 32317 4399 32320
rect 4341 32311 4399 32317
rect 5902 32308 5908 32320
rect 5960 32348 5966 32360
rect 6196 32357 6224 32388
rect 7377 32385 7389 32388
rect 7423 32385 7435 32419
rect 7377 32379 7435 32385
rect 8389 32419 8447 32425
rect 8389 32385 8401 32419
rect 8435 32416 8447 32419
rect 8570 32416 8576 32428
rect 8435 32388 8576 32416
rect 8435 32385 8447 32388
rect 8389 32379 8447 32385
rect 8570 32376 8576 32388
rect 8628 32416 8634 32428
rect 9401 32419 9459 32425
rect 9401 32416 9413 32419
rect 8628 32388 9413 32416
rect 8628 32376 8634 32388
rect 9401 32385 9413 32388
rect 9447 32385 9459 32419
rect 11054 32416 11060 32428
rect 11015 32388 11060 32416
rect 9401 32379 9459 32385
rect 11054 32376 11060 32388
rect 11112 32376 11118 32428
rect 12437 32419 12495 32425
rect 12437 32385 12449 32419
rect 12483 32416 12495 32419
rect 12802 32416 12808 32428
rect 12483 32388 12808 32416
rect 12483 32385 12495 32388
rect 12437 32379 12495 32385
rect 12802 32376 12808 32388
rect 12860 32376 12866 32428
rect 6181 32351 6239 32357
rect 6181 32348 6193 32351
rect 5960 32320 6193 32348
rect 5960 32308 5966 32320
rect 6181 32317 6193 32320
rect 6227 32317 6239 32351
rect 6181 32311 6239 32317
rect 6914 32308 6920 32360
rect 6972 32348 6978 32360
rect 7193 32351 7251 32357
rect 7193 32348 7205 32351
rect 6972 32320 7205 32348
rect 6972 32308 6978 32320
rect 7193 32317 7205 32320
rect 7239 32348 7251 32351
rect 7926 32348 7932 32360
rect 7239 32320 7932 32348
rect 7239 32317 7251 32320
rect 7193 32311 7251 32317
rect 7926 32308 7932 32320
rect 7984 32308 7990 32360
rect 9306 32348 9312 32360
rect 9267 32320 9312 32348
rect 9306 32308 9312 32320
rect 9364 32308 9370 32360
rect 10318 32308 10324 32360
rect 10376 32348 10382 32360
rect 10873 32351 10931 32357
rect 10873 32348 10885 32351
rect 10376 32320 10885 32348
rect 10376 32308 10382 32320
rect 10873 32317 10885 32320
rect 10919 32317 10931 32351
rect 10873 32311 10931 32317
rect 6546 32240 6552 32292
rect 6604 32280 6610 32292
rect 6730 32280 6736 32292
rect 6604 32252 6736 32280
rect 6604 32240 6610 32252
rect 6730 32240 6736 32252
rect 6788 32280 6794 32292
rect 7285 32283 7343 32289
rect 7285 32280 7297 32283
rect 6788 32252 7297 32280
rect 6788 32240 6794 32252
rect 7285 32249 7297 32252
rect 7331 32249 7343 32283
rect 7285 32243 7343 32249
rect 8573 32283 8631 32289
rect 8573 32249 8585 32283
rect 8619 32280 8631 32283
rect 8662 32280 8668 32292
rect 8619 32252 8668 32280
rect 8619 32249 8631 32252
rect 8573 32243 8631 32249
rect 8662 32240 8668 32252
rect 8720 32280 8726 32292
rect 9217 32283 9275 32289
rect 9217 32280 9229 32283
rect 8720 32252 9229 32280
rect 8720 32240 8726 32252
rect 9217 32249 9229 32252
rect 9263 32249 9275 32283
rect 9217 32243 9275 32249
rect 1673 32215 1731 32221
rect 1673 32181 1685 32215
rect 1719 32212 1731 32215
rect 1762 32212 1768 32224
rect 1719 32184 1768 32212
rect 1719 32181 1731 32184
rect 1673 32175 1731 32181
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 4709 32215 4767 32221
rect 4709 32181 4721 32215
rect 4755 32212 4767 32215
rect 5537 32215 5595 32221
rect 5537 32212 5549 32215
rect 4755 32184 5549 32212
rect 4755 32181 4767 32184
rect 4709 32175 4767 32181
rect 5537 32181 5549 32184
rect 5583 32212 5595 32215
rect 5626 32212 5632 32224
rect 5583 32184 5632 32212
rect 5583 32181 5595 32184
rect 5537 32175 5595 32181
rect 5626 32172 5632 32184
rect 5684 32172 5690 32224
rect 7374 32172 7380 32224
rect 7432 32212 7438 32224
rect 7837 32215 7895 32221
rect 7837 32212 7849 32215
rect 7432 32184 7849 32212
rect 7432 32172 7438 32184
rect 7837 32181 7849 32184
rect 7883 32181 7895 32215
rect 8846 32212 8852 32224
rect 8807 32184 8852 32212
rect 7837 32175 7895 32181
rect 8846 32172 8852 32184
rect 8904 32172 8910 32224
rect 10962 32212 10968 32224
rect 10923 32184 10968 32212
rect 10962 32172 10968 32184
rect 11020 32172 11026 32224
rect 11974 32172 11980 32224
rect 12032 32212 12038 32224
rect 12618 32212 12624 32224
rect 12032 32184 12624 32212
rect 12032 32172 12038 32184
rect 12618 32172 12624 32184
rect 12676 32172 12682 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 4801 32011 4859 32017
rect 4801 31977 4813 32011
rect 4847 32008 4859 32011
rect 5534 32008 5540 32020
rect 4847 31980 5540 32008
rect 4847 31977 4859 31980
rect 4801 31971 4859 31977
rect 5534 31968 5540 31980
rect 5592 31968 5598 32020
rect 5902 31968 5908 32020
rect 5960 32008 5966 32020
rect 6273 32011 6331 32017
rect 6273 32008 6285 32011
rect 5960 31980 6285 32008
rect 5960 31968 5966 31980
rect 6273 31977 6285 31980
rect 6319 31977 6331 32011
rect 6914 32008 6920 32020
rect 6875 31980 6920 32008
rect 6273 31971 6331 31977
rect 1670 31940 1676 31952
rect 1631 31912 1676 31940
rect 1670 31900 1676 31912
rect 1728 31900 1734 31952
rect 5626 31940 5632 31952
rect 4908 31912 5632 31940
rect 4908 31881 4936 31912
rect 5626 31900 5632 31912
rect 5684 31900 5690 31952
rect 6288 31940 6316 31971
rect 6914 31968 6920 31980
rect 6972 31968 6978 32020
rect 8294 31968 8300 32020
rect 8352 32008 8358 32020
rect 8757 32011 8815 32017
rect 8757 32008 8769 32011
rect 8352 31980 8769 32008
rect 8352 31968 8358 31980
rect 8757 31977 8769 31980
rect 8803 31977 8815 32011
rect 9490 32008 9496 32020
rect 9451 31980 9496 32008
rect 8757 31971 8815 31977
rect 9490 31968 9496 31980
rect 9548 31968 9554 32020
rect 10229 32011 10287 32017
rect 10229 31977 10241 32011
rect 10275 32008 10287 32011
rect 10873 32011 10931 32017
rect 10873 32008 10885 32011
rect 10275 31980 10885 32008
rect 10275 31977 10287 31980
rect 10229 31971 10287 31977
rect 10873 31977 10885 31980
rect 10919 32008 10931 32011
rect 11054 32008 11060 32020
rect 10919 31980 11060 32008
rect 10919 31977 10931 31980
rect 10873 31971 10931 31977
rect 11054 31968 11060 31980
rect 11112 31968 11118 32020
rect 11514 32008 11520 32020
rect 11475 31980 11520 32008
rect 11514 31968 11520 31980
rect 11572 31968 11578 32020
rect 7190 31940 7196 31952
rect 6288 31912 7196 31940
rect 7190 31900 7196 31912
rect 7248 31900 7254 31952
rect 7466 31900 7472 31952
rect 7524 31940 7530 31952
rect 7644 31943 7702 31949
rect 7644 31940 7656 31943
rect 7524 31912 7656 31940
rect 7524 31900 7530 31912
rect 7644 31909 7656 31912
rect 7690 31940 7702 31943
rect 8570 31940 8576 31952
rect 7690 31912 8576 31940
rect 7690 31909 7702 31912
rect 7644 31903 7702 31909
rect 8570 31900 8576 31912
rect 8628 31900 8634 31952
rect 9582 31900 9588 31952
rect 9640 31940 9646 31952
rect 10505 31943 10563 31949
rect 10505 31940 10517 31943
rect 9640 31912 10517 31940
rect 9640 31900 9646 31912
rect 10505 31909 10517 31912
rect 10551 31940 10563 31943
rect 10962 31940 10968 31952
rect 10551 31912 10968 31940
rect 10551 31909 10563 31912
rect 10505 31903 10563 31909
rect 10962 31900 10968 31912
rect 11020 31900 11026 31952
rect 11072 31940 11100 31968
rect 12069 31943 12127 31949
rect 12069 31940 12081 31943
rect 11072 31912 12081 31940
rect 12069 31909 12081 31912
rect 12115 31909 12127 31943
rect 12069 31903 12127 31909
rect 5166 31881 5172 31884
rect 1397 31875 1455 31881
rect 1397 31841 1409 31875
rect 1443 31872 1455 31875
rect 4893 31875 4951 31881
rect 4893 31872 4905 31875
rect 1443 31844 1716 31872
rect 1443 31841 1455 31844
rect 1397 31835 1455 31841
rect 1688 31816 1716 31844
rect 3804 31844 4905 31872
rect 1670 31764 1676 31816
rect 1728 31764 1734 31816
rect 3418 31628 3424 31680
rect 3476 31668 3482 31680
rect 3697 31671 3755 31677
rect 3697 31668 3709 31671
rect 3476 31640 3709 31668
rect 3476 31628 3482 31640
rect 3697 31637 3709 31640
rect 3743 31668 3755 31671
rect 3804 31668 3832 31844
rect 4893 31841 4905 31844
rect 4939 31841 4951 31875
rect 4893 31835 4951 31841
rect 5160 31835 5172 31881
rect 5224 31872 5230 31884
rect 5224 31844 5260 31872
rect 5166 31832 5172 31835
rect 5224 31832 5230 31844
rect 6546 31832 6552 31884
rect 6604 31872 6610 31884
rect 7374 31872 7380 31884
rect 6604 31844 7380 31872
rect 6604 31832 6610 31844
rect 7374 31832 7380 31844
rect 7432 31832 7438 31884
rect 11425 31875 11483 31881
rect 11425 31841 11437 31875
rect 11471 31872 11483 31875
rect 12342 31872 12348 31884
rect 11471 31844 12348 31872
rect 11471 31841 11483 31844
rect 11425 31835 11483 31841
rect 12342 31832 12348 31844
rect 12400 31832 12406 31884
rect 9677 31807 9735 31813
rect 9677 31773 9689 31807
rect 9723 31804 9735 31807
rect 9950 31804 9956 31816
rect 9723 31776 9956 31804
rect 9723 31773 9735 31776
rect 9677 31767 9735 31773
rect 9950 31764 9956 31776
rect 10008 31764 10014 31816
rect 11609 31807 11667 31813
rect 11609 31773 11621 31807
rect 11655 31804 11667 31807
rect 14918 31804 14924 31816
rect 11655 31776 11689 31804
rect 14752 31776 14924 31804
rect 11655 31773 11667 31776
rect 11609 31767 11667 31773
rect 11422 31696 11428 31748
rect 11480 31736 11486 31748
rect 11624 31736 11652 31767
rect 14752 31748 14780 31776
rect 14918 31764 14924 31776
rect 14976 31764 14982 31816
rect 11480 31708 11652 31736
rect 11480 31696 11486 31708
rect 14734 31696 14740 31748
rect 14792 31696 14798 31748
rect 3743 31640 3832 31668
rect 3743 31637 3755 31640
rect 3697 31631 3755 31637
rect 10502 31628 10508 31680
rect 10560 31668 10566 31680
rect 11057 31671 11115 31677
rect 11057 31668 11069 31671
rect 10560 31640 11069 31668
rect 10560 31628 10566 31640
rect 11057 31637 11069 31640
rect 11103 31637 11115 31671
rect 11057 31631 11115 31637
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 5626 31424 5632 31476
rect 5684 31464 5690 31476
rect 5813 31467 5871 31473
rect 5813 31464 5825 31467
rect 5684 31436 5825 31464
rect 5684 31424 5690 31436
rect 5813 31433 5825 31436
rect 5859 31464 5871 31467
rect 6546 31464 6552 31476
rect 5859 31436 6552 31464
rect 5859 31433 5871 31436
rect 5813 31427 5871 31433
rect 6546 31424 6552 31436
rect 6604 31424 6610 31476
rect 7193 31467 7251 31473
rect 7193 31433 7205 31467
rect 7239 31464 7251 31467
rect 7466 31464 7472 31476
rect 7239 31436 7472 31464
rect 7239 31433 7251 31436
rect 7193 31427 7251 31433
rect 7466 31424 7472 31436
rect 7524 31424 7530 31476
rect 11514 31464 11520 31476
rect 11475 31436 11520 31464
rect 11514 31424 11520 31436
rect 11572 31424 11578 31476
rect 11977 31467 12035 31473
rect 11977 31433 11989 31467
rect 12023 31464 12035 31467
rect 12342 31464 12348 31476
rect 12023 31436 12348 31464
rect 12023 31433 12035 31436
rect 11977 31427 12035 31433
rect 12342 31424 12348 31436
rect 12400 31424 12406 31476
rect 7561 31331 7619 31337
rect 7561 31297 7573 31331
rect 7607 31328 7619 31331
rect 8018 31328 8024 31340
rect 7607 31300 8024 31328
rect 7607 31297 7619 31300
rect 7561 31291 7619 31297
rect 8018 31288 8024 31300
rect 8076 31328 8082 31340
rect 8205 31331 8263 31337
rect 8205 31328 8217 31331
rect 8076 31300 8217 31328
rect 8076 31288 8082 31300
rect 8205 31297 8217 31300
rect 8251 31297 8263 31331
rect 8205 31291 8263 31297
rect 10045 31331 10103 31337
rect 10045 31297 10057 31331
rect 10091 31328 10103 31331
rect 10689 31331 10747 31337
rect 10689 31328 10701 31331
rect 10091 31300 10701 31328
rect 10091 31297 10103 31300
rect 10045 31291 10103 31297
rect 10689 31297 10701 31300
rect 10735 31328 10747 31331
rect 11514 31328 11520 31340
rect 10735 31300 11520 31328
rect 10735 31297 10747 31300
rect 10689 31291 10747 31297
rect 11514 31288 11520 31300
rect 11572 31288 11578 31340
rect 1670 31260 1676 31272
rect 1631 31232 1676 31260
rect 1670 31220 1676 31232
rect 1728 31220 1734 31272
rect 3418 31220 3424 31272
rect 3476 31260 3482 31272
rect 3697 31263 3755 31269
rect 3697 31260 3709 31263
rect 3476 31232 3709 31260
rect 3476 31220 3482 31232
rect 3697 31229 3709 31232
rect 3743 31229 3755 31263
rect 3697 31223 3755 31229
rect 9677 31263 9735 31269
rect 9677 31229 9689 31263
rect 9723 31260 9735 31263
rect 10502 31260 10508 31272
rect 9723 31232 10508 31260
rect 9723 31229 9735 31232
rect 9677 31223 9735 31229
rect 10502 31220 10508 31232
rect 10560 31220 10566 31272
rect 10597 31263 10655 31269
rect 10597 31229 10609 31263
rect 10643 31260 10655 31263
rect 10778 31260 10784 31272
rect 10643 31232 10784 31260
rect 10643 31229 10655 31232
rect 10597 31223 10655 31229
rect 10778 31220 10784 31232
rect 10836 31220 10842 31272
rect 3605 31195 3663 31201
rect 3605 31161 3617 31195
rect 3651 31192 3663 31195
rect 3964 31195 4022 31201
rect 3964 31192 3976 31195
rect 3651 31164 3976 31192
rect 3651 31161 3663 31164
rect 3605 31155 3663 31161
rect 3964 31161 3976 31164
rect 4010 31192 4022 31195
rect 4338 31192 4344 31204
rect 4010 31164 4344 31192
rect 4010 31161 4022 31164
rect 3964 31155 4022 31161
rect 4338 31152 4344 31164
rect 4396 31152 4402 31204
rect 8018 31192 8024 31204
rect 7931 31164 8024 31192
rect 8018 31152 8024 31164
rect 8076 31192 8082 31204
rect 8665 31195 8723 31201
rect 8665 31192 8677 31195
rect 8076 31164 8677 31192
rect 8076 31152 8082 31164
rect 8665 31161 8677 31164
rect 8711 31161 8723 31195
rect 8665 31155 8723 31161
rect 4154 31084 4160 31136
rect 4212 31124 4218 31136
rect 5077 31127 5135 31133
rect 5077 31124 5089 31127
rect 4212 31096 5089 31124
rect 4212 31084 4218 31096
rect 5077 31093 5089 31096
rect 5123 31124 5135 31127
rect 5166 31124 5172 31136
rect 5123 31096 5172 31124
rect 5123 31093 5135 31096
rect 5077 31087 5135 31093
rect 5166 31084 5172 31096
rect 5224 31124 5230 31136
rect 5353 31127 5411 31133
rect 5353 31124 5365 31127
rect 5224 31096 5365 31124
rect 5224 31084 5230 31096
rect 5353 31093 5365 31096
rect 5399 31093 5411 31127
rect 5353 31087 5411 31093
rect 6914 31084 6920 31136
rect 6972 31124 6978 31136
rect 7653 31127 7711 31133
rect 7653 31124 7665 31127
rect 6972 31096 7665 31124
rect 6972 31084 6978 31096
rect 7653 31093 7665 31096
rect 7699 31093 7711 31127
rect 8110 31124 8116 31136
rect 8071 31096 8116 31124
rect 7653 31087 7711 31093
rect 8110 31084 8116 31096
rect 8168 31084 8174 31136
rect 10134 31124 10140 31136
rect 10095 31096 10140 31124
rect 10134 31084 10140 31096
rect 10192 31084 10198 31136
rect 11238 31124 11244 31136
rect 11199 31096 11244 31124
rect 11238 31084 11244 31096
rect 11296 31124 11302 31136
rect 11422 31124 11428 31136
rect 11296 31096 11428 31124
rect 11296 31084 11302 31096
rect 11422 31084 11428 31096
rect 11480 31084 11486 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 7009 30923 7067 30929
rect 7009 30889 7021 30923
rect 7055 30920 7067 30923
rect 7282 30920 7288 30932
rect 7055 30892 7288 30920
rect 7055 30889 7067 30892
rect 7009 30883 7067 30889
rect 7282 30880 7288 30892
rect 7340 30880 7346 30932
rect 8110 30920 8116 30932
rect 8071 30892 8116 30920
rect 8110 30880 8116 30892
rect 8168 30880 8174 30932
rect 10229 30923 10287 30929
rect 10229 30889 10241 30923
rect 10275 30920 10287 30923
rect 10778 30920 10784 30932
rect 10275 30892 10784 30920
rect 10275 30889 10287 30892
rect 10229 30883 10287 30889
rect 10778 30880 10784 30892
rect 10836 30880 10842 30932
rect 11514 30880 11520 30932
rect 11572 30920 11578 30932
rect 11793 30923 11851 30929
rect 11793 30920 11805 30923
rect 11572 30892 11805 30920
rect 11572 30880 11578 30892
rect 11793 30889 11805 30892
rect 11839 30889 11851 30923
rect 11793 30883 11851 30889
rect 10680 30855 10738 30861
rect 10680 30821 10692 30855
rect 10726 30852 10738 30855
rect 11238 30852 11244 30864
rect 10726 30824 11244 30852
rect 10726 30821 10738 30824
rect 10680 30815 10738 30821
rect 11238 30812 11244 30824
rect 11296 30812 11302 30864
rect 3881 30787 3939 30793
rect 3881 30753 3893 30787
rect 3927 30784 3939 30787
rect 4430 30784 4436 30796
rect 3927 30756 4436 30784
rect 3927 30753 3939 30756
rect 3881 30747 3939 30753
rect 4430 30744 4436 30756
rect 4488 30744 4494 30796
rect 4525 30787 4583 30793
rect 4525 30753 4537 30787
rect 4571 30784 4583 30787
rect 4982 30784 4988 30796
rect 4571 30756 4988 30784
rect 4571 30753 4583 30756
rect 4525 30747 4583 30753
rect 4982 30744 4988 30756
rect 5040 30744 5046 30796
rect 7098 30744 7104 30796
rect 7156 30784 7162 30796
rect 7374 30784 7380 30796
rect 7156 30756 7380 30784
rect 7156 30744 7162 30756
rect 7374 30744 7380 30756
rect 7432 30744 7438 30796
rect 9674 30744 9680 30796
rect 9732 30784 9738 30796
rect 10226 30784 10232 30796
rect 9732 30756 10232 30784
rect 9732 30744 9738 30756
rect 10226 30744 10232 30756
rect 10284 30784 10290 30796
rect 10413 30787 10471 30793
rect 10413 30784 10425 30787
rect 10284 30756 10425 30784
rect 10284 30744 10290 30756
rect 10413 30753 10425 30756
rect 10459 30753 10471 30787
rect 10413 30747 10471 30753
rect 4338 30676 4344 30728
rect 4396 30716 4402 30728
rect 4617 30719 4675 30725
rect 4617 30716 4629 30719
rect 4396 30688 4629 30716
rect 4396 30676 4402 30688
rect 4617 30685 4629 30688
rect 4663 30685 4675 30719
rect 5626 30716 5632 30728
rect 5587 30688 5632 30716
rect 4617 30679 4675 30685
rect 5626 30676 5632 30688
rect 5684 30676 5690 30728
rect 7190 30676 7196 30728
rect 7248 30716 7254 30728
rect 7248 30688 7293 30716
rect 7248 30676 7254 30688
rect 2958 30580 2964 30592
rect 2919 30552 2964 30580
rect 2958 30540 2964 30552
rect 3016 30540 3022 30592
rect 4062 30580 4068 30592
rect 4023 30552 4068 30580
rect 4062 30540 4068 30552
rect 4120 30540 4126 30592
rect 5169 30583 5227 30589
rect 5169 30549 5181 30583
rect 5215 30580 5227 30583
rect 5258 30580 5264 30592
rect 5215 30552 5264 30580
rect 5215 30549 5227 30552
rect 5169 30543 5227 30549
rect 5258 30540 5264 30552
rect 5316 30540 5322 30592
rect 5534 30580 5540 30592
rect 5495 30552 5540 30580
rect 5534 30540 5540 30552
rect 5592 30540 5598 30592
rect 6638 30580 6644 30592
rect 6599 30552 6644 30580
rect 6638 30540 6644 30552
rect 6696 30540 6702 30592
rect 7745 30583 7803 30589
rect 7745 30549 7757 30583
rect 7791 30580 7803 30583
rect 7834 30580 7840 30592
rect 7791 30552 7840 30580
rect 7791 30549 7803 30552
rect 7745 30543 7803 30549
rect 7834 30540 7840 30552
rect 7892 30540 7898 30592
rect 8754 30540 8760 30592
rect 8812 30580 8818 30592
rect 9033 30583 9091 30589
rect 9033 30580 9045 30583
rect 8812 30552 9045 30580
rect 8812 30540 8818 30552
rect 9033 30549 9045 30552
rect 9079 30580 9091 30583
rect 9306 30580 9312 30592
rect 9079 30552 9312 30580
rect 9079 30549 9091 30552
rect 9033 30543 9091 30549
rect 9306 30540 9312 30552
rect 9364 30540 9370 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 7190 30376 7196 30388
rect 6840 30348 7196 30376
rect 2222 30308 2228 30320
rect 1412 30280 2228 30308
rect 1412 30181 1440 30280
rect 2222 30268 2228 30280
rect 2280 30268 2286 30320
rect 6273 30311 6331 30317
rect 6273 30277 6285 30311
rect 6319 30308 6331 30311
rect 6840 30308 6868 30348
rect 7190 30336 7196 30348
rect 7248 30336 7254 30388
rect 7377 30379 7435 30385
rect 7377 30345 7389 30379
rect 7423 30376 7435 30379
rect 8110 30376 8116 30388
rect 7423 30348 8116 30376
rect 7423 30345 7435 30348
rect 7377 30339 7435 30345
rect 8110 30336 8116 30348
rect 8168 30336 8174 30388
rect 9784 30348 10088 30376
rect 6319 30280 6868 30308
rect 8481 30311 8539 30317
rect 6319 30277 6331 30280
rect 6273 30271 6331 30277
rect 8481 30277 8493 30311
rect 8527 30308 8539 30311
rect 8570 30308 8576 30320
rect 8527 30280 8576 30308
rect 8527 30277 8539 30280
rect 8481 30271 8539 30277
rect 8570 30268 8576 30280
rect 8628 30308 8634 30320
rect 9784 30308 9812 30348
rect 9950 30308 9956 30320
rect 8628 30280 9812 30308
rect 9911 30280 9956 30308
rect 8628 30268 8634 30280
rect 1578 30240 1584 30252
rect 1539 30212 1584 30240
rect 1578 30200 1584 30212
rect 1636 30200 1642 30252
rect 4617 30243 4675 30249
rect 4617 30209 4629 30243
rect 4663 30240 4675 30243
rect 5350 30240 5356 30252
rect 4663 30212 5356 30240
rect 4663 30209 4675 30212
rect 4617 30203 4675 30209
rect 5350 30200 5356 30212
rect 5408 30240 5414 30252
rect 5629 30243 5687 30249
rect 5629 30240 5641 30243
rect 5408 30212 5641 30240
rect 5408 30200 5414 30212
rect 5629 30209 5641 30212
rect 5675 30209 5687 30243
rect 5629 30203 5687 30209
rect 6641 30243 6699 30249
rect 6641 30209 6653 30243
rect 6687 30240 6699 30243
rect 7098 30240 7104 30252
rect 6687 30212 7104 30240
rect 6687 30209 6699 30212
rect 6641 30203 6699 30209
rect 7098 30200 7104 30212
rect 7156 30240 7162 30252
rect 7282 30240 7288 30252
rect 7156 30212 7288 30240
rect 7156 30200 7162 30212
rect 7282 30200 7288 30212
rect 7340 30200 7346 30252
rect 8021 30243 8079 30249
rect 8021 30209 8033 30243
rect 8067 30240 8079 30243
rect 8202 30240 8208 30252
rect 8067 30212 8208 30240
rect 8067 30209 8079 30212
rect 8021 30203 8079 30209
rect 8202 30200 8208 30212
rect 8260 30200 8266 30252
rect 8386 30200 8392 30252
rect 8444 30240 8450 30252
rect 9508 30249 9536 30280
rect 9950 30268 9956 30280
rect 10008 30268 10014 30320
rect 8757 30243 8815 30249
rect 8757 30240 8769 30243
rect 8444 30212 8769 30240
rect 8444 30200 8450 30212
rect 8757 30209 8769 30212
rect 8803 30240 8815 30243
rect 9493 30243 9551 30249
rect 8803 30212 9260 30240
rect 8803 30209 8815 30212
rect 8757 30203 8815 30209
rect 1397 30175 1455 30181
rect 1397 30141 1409 30175
rect 1443 30141 1455 30175
rect 1397 30135 1455 30141
rect 2869 30175 2927 30181
rect 2869 30141 2881 30175
rect 2915 30172 2927 30175
rect 2958 30172 2964 30184
rect 2915 30144 2964 30172
rect 2915 30141 2927 30144
rect 2869 30135 2927 30141
rect 2958 30132 2964 30144
rect 3016 30172 3022 30184
rect 3418 30172 3424 30184
rect 3016 30144 3424 30172
rect 3016 30132 3022 30144
rect 3418 30132 3424 30144
rect 3476 30132 3482 30184
rect 2777 30107 2835 30113
rect 2777 30073 2789 30107
rect 2823 30104 2835 30107
rect 3136 30107 3194 30113
rect 3136 30104 3148 30107
rect 2823 30076 3148 30104
rect 2823 30073 2835 30076
rect 2777 30067 2835 30073
rect 3136 30073 3148 30076
rect 3182 30104 3194 30107
rect 3510 30104 3516 30116
rect 3182 30076 3516 30104
rect 3182 30073 3194 30076
rect 3136 30067 3194 30073
rect 3510 30064 3516 30076
rect 3568 30064 3574 30116
rect 5445 30107 5503 30113
rect 5445 30104 5457 30107
rect 4908 30076 5457 30104
rect 4908 30048 4936 30076
rect 5445 30073 5457 30076
rect 5491 30104 5503 30107
rect 5718 30104 5724 30116
rect 5491 30076 5724 30104
rect 5491 30073 5503 30076
rect 5445 30067 5503 30073
rect 5718 30064 5724 30076
rect 5776 30064 5782 30116
rect 7742 30104 7748 30116
rect 7655 30076 7748 30104
rect 7742 30064 7748 30076
rect 7800 30104 7806 30116
rect 7800 30076 8984 30104
rect 7800 30064 7806 30076
rect 4249 30039 4307 30045
rect 4249 30005 4261 30039
rect 4295 30036 4307 30039
rect 4338 30036 4344 30048
rect 4295 30008 4344 30036
rect 4295 30005 4307 30008
rect 4249 29999 4307 30005
rect 4338 29996 4344 30008
rect 4396 29996 4402 30048
rect 4890 30036 4896 30048
rect 4851 30008 4896 30036
rect 4890 29996 4896 30008
rect 4948 29996 4954 30048
rect 4982 29996 4988 30048
rect 5040 30036 5046 30048
rect 5077 30039 5135 30045
rect 5077 30036 5089 30039
rect 5040 30008 5089 30036
rect 5040 29996 5046 30008
rect 5077 30005 5089 30008
rect 5123 30005 5135 30039
rect 5077 29999 5135 30005
rect 5258 29996 5264 30048
rect 5316 30036 5322 30048
rect 5537 30039 5595 30045
rect 5537 30036 5549 30039
rect 5316 30008 5549 30036
rect 5316 29996 5322 30008
rect 5537 30005 5549 30008
rect 5583 30005 5595 30039
rect 5537 29999 5595 30005
rect 7101 30039 7159 30045
rect 7101 30005 7113 30039
rect 7147 30036 7159 30039
rect 7374 30036 7380 30048
rect 7147 30008 7380 30036
rect 7147 30005 7159 30008
rect 7101 29999 7159 30005
rect 7374 29996 7380 30008
rect 7432 29996 7438 30048
rect 7834 30036 7840 30048
rect 7795 30008 7840 30036
rect 7834 29996 7840 30008
rect 7892 29996 7898 30048
rect 8956 30045 8984 30076
rect 8941 30039 8999 30045
rect 8941 30005 8953 30039
rect 8987 30005 8999 30039
rect 9232 30036 9260 30212
rect 9493 30209 9505 30243
rect 9539 30209 9551 30243
rect 9493 30203 9551 30209
rect 9306 30132 9312 30184
rect 9364 30172 9370 30184
rect 9401 30175 9459 30181
rect 9401 30172 9413 30175
rect 9364 30144 9413 30172
rect 9364 30132 9370 30144
rect 9401 30141 9413 30144
rect 9447 30141 9459 30175
rect 9968 30172 9996 30268
rect 10060 30240 10088 30348
rect 11238 30336 11244 30388
rect 11296 30376 11302 30388
rect 11885 30379 11943 30385
rect 11885 30376 11897 30379
rect 11296 30348 11897 30376
rect 11296 30336 11302 30348
rect 11885 30345 11897 30348
rect 11931 30345 11943 30379
rect 11885 30339 11943 30345
rect 10594 30240 10600 30252
rect 10060 30212 10600 30240
rect 10594 30200 10600 30212
rect 10652 30240 10658 30252
rect 11057 30243 11115 30249
rect 11057 30240 11069 30243
rect 10652 30212 11069 30240
rect 10652 30200 10658 30212
rect 11057 30209 11069 30212
rect 11103 30240 11115 30243
rect 11517 30243 11575 30249
rect 11517 30240 11529 30243
rect 11103 30212 11529 30240
rect 11103 30209 11115 30212
rect 11057 30203 11115 30209
rect 11517 30209 11529 30212
rect 11563 30209 11575 30243
rect 11517 30203 11575 30209
rect 10873 30175 10931 30181
rect 10873 30172 10885 30175
rect 9968 30144 10885 30172
rect 9401 30135 9459 30141
rect 10873 30141 10885 30144
rect 10919 30141 10931 30175
rect 10873 30135 10931 30141
rect 10413 30107 10471 30113
rect 10413 30073 10425 30107
rect 10459 30104 10471 30107
rect 10459 30076 11008 30104
rect 10459 30073 10471 30076
rect 10413 30067 10471 30073
rect 10980 30048 11008 30076
rect 9309 30039 9367 30045
rect 9309 30036 9321 30039
rect 9232 30008 9321 30036
rect 8941 29999 8999 30005
rect 9309 30005 9321 30008
rect 9355 30036 9367 30039
rect 10134 30036 10140 30048
rect 9355 30008 10140 30036
rect 9355 30005 9367 30008
rect 9309 29999 9367 30005
rect 10134 29996 10140 30008
rect 10192 29996 10198 30048
rect 10502 30036 10508 30048
rect 10463 30008 10508 30036
rect 10502 29996 10508 30008
rect 10560 29996 10566 30048
rect 10962 30036 10968 30048
rect 10923 30008 10968 30036
rect 10962 29996 10968 30008
rect 11020 29996 11026 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 2774 29792 2780 29844
rect 2832 29832 2838 29844
rect 4062 29832 4068 29844
rect 2832 29804 4068 29832
rect 2832 29792 2838 29804
rect 4062 29792 4068 29804
rect 4120 29792 4126 29844
rect 4430 29792 4436 29844
rect 4488 29832 4494 29844
rect 4709 29835 4767 29841
rect 4709 29832 4721 29835
rect 4488 29804 4721 29832
rect 4488 29792 4494 29804
rect 4709 29801 4721 29804
rect 4755 29801 4767 29835
rect 4709 29795 4767 29801
rect 5534 29792 5540 29844
rect 5592 29832 5598 29844
rect 6273 29835 6331 29841
rect 6273 29832 6285 29835
rect 5592 29804 6285 29832
rect 5592 29792 5598 29804
rect 6273 29801 6285 29804
rect 6319 29801 6331 29835
rect 6273 29795 6331 29801
rect 6638 29792 6644 29844
rect 6696 29832 6702 29844
rect 6733 29835 6791 29841
rect 6733 29832 6745 29835
rect 6696 29804 6745 29832
rect 6696 29792 6702 29804
rect 6733 29801 6745 29804
rect 6779 29801 6791 29835
rect 7742 29832 7748 29844
rect 7703 29804 7748 29832
rect 6733 29795 6791 29801
rect 7742 29792 7748 29804
rect 7800 29792 7806 29844
rect 8018 29832 8024 29844
rect 7979 29804 8024 29832
rect 8018 29792 8024 29804
rect 8076 29792 8082 29844
rect 8294 29792 8300 29844
rect 8352 29832 8358 29844
rect 8481 29835 8539 29841
rect 8481 29832 8493 29835
rect 8352 29804 8493 29832
rect 8352 29792 8358 29804
rect 8481 29801 8493 29804
rect 8527 29832 8539 29835
rect 8846 29832 8852 29844
rect 8527 29804 8852 29832
rect 8527 29801 8539 29804
rect 8481 29795 8539 29801
rect 8846 29792 8852 29804
rect 8904 29792 8910 29844
rect 10226 29832 10232 29844
rect 10187 29804 10232 29832
rect 10226 29792 10232 29804
rect 10284 29832 10290 29844
rect 10413 29835 10471 29841
rect 10413 29832 10425 29835
rect 10284 29804 10425 29832
rect 10284 29792 10290 29804
rect 10413 29801 10425 29804
rect 10459 29832 10471 29835
rect 11238 29832 11244 29844
rect 10459 29804 11244 29832
rect 10459 29801 10471 29804
rect 10413 29795 10471 29801
rect 3881 29767 3939 29773
rect 3881 29733 3893 29767
rect 3927 29764 3939 29767
rect 4982 29764 4988 29776
rect 3927 29736 4988 29764
rect 3927 29733 3939 29736
rect 3881 29727 3939 29733
rect 4982 29724 4988 29736
rect 5040 29724 5046 29776
rect 5077 29767 5135 29773
rect 5077 29733 5089 29767
rect 5123 29764 5135 29767
rect 5166 29764 5172 29776
rect 5123 29736 5172 29764
rect 5123 29733 5135 29736
rect 5077 29727 5135 29733
rect 5166 29724 5172 29736
rect 5224 29764 5230 29776
rect 5626 29764 5632 29776
rect 5224 29736 5632 29764
rect 5224 29724 5230 29736
rect 5626 29724 5632 29736
rect 5684 29724 5690 29776
rect 8389 29767 8447 29773
rect 8389 29733 8401 29767
rect 8435 29764 8447 29767
rect 8570 29764 8576 29776
rect 8435 29736 8576 29764
rect 8435 29733 8447 29736
rect 8389 29727 8447 29733
rect 8570 29724 8576 29736
rect 8628 29764 8634 29776
rect 10502 29764 10508 29776
rect 8628 29736 10508 29764
rect 8628 29724 8634 29736
rect 10502 29724 10508 29736
rect 10560 29724 10566 29776
rect 2866 29696 2872 29708
rect 2827 29668 2872 29696
rect 2866 29656 2872 29668
rect 2924 29656 2930 29708
rect 5442 29656 5448 29708
rect 5500 29696 5506 29708
rect 6089 29699 6147 29705
rect 6089 29696 6101 29699
rect 5500 29668 6101 29696
rect 5500 29656 5506 29668
rect 5644 29640 5672 29668
rect 6089 29665 6101 29668
rect 6135 29665 6147 29699
rect 6089 29659 6147 29665
rect 6270 29656 6276 29708
rect 6328 29696 6334 29708
rect 10888 29705 10916 29804
rect 11238 29792 11244 29804
rect 11296 29792 11302 29844
rect 10962 29724 10968 29776
rect 11020 29764 11026 29776
rect 11140 29767 11198 29773
rect 11140 29764 11152 29767
rect 11020 29736 11152 29764
rect 11020 29724 11026 29736
rect 11140 29733 11152 29736
rect 11186 29764 11198 29767
rect 11514 29764 11520 29776
rect 11186 29736 11520 29764
rect 11186 29733 11198 29736
rect 11140 29727 11198 29733
rect 11514 29724 11520 29736
rect 11572 29724 11578 29776
rect 6641 29699 6699 29705
rect 6641 29696 6653 29699
rect 6328 29668 6653 29696
rect 6328 29656 6334 29668
rect 6641 29665 6653 29668
rect 6687 29665 6699 29699
rect 10597 29699 10655 29705
rect 10597 29696 10609 29699
rect 6641 29659 6699 29665
rect 10520 29668 10609 29696
rect 10520 29640 10548 29668
rect 10597 29665 10609 29668
rect 10643 29665 10655 29699
rect 10597 29659 10655 29665
rect 10873 29699 10931 29705
rect 10873 29665 10885 29699
rect 10919 29665 10931 29699
rect 10873 29659 10931 29665
rect 2958 29628 2964 29640
rect 2919 29600 2964 29628
rect 2958 29588 2964 29600
rect 3016 29628 3022 29640
rect 4154 29628 4160 29640
rect 3016 29600 4160 29628
rect 3016 29588 3022 29600
rect 4154 29588 4160 29600
rect 4212 29588 4218 29640
rect 5074 29588 5080 29640
rect 5132 29628 5138 29640
rect 5169 29631 5227 29637
rect 5169 29628 5181 29631
rect 5132 29600 5181 29628
rect 5132 29588 5138 29600
rect 5169 29597 5181 29600
rect 5215 29597 5227 29631
rect 5169 29591 5227 29597
rect 5353 29631 5411 29637
rect 5353 29597 5365 29631
rect 5399 29597 5411 29631
rect 5353 29591 5411 29597
rect 5368 29560 5396 29591
rect 5626 29588 5632 29640
rect 5684 29588 5690 29640
rect 6917 29631 6975 29637
rect 6917 29597 6929 29631
rect 6963 29628 6975 29631
rect 7006 29628 7012 29640
rect 6963 29600 7012 29628
rect 6963 29597 6975 29600
rect 6917 29591 6975 29597
rect 7006 29588 7012 29600
rect 7064 29588 7070 29640
rect 7469 29631 7527 29637
rect 7469 29597 7481 29631
rect 7515 29628 7527 29631
rect 8202 29628 8208 29640
rect 7515 29600 8208 29628
rect 7515 29597 7527 29600
rect 7469 29591 7527 29597
rect 8202 29588 8208 29600
rect 8260 29628 8266 29640
rect 8573 29631 8631 29637
rect 8573 29628 8585 29631
rect 8260 29600 8585 29628
rect 8260 29588 8266 29600
rect 8573 29597 8585 29600
rect 8619 29597 8631 29631
rect 8573 29591 8631 29597
rect 10502 29588 10508 29640
rect 10560 29588 10566 29640
rect 5442 29560 5448 29572
rect 5368 29532 5448 29560
rect 5442 29520 5448 29532
rect 5500 29520 5506 29572
rect 8754 29520 8760 29572
rect 8812 29560 8818 29572
rect 9582 29560 9588 29572
rect 8812 29532 9588 29560
rect 8812 29520 8818 29532
rect 9582 29520 9588 29532
rect 9640 29520 9646 29572
rect 1394 29452 1400 29504
rect 1452 29492 1458 29504
rect 2409 29495 2467 29501
rect 2409 29492 2421 29495
rect 1452 29464 2421 29492
rect 1452 29452 1458 29464
rect 2409 29461 2421 29464
rect 2455 29461 2467 29495
rect 3510 29492 3516 29504
rect 3471 29464 3516 29492
rect 2409 29455 2467 29461
rect 3510 29452 3516 29464
rect 3568 29452 3574 29504
rect 4338 29492 4344 29504
rect 4251 29464 4344 29492
rect 4338 29452 4344 29464
rect 4396 29492 4402 29504
rect 4614 29492 4620 29504
rect 4396 29464 4620 29492
rect 4396 29452 4402 29464
rect 4614 29452 4620 29464
rect 4672 29452 4678 29504
rect 5810 29492 5816 29504
rect 5771 29464 5816 29492
rect 5810 29452 5816 29464
rect 5868 29452 5874 29504
rect 9217 29495 9275 29501
rect 9217 29461 9229 29495
rect 9263 29492 9275 29495
rect 9490 29492 9496 29504
rect 9263 29464 9496 29492
rect 9263 29461 9275 29464
rect 9217 29455 9275 29461
rect 9490 29452 9496 29464
rect 9548 29452 9554 29504
rect 11514 29452 11520 29504
rect 11572 29492 11578 29504
rect 12253 29495 12311 29501
rect 12253 29492 12265 29495
rect 11572 29464 12265 29492
rect 11572 29452 11578 29464
rect 12253 29461 12265 29464
rect 12299 29461 12311 29495
rect 12253 29455 12311 29461
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 1578 29288 1584 29300
rect 1539 29260 1584 29288
rect 1578 29248 1584 29260
rect 1636 29248 1642 29300
rect 2501 29291 2559 29297
rect 2501 29257 2513 29291
rect 2547 29288 2559 29291
rect 2958 29288 2964 29300
rect 2547 29260 2964 29288
rect 2547 29257 2559 29260
rect 2501 29251 2559 29257
rect 2958 29248 2964 29260
rect 3016 29248 3022 29300
rect 4801 29291 4859 29297
rect 4801 29257 4813 29291
rect 4847 29288 4859 29291
rect 5074 29288 5080 29300
rect 4847 29260 5080 29288
rect 4847 29257 4859 29260
rect 4801 29251 4859 29257
rect 5074 29248 5080 29260
rect 5132 29248 5138 29300
rect 7006 29288 7012 29300
rect 6967 29260 7012 29288
rect 7006 29248 7012 29260
rect 7064 29248 7070 29300
rect 8113 29291 8171 29297
rect 8113 29257 8125 29291
rect 8159 29288 8171 29291
rect 8202 29288 8208 29300
rect 8159 29260 8208 29288
rect 8159 29257 8171 29260
rect 8113 29251 8171 29257
rect 8202 29248 8208 29260
rect 8260 29248 8266 29300
rect 10962 29288 10968 29300
rect 10923 29260 10968 29288
rect 10962 29248 10968 29260
rect 11020 29248 11026 29300
rect 11238 29288 11244 29300
rect 11199 29260 11244 29288
rect 11238 29248 11244 29260
rect 11296 29248 11302 29300
rect 3421 29223 3479 29229
rect 3421 29189 3433 29223
rect 3467 29220 3479 29223
rect 4154 29220 4160 29232
rect 3467 29192 4160 29220
rect 3467 29189 3479 29192
rect 3421 29183 3479 29189
rect 4154 29180 4160 29192
rect 4212 29180 4218 29232
rect 5169 29223 5227 29229
rect 5169 29189 5181 29223
rect 5215 29220 5227 29223
rect 5350 29220 5356 29232
rect 5215 29192 5356 29220
rect 5215 29189 5227 29192
rect 5169 29183 5227 29189
rect 5350 29180 5356 29192
rect 5408 29180 5414 29232
rect 9125 29223 9183 29229
rect 9125 29189 9137 29223
rect 9171 29220 9183 29223
rect 9582 29220 9588 29232
rect 9171 29192 9588 29220
rect 9171 29189 9183 29192
rect 9125 29183 9183 29189
rect 9582 29180 9588 29192
rect 9640 29180 9646 29232
rect 2038 29152 2044 29164
rect 1412 29124 2044 29152
rect 1412 29093 1440 29124
rect 2038 29112 2044 29124
rect 2096 29112 2102 29164
rect 3510 29112 3516 29164
rect 3568 29152 3574 29164
rect 4065 29155 4123 29161
rect 4065 29152 4077 29155
rect 3568 29124 4077 29152
rect 3568 29112 3574 29124
rect 4065 29121 4077 29124
rect 4111 29152 4123 29155
rect 4338 29152 4344 29164
rect 4111 29124 4344 29152
rect 4111 29121 4123 29124
rect 4065 29115 4123 29121
rect 4338 29112 4344 29124
rect 4396 29152 4402 29164
rect 5442 29152 5448 29164
rect 4396 29124 5448 29152
rect 4396 29112 4402 29124
rect 5442 29112 5448 29124
rect 5500 29112 5506 29164
rect 5626 29152 5632 29164
rect 5587 29124 5632 29152
rect 5626 29112 5632 29124
rect 5684 29112 5690 29164
rect 5810 29152 5816 29164
rect 5771 29124 5816 29152
rect 5810 29112 5816 29124
rect 5868 29112 5874 29164
rect 9490 29112 9496 29164
rect 9548 29152 9554 29164
rect 9677 29155 9735 29161
rect 9677 29152 9689 29155
rect 9548 29124 9689 29152
rect 9548 29112 9554 29124
rect 9677 29121 9689 29124
rect 9723 29121 9735 29155
rect 9677 29115 9735 29121
rect 1397 29087 1455 29093
rect 1397 29053 1409 29087
rect 1443 29053 1455 29087
rect 5534 29084 5540 29096
rect 5495 29056 5540 29084
rect 1397 29047 1455 29053
rect 5534 29044 5540 29056
rect 5592 29044 5598 29096
rect 8481 29087 8539 29093
rect 8481 29053 8493 29087
rect 8527 29084 8539 29087
rect 8846 29084 8852 29096
rect 8527 29056 8852 29084
rect 8527 29053 8539 29056
rect 8481 29047 8539 29053
rect 8846 29044 8852 29056
rect 8904 29084 8910 29096
rect 10137 29087 10195 29093
rect 10137 29084 10149 29087
rect 8904 29056 10149 29084
rect 8904 29044 8910 29056
rect 10137 29053 10149 29056
rect 10183 29053 10195 29087
rect 10137 29047 10195 29053
rect 3234 28976 3240 29028
rect 3292 29016 3298 29028
rect 3329 29019 3387 29025
rect 3329 29016 3341 29019
rect 3292 28988 3341 29016
rect 3292 28976 3298 28988
rect 3329 28985 3341 28988
rect 3375 29016 3387 29019
rect 3789 29019 3847 29025
rect 3789 29016 3801 29019
rect 3375 28988 3801 29016
rect 3375 28985 3387 28988
rect 3329 28979 3387 28985
rect 3789 28985 3801 28988
rect 3835 29016 3847 29019
rect 3970 29016 3976 29028
rect 3835 28988 3976 29016
rect 3835 28985 3847 28988
rect 3789 28979 3847 28985
rect 3970 28976 3976 28988
rect 4028 28976 4034 29028
rect 5994 28976 6000 29028
rect 6052 29016 6058 29028
rect 6270 29016 6276 29028
rect 6052 28988 6276 29016
rect 6052 28976 6058 28988
rect 6270 28976 6276 28988
rect 6328 28976 6334 29028
rect 8938 29016 8944 29028
rect 8899 28988 8944 29016
rect 8938 28976 8944 28988
rect 8996 29016 9002 29028
rect 9585 29019 9643 29025
rect 9585 29016 9597 29019
rect 8996 28988 9597 29016
rect 8996 28976 9002 28988
rect 9585 28985 9597 28988
rect 9631 29016 9643 29019
rect 9674 29016 9680 29028
rect 9631 28988 9680 29016
rect 9631 28985 9643 28988
rect 9585 28979 9643 28985
rect 9674 28976 9680 28988
rect 9732 28976 9738 29028
rect 10042 28976 10048 29028
rect 10100 29016 10106 29028
rect 10318 29016 10324 29028
rect 10100 28988 10324 29016
rect 10100 28976 10106 28988
rect 10318 28976 10324 28988
rect 10376 28976 10382 29028
rect 10502 29016 10508 29028
rect 10463 28988 10508 29016
rect 10502 28976 10508 28988
rect 10560 28976 10566 29028
rect 11974 28976 11980 29028
rect 12032 29016 12038 29028
rect 12066 29016 12072 29028
rect 12032 28988 12072 29016
rect 12032 28976 12038 28988
rect 12066 28976 12072 28988
rect 12124 28976 12130 29028
rect 2866 28948 2872 28960
rect 2827 28920 2872 28948
rect 2866 28908 2872 28920
rect 2924 28908 2930 28960
rect 3510 28908 3516 28960
rect 3568 28948 3574 28960
rect 3881 28951 3939 28957
rect 3881 28948 3893 28951
rect 3568 28920 3893 28948
rect 3568 28908 3574 28920
rect 3881 28917 3893 28920
rect 3927 28948 3939 28951
rect 6914 28948 6920 28960
rect 3927 28920 6920 28948
rect 3927 28917 3939 28920
rect 3881 28911 3939 28917
rect 6914 28908 6920 28920
rect 6972 28908 6978 28960
rect 7285 28951 7343 28957
rect 7285 28917 7297 28951
rect 7331 28948 7343 28951
rect 7466 28948 7472 28960
rect 7331 28920 7472 28948
rect 7331 28917 7343 28920
rect 7285 28911 7343 28917
rect 7466 28908 7472 28920
rect 7524 28908 7530 28960
rect 8297 28951 8355 28957
rect 8297 28917 8309 28951
rect 8343 28948 8355 28951
rect 8386 28948 8392 28960
rect 8343 28920 8392 28948
rect 8343 28917 8355 28920
rect 8297 28911 8355 28917
rect 8386 28908 8392 28920
rect 8444 28908 8450 28960
rect 9214 28908 9220 28960
rect 9272 28948 9278 28960
rect 9493 28951 9551 28957
rect 9493 28948 9505 28951
rect 9272 28920 9505 28948
rect 9272 28908 9278 28920
rect 9493 28917 9505 28920
rect 9539 28917 9551 28951
rect 9493 28911 9551 28917
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 2501 28747 2559 28753
rect 2501 28713 2513 28747
rect 2547 28744 2559 28747
rect 2774 28744 2780 28756
rect 2547 28716 2780 28744
rect 2547 28713 2559 28716
rect 2501 28707 2559 28713
rect 2774 28704 2780 28716
rect 2832 28704 2838 28756
rect 2866 28704 2872 28756
rect 2924 28744 2930 28756
rect 4065 28747 4123 28753
rect 4065 28744 4077 28747
rect 2924 28716 4077 28744
rect 2924 28704 2930 28716
rect 4065 28713 4077 28716
rect 4111 28713 4123 28747
rect 4065 28707 4123 28713
rect 4154 28704 4160 28756
rect 4212 28744 4218 28756
rect 4433 28747 4491 28753
rect 4433 28744 4445 28747
rect 4212 28716 4445 28744
rect 4212 28704 4218 28716
rect 4433 28713 4445 28716
rect 4479 28713 4491 28747
rect 5166 28744 5172 28756
rect 5127 28716 5172 28744
rect 4433 28707 4491 28713
rect 5166 28704 5172 28716
rect 5224 28704 5230 28756
rect 6365 28747 6423 28753
rect 6365 28713 6377 28747
rect 6411 28744 6423 28747
rect 6638 28744 6644 28756
rect 6411 28716 6644 28744
rect 6411 28713 6423 28716
rect 6365 28707 6423 28713
rect 6638 28704 6644 28716
rect 6696 28704 6702 28756
rect 7006 28744 7012 28756
rect 6967 28716 7012 28744
rect 7006 28704 7012 28716
rect 7064 28704 7070 28756
rect 8202 28744 8208 28756
rect 8163 28716 8208 28744
rect 8202 28704 8208 28716
rect 8260 28704 8266 28756
rect 8570 28744 8576 28756
rect 8531 28716 8576 28744
rect 8570 28704 8576 28716
rect 8628 28704 8634 28756
rect 9953 28747 10011 28753
rect 9953 28713 9965 28747
rect 9999 28744 10011 28747
rect 10226 28744 10232 28756
rect 9999 28716 10232 28744
rect 9999 28713 10011 28716
rect 9953 28707 10011 28713
rect 10226 28704 10232 28716
rect 10284 28704 10290 28756
rect 3510 28676 3516 28688
rect 3471 28648 3516 28676
rect 3510 28636 3516 28648
rect 3568 28636 3574 28688
rect 4982 28636 4988 28688
rect 5040 28676 5046 28688
rect 7098 28676 7104 28688
rect 5040 28648 7104 28676
rect 5040 28636 5046 28648
rect 7098 28636 7104 28648
rect 7156 28636 7162 28688
rect 7466 28676 7472 28688
rect 7427 28648 7472 28676
rect 7466 28636 7472 28648
rect 7524 28636 7530 28688
rect 4525 28611 4583 28617
rect 4525 28608 4537 28611
rect 4448 28580 4537 28608
rect 4448 28472 4476 28580
rect 4525 28577 4537 28580
rect 4571 28577 4583 28611
rect 4525 28571 4583 28577
rect 5442 28568 5448 28620
rect 5500 28608 5506 28620
rect 5537 28611 5595 28617
rect 5537 28608 5549 28611
rect 5500 28580 5549 28608
rect 5500 28568 5506 28580
rect 5537 28577 5549 28580
rect 5583 28608 5595 28611
rect 5718 28608 5724 28620
rect 5583 28580 5724 28608
rect 5583 28577 5595 28580
rect 5537 28571 5595 28577
rect 5718 28568 5724 28580
rect 5776 28568 5782 28620
rect 5902 28608 5908 28620
rect 5863 28580 5908 28608
rect 5902 28568 5908 28580
rect 5960 28568 5966 28620
rect 7558 28608 7564 28620
rect 7519 28580 7564 28608
rect 7558 28568 7564 28580
rect 7616 28568 7622 28620
rect 10689 28611 10747 28617
rect 10689 28608 10701 28611
rect 9508 28580 10701 28608
rect 4614 28540 4620 28552
rect 4575 28512 4620 28540
rect 4614 28500 4620 28512
rect 4672 28500 4678 28552
rect 7006 28500 7012 28552
rect 7064 28540 7070 28552
rect 7653 28543 7711 28549
rect 7653 28540 7665 28543
rect 7064 28512 7665 28540
rect 7064 28500 7070 28512
rect 7653 28509 7665 28512
rect 7699 28540 7711 28543
rect 7742 28540 7748 28552
rect 7699 28512 7748 28540
rect 7699 28509 7711 28512
rect 7653 28503 7711 28509
rect 7742 28500 7748 28512
rect 7800 28500 7806 28552
rect 7926 28500 7932 28552
rect 7984 28540 7990 28552
rect 9125 28543 9183 28549
rect 9125 28540 9137 28543
rect 7984 28512 9137 28540
rect 7984 28500 7990 28512
rect 9125 28509 9137 28512
rect 9171 28540 9183 28543
rect 9214 28540 9220 28552
rect 9171 28512 9220 28540
rect 9171 28509 9183 28512
rect 9125 28503 9183 28509
rect 9214 28500 9220 28512
rect 9272 28540 9278 28552
rect 9508 28540 9536 28580
rect 10689 28577 10701 28580
rect 10735 28608 10747 28611
rect 11054 28608 11060 28620
rect 10735 28580 11060 28608
rect 10735 28577 10747 28580
rect 10689 28571 10747 28577
rect 11054 28568 11060 28580
rect 11112 28568 11118 28620
rect 9272 28512 9536 28540
rect 9272 28500 9278 28512
rect 9674 28500 9680 28552
rect 9732 28540 9738 28552
rect 10778 28540 10784 28552
rect 9732 28512 10784 28540
rect 9732 28500 9738 28512
rect 10778 28500 10784 28512
rect 10836 28500 10842 28552
rect 10965 28543 11023 28549
rect 10965 28509 10977 28543
rect 11011 28540 11023 28543
rect 11514 28540 11520 28552
rect 11011 28512 11520 28540
rect 11011 28509 11023 28512
rect 10965 28503 11023 28509
rect 11514 28500 11520 28512
rect 11572 28500 11578 28552
rect 4522 28472 4528 28484
rect 4448 28444 4528 28472
rect 4522 28432 4528 28444
rect 4580 28432 4586 28484
rect 5534 28432 5540 28484
rect 5592 28472 5598 28484
rect 7101 28475 7159 28481
rect 7101 28472 7113 28475
rect 5592 28444 7113 28472
rect 5592 28432 5598 28444
rect 7101 28441 7113 28444
rect 7147 28441 7159 28475
rect 7101 28435 7159 28441
rect 3881 28407 3939 28413
rect 3881 28373 3893 28407
rect 3927 28404 3939 28407
rect 4062 28404 4068 28416
rect 3927 28376 4068 28404
rect 3927 28373 3939 28376
rect 3881 28367 3939 28373
rect 4062 28364 4068 28376
rect 4120 28364 4126 28416
rect 5258 28364 5264 28416
rect 5316 28404 5322 28416
rect 5721 28407 5779 28413
rect 5721 28404 5733 28407
rect 5316 28376 5733 28404
rect 5316 28364 5322 28376
rect 5721 28373 5733 28376
rect 5767 28373 5779 28407
rect 5721 28367 5779 28373
rect 6914 28364 6920 28416
rect 6972 28404 6978 28416
rect 8110 28404 8116 28416
rect 6972 28376 8116 28404
rect 6972 28364 6978 28376
rect 8110 28364 8116 28376
rect 8168 28364 8174 28416
rect 10318 28404 10324 28416
rect 10279 28376 10324 28404
rect 10318 28364 10324 28376
rect 10376 28364 10382 28416
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 2038 28200 2044 28212
rect 1999 28172 2044 28200
rect 2038 28160 2044 28172
rect 2096 28160 2102 28212
rect 3326 28160 3332 28212
rect 3384 28200 3390 28212
rect 3421 28203 3479 28209
rect 3421 28200 3433 28203
rect 3384 28172 3433 28200
rect 3384 28160 3390 28172
rect 3421 28169 3433 28172
rect 3467 28169 3479 28203
rect 4614 28200 4620 28212
rect 4575 28172 4620 28200
rect 3421 28163 3479 28169
rect 1581 28135 1639 28141
rect 1581 28101 1593 28135
rect 1627 28132 1639 28135
rect 2590 28132 2596 28144
rect 1627 28104 2596 28132
rect 1627 28101 1639 28104
rect 1581 28095 1639 28101
rect 2590 28092 2596 28104
rect 2648 28092 2654 28144
rect 1397 27999 1455 28005
rect 1397 27965 1409 27999
rect 1443 27996 1455 27999
rect 2038 27996 2044 28008
rect 1443 27968 2044 27996
rect 1443 27965 1455 27968
rect 1397 27959 1455 27965
rect 2038 27956 2044 27968
rect 2096 27956 2102 28008
rect 3436 27996 3464 28163
rect 4614 28160 4620 28172
rect 4672 28160 4678 28212
rect 6641 28203 6699 28209
rect 6641 28169 6653 28203
rect 6687 28200 6699 28203
rect 6822 28200 6828 28212
rect 6687 28172 6828 28200
rect 6687 28169 6699 28172
rect 6641 28163 6699 28169
rect 6822 28160 6828 28172
rect 6880 28200 6886 28212
rect 6880 28172 7328 28200
rect 6880 28160 6886 28172
rect 7009 28135 7067 28141
rect 7009 28132 7021 28135
rect 5644 28104 7021 28132
rect 5644 28076 5672 28104
rect 7009 28101 7021 28104
rect 7055 28101 7067 28135
rect 7009 28095 7067 28101
rect 3694 28024 3700 28076
rect 3752 28064 3758 28076
rect 4249 28067 4307 28073
rect 4249 28064 4261 28067
rect 3752 28036 4261 28064
rect 3752 28024 3758 28036
rect 4249 28033 4261 28036
rect 4295 28064 4307 28067
rect 4338 28064 4344 28076
rect 4295 28036 4344 28064
rect 4295 28033 4307 28036
rect 4249 28027 4307 28033
rect 4338 28024 4344 28036
rect 4396 28024 4402 28076
rect 5626 28064 5632 28076
rect 5539 28036 5632 28064
rect 5626 28024 5632 28036
rect 5684 28024 5690 28076
rect 5810 28064 5816 28076
rect 5723 28036 5816 28064
rect 5810 28024 5816 28036
rect 5868 28064 5874 28076
rect 6730 28064 6736 28076
rect 5868 28036 6736 28064
rect 5868 28024 5874 28036
rect 6730 28024 6736 28036
rect 6788 28024 6794 28076
rect 3973 27999 4031 28005
rect 3973 27996 3985 27999
rect 3436 27968 3985 27996
rect 3973 27965 3985 27968
rect 4019 27965 4031 27999
rect 5534 27996 5540 28008
rect 5495 27968 5540 27996
rect 3973 27959 4031 27965
rect 5534 27956 5540 27968
rect 5592 27956 5598 28008
rect 3145 27931 3203 27937
rect 3145 27897 3157 27931
rect 3191 27928 3203 27931
rect 4062 27928 4068 27940
rect 3191 27900 4068 27928
rect 3191 27897 3203 27900
rect 3145 27891 3203 27897
rect 4062 27888 4068 27900
rect 4120 27888 4126 27940
rect 5077 27931 5135 27937
rect 5077 27897 5089 27931
rect 5123 27928 5135 27931
rect 5828 27928 5856 28024
rect 7300 27996 7328 28172
rect 7466 28160 7472 28212
rect 7524 28200 7530 28212
rect 8021 28203 8079 28209
rect 8021 28200 8033 28203
rect 7524 28172 8033 28200
rect 7524 28160 7530 28172
rect 8021 28169 8033 28172
rect 8067 28169 8079 28203
rect 8021 28163 8079 28169
rect 10413 28203 10471 28209
rect 10413 28169 10425 28203
rect 10459 28200 10471 28203
rect 10594 28200 10600 28212
rect 10459 28172 10600 28200
rect 10459 28169 10471 28172
rect 10413 28163 10471 28169
rect 10594 28160 10600 28172
rect 10652 28160 10658 28212
rect 10778 28200 10784 28212
rect 10739 28172 10784 28200
rect 10778 28160 10784 28172
rect 10836 28160 10842 28212
rect 11054 28200 11060 28212
rect 11015 28172 11060 28200
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 11514 28200 11520 28212
rect 11475 28172 11520 28200
rect 11514 28160 11520 28172
rect 11572 28160 11578 28212
rect 8110 28092 8116 28144
rect 8168 28132 8174 28144
rect 8754 28132 8760 28144
rect 8168 28104 8760 28132
rect 8168 28092 8174 28104
rect 8754 28092 8760 28104
rect 8812 28092 8818 28144
rect 7466 28064 7472 28076
rect 7427 28036 7472 28064
rect 7466 28024 7472 28036
rect 7524 28024 7530 28076
rect 7653 28067 7711 28073
rect 7653 28033 7665 28067
rect 7699 28064 7711 28067
rect 7742 28064 7748 28076
rect 7699 28036 7748 28064
rect 7699 28033 7711 28036
rect 7653 28027 7711 28033
rect 7742 28024 7748 28036
rect 7800 28064 7806 28076
rect 8481 28067 8539 28073
rect 8481 28064 8493 28067
rect 7800 28036 8493 28064
rect 7800 28024 7806 28036
rect 8481 28033 8493 28036
rect 8527 28033 8539 28067
rect 8481 28027 8539 28033
rect 7377 27999 7435 28005
rect 7377 27996 7389 27999
rect 7300 27968 7389 27996
rect 7377 27965 7389 27968
rect 7423 27996 7435 27999
rect 8202 27996 8208 28008
rect 7423 27968 8208 27996
rect 7423 27965 7435 27968
rect 7377 27959 7435 27965
rect 8202 27956 8208 27968
rect 8260 27956 8266 28008
rect 8386 27956 8392 28008
rect 8444 27996 8450 28008
rect 8941 27999 8999 28005
rect 8941 27996 8953 27999
rect 8444 27968 8953 27996
rect 8444 27956 8450 27968
rect 8941 27965 8953 27968
rect 8987 27965 8999 27999
rect 8941 27959 8999 27965
rect 9033 27999 9091 28005
rect 9033 27965 9045 27999
rect 9079 27996 9091 27999
rect 10226 27996 10232 28008
rect 9079 27968 10232 27996
rect 9079 27965 9091 27968
rect 9033 27959 9091 27965
rect 5123 27900 5856 27928
rect 6273 27931 6331 27937
rect 5123 27897 5135 27900
rect 5077 27891 5135 27897
rect 6273 27897 6285 27931
rect 6319 27928 6331 27931
rect 7558 27928 7564 27940
rect 6319 27900 7564 27928
rect 6319 27897 6331 27900
rect 6273 27891 6331 27897
rect 7558 27888 7564 27900
rect 7616 27888 7622 27940
rect 8956 27928 8984 27959
rect 10226 27956 10232 27968
rect 10284 27956 10290 28008
rect 9300 27931 9358 27937
rect 8956 27900 9260 27928
rect 9232 27872 9260 27900
rect 9300 27897 9312 27931
rect 9346 27928 9358 27931
rect 9490 27928 9496 27940
rect 9346 27900 9496 27928
rect 9346 27897 9358 27900
rect 9300 27891 9358 27897
rect 9490 27888 9496 27900
rect 9548 27888 9554 27940
rect 3605 27863 3663 27869
rect 3605 27829 3617 27863
rect 3651 27860 3663 27863
rect 4522 27860 4528 27872
rect 3651 27832 4528 27860
rect 3651 27829 3663 27832
rect 3605 27823 3663 27829
rect 4522 27820 4528 27832
rect 4580 27820 4586 27872
rect 5169 27863 5227 27869
rect 5169 27829 5181 27863
rect 5215 27860 5227 27863
rect 5442 27860 5448 27872
rect 5215 27832 5448 27860
rect 5215 27829 5227 27832
rect 5169 27823 5227 27829
rect 5442 27820 5448 27832
rect 5500 27820 5506 27872
rect 8754 27860 8760 27872
rect 8715 27832 8760 27860
rect 8754 27820 8760 27832
rect 8812 27820 8818 27872
rect 9214 27820 9220 27872
rect 9272 27820 9278 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 3694 27656 3700 27668
rect 3655 27628 3700 27656
rect 3694 27616 3700 27628
rect 3752 27616 3758 27668
rect 4341 27659 4399 27665
rect 4341 27625 4353 27659
rect 4387 27656 4399 27659
rect 4522 27656 4528 27668
rect 4387 27628 4528 27656
rect 4387 27625 4399 27628
rect 4341 27619 4399 27625
rect 4522 27616 4528 27628
rect 4580 27616 4586 27668
rect 5626 27656 5632 27668
rect 5552 27628 5632 27656
rect 4154 27548 4160 27600
rect 4212 27588 4218 27600
rect 4617 27591 4675 27597
rect 4617 27588 4629 27591
rect 4212 27560 4629 27588
rect 4212 27548 4218 27560
rect 4617 27557 4629 27560
rect 4663 27557 4675 27591
rect 4617 27551 4675 27557
rect 5077 27591 5135 27597
rect 5077 27557 5089 27591
rect 5123 27588 5135 27591
rect 5552 27588 5580 27628
rect 5626 27616 5632 27628
rect 5684 27616 5690 27668
rect 7098 27656 7104 27668
rect 7011 27628 7104 27656
rect 7098 27616 7104 27628
rect 7156 27656 7162 27668
rect 7466 27656 7472 27668
rect 7156 27628 7472 27656
rect 7156 27616 7162 27628
rect 7466 27616 7472 27628
rect 7524 27616 7530 27668
rect 8757 27659 8815 27665
rect 8757 27625 8769 27659
rect 8803 27656 8815 27659
rect 9125 27659 9183 27665
rect 9125 27656 9137 27659
rect 8803 27628 9137 27656
rect 8803 27625 8815 27628
rect 8757 27619 8815 27625
rect 9125 27625 9137 27628
rect 9171 27656 9183 27659
rect 9490 27656 9496 27668
rect 9171 27628 9496 27656
rect 9171 27625 9183 27628
rect 9125 27619 9183 27625
rect 9490 27616 9496 27628
rect 9548 27616 9554 27668
rect 10318 27616 10324 27668
rect 10376 27656 10382 27668
rect 10778 27656 10784 27668
rect 10376 27628 10784 27656
rect 10376 27616 10382 27628
rect 10778 27616 10784 27628
rect 10836 27656 10842 27668
rect 10965 27659 11023 27665
rect 10965 27656 10977 27659
rect 10836 27628 10977 27656
rect 10836 27616 10842 27628
rect 10965 27625 10977 27628
rect 11011 27625 11023 27659
rect 10965 27619 11023 27625
rect 5123 27560 5580 27588
rect 5123 27557 5135 27560
rect 5077 27551 5135 27557
rect 11514 27548 11520 27600
rect 11572 27588 11578 27600
rect 11762 27591 11820 27597
rect 11762 27588 11774 27591
rect 11572 27560 11774 27588
rect 11572 27548 11578 27560
rect 11762 27557 11774 27560
rect 11808 27557 11820 27591
rect 11762 27551 11820 27557
rect 5169 27523 5227 27529
rect 5169 27489 5181 27523
rect 5215 27520 5227 27523
rect 5258 27520 5264 27532
rect 5215 27492 5264 27520
rect 5215 27489 5227 27492
rect 5169 27483 5227 27489
rect 5258 27480 5264 27492
rect 5316 27480 5322 27532
rect 5436 27523 5494 27529
rect 5436 27489 5448 27523
rect 5482 27520 5494 27523
rect 6822 27520 6828 27532
rect 5482 27492 6828 27520
rect 5482 27489 5494 27492
rect 5436 27483 5494 27489
rect 6822 27480 6828 27492
rect 6880 27480 6886 27532
rect 7190 27480 7196 27532
rect 7248 27520 7254 27532
rect 7633 27523 7691 27529
rect 7633 27520 7645 27523
rect 7248 27492 7645 27520
rect 7248 27480 7254 27492
rect 7633 27489 7645 27492
rect 7679 27489 7691 27523
rect 7633 27483 7691 27489
rect 9122 27480 9128 27532
rect 9180 27520 9186 27532
rect 9766 27520 9772 27532
rect 9180 27492 9772 27520
rect 9180 27480 9186 27492
rect 9766 27480 9772 27492
rect 9824 27520 9830 27532
rect 10321 27523 10379 27529
rect 10321 27520 10333 27523
rect 9824 27492 10333 27520
rect 9824 27480 9830 27492
rect 10321 27489 10333 27492
rect 10367 27489 10379 27523
rect 11532 27520 11560 27548
rect 10321 27483 10379 27489
rect 10612 27492 11560 27520
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27421 7435 27455
rect 7377 27415 7435 27421
rect 4614 27276 4620 27328
rect 4672 27316 4678 27328
rect 4890 27316 4896 27328
rect 4672 27288 4896 27316
rect 4672 27276 4678 27288
rect 4890 27276 4896 27288
rect 4948 27276 4954 27328
rect 6549 27319 6607 27325
rect 6549 27285 6561 27319
rect 6595 27316 6607 27319
rect 6730 27316 6736 27328
rect 6595 27288 6736 27316
rect 6595 27285 6607 27288
rect 6549 27279 6607 27285
rect 6730 27276 6736 27288
rect 6788 27276 6794 27328
rect 7392 27316 7420 27415
rect 10226 27412 10232 27464
rect 10284 27452 10290 27464
rect 10612 27461 10640 27492
rect 10413 27455 10471 27461
rect 10413 27452 10425 27455
rect 10284 27424 10425 27452
rect 10284 27412 10290 27424
rect 10413 27421 10425 27424
rect 10459 27421 10471 27455
rect 10413 27415 10471 27421
rect 10597 27455 10655 27461
rect 10597 27421 10609 27455
rect 10643 27421 10655 27455
rect 10597 27415 10655 27421
rect 11422 27412 11428 27464
rect 11480 27452 11486 27464
rect 11517 27455 11575 27461
rect 11517 27452 11529 27455
rect 11480 27424 11529 27452
rect 11480 27412 11486 27424
rect 11517 27421 11529 27424
rect 11563 27421 11575 27455
rect 11517 27415 11575 27421
rect 7558 27316 7564 27328
rect 7392 27288 7564 27316
rect 7558 27276 7564 27288
rect 7616 27276 7622 27328
rect 9306 27276 9312 27328
rect 9364 27316 9370 27328
rect 9401 27319 9459 27325
rect 9401 27316 9413 27319
rect 9364 27288 9413 27316
rect 9364 27276 9370 27288
rect 9401 27285 9413 27288
rect 9447 27285 9459 27319
rect 9401 27279 9459 27285
rect 9953 27319 10011 27325
rect 9953 27285 9965 27319
rect 9999 27316 10011 27319
rect 10686 27316 10692 27328
rect 9999 27288 10692 27316
rect 9999 27285 10011 27288
rect 9953 27279 10011 27285
rect 10686 27276 10692 27288
rect 10744 27276 10750 27328
rect 12894 27316 12900 27328
rect 12855 27288 12900 27316
rect 12894 27276 12900 27288
rect 12952 27276 12958 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 3418 27112 3424 27124
rect 3331 27084 3424 27112
rect 3418 27072 3424 27084
rect 3476 27112 3482 27124
rect 5258 27112 5264 27124
rect 3476 27084 5264 27112
rect 3476 27072 3482 27084
rect 5258 27072 5264 27084
rect 5316 27072 5322 27124
rect 5629 27115 5687 27121
rect 5629 27081 5641 27115
rect 5675 27112 5687 27115
rect 5718 27112 5724 27124
rect 5675 27084 5724 27112
rect 5675 27081 5687 27084
rect 5629 27075 5687 27081
rect 5718 27072 5724 27084
rect 5776 27072 5782 27124
rect 5902 27072 5908 27124
rect 5960 27112 5966 27124
rect 6457 27115 6515 27121
rect 6457 27112 6469 27115
rect 5960 27084 6469 27112
rect 5960 27072 5966 27084
rect 6457 27081 6469 27084
rect 6503 27112 6515 27115
rect 6638 27112 6644 27124
rect 6503 27084 6644 27112
rect 6503 27081 6515 27084
rect 6457 27075 6515 27081
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 6822 27072 6828 27124
rect 6880 27072 6886 27124
rect 9309 27115 9367 27121
rect 9309 27081 9321 27115
rect 9355 27112 9367 27115
rect 11514 27112 11520 27124
rect 9355 27084 11520 27112
rect 9355 27081 9367 27084
rect 9309 27075 9367 27081
rect 11514 27072 11520 27084
rect 11572 27072 11578 27124
rect 5997 27047 6055 27053
rect 5997 27013 6009 27047
rect 6043 27044 6055 27047
rect 6840 27044 6868 27072
rect 6043 27016 6868 27044
rect 6043 27013 6055 27016
rect 5997 27007 6055 27013
rect 3789 26979 3847 26985
rect 3789 26945 3801 26979
rect 3835 26976 3847 26979
rect 4154 26976 4160 26988
rect 3835 26948 4160 26976
rect 3835 26945 3847 26948
rect 3789 26939 3847 26945
rect 4154 26936 4160 26948
rect 4212 26976 4218 26988
rect 4249 26979 4307 26985
rect 4249 26976 4261 26979
rect 4212 26948 4261 26976
rect 4212 26936 4218 26948
rect 4249 26945 4261 26948
rect 4295 26945 4307 26979
rect 4249 26939 4307 26945
rect 6178 26936 6184 26988
rect 6236 26936 6242 26988
rect 10778 26936 10784 26988
rect 10836 26976 10842 26988
rect 10873 26979 10931 26985
rect 10873 26976 10885 26979
rect 10836 26948 10885 26976
rect 10836 26936 10842 26948
rect 10873 26945 10885 26948
rect 10919 26945 10931 26979
rect 10873 26939 10931 26945
rect 10962 26936 10968 26988
rect 11020 26976 11026 26988
rect 11020 26948 11065 26976
rect 11020 26936 11026 26948
rect 5994 26868 6000 26920
rect 6052 26908 6058 26920
rect 6196 26908 6224 26936
rect 6052 26880 6224 26908
rect 6365 26911 6423 26917
rect 6052 26868 6058 26880
rect 6365 26877 6377 26911
rect 6411 26908 6423 26911
rect 6641 26911 6699 26917
rect 6641 26908 6653 26911
rect 6411 26880 6653 26908
rect 6411 26877 6423 26880
rect 6365 26871 6423 26877
rect 6641 26877 6653 26880
rect 6687 26908 6699 26911
rect 6822 26908 6828 26920
rect 6687 26880 6828 26908
rect 6687 26877 6699 26880
rect 6641 26871 6699 26877
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 7466 26908 7472 26920
rect 7427 26880 7472 26908
rect 7466 26868 7472 26880
rect 7524 26868 7530 26920
rect 12802 26868 12808 26920
rect 12860 26908 12866 26920
rect 13354 26908 13360 26920
rect 12860 26880 13360 26908
rect 12860 26868 12866 26880
rect 13354 26868 13360 26880
rect 13412 26868 13418 26920
rect 4157 26843 4215 26849
rect 4157 26809 4169 26843
rect 4203 26840 4215 26843
rect 4516 26843 4574 26849
rect 4516 26840 4528 26843
rect 4203 26812 4528 26840
rect 4203 26809 4215 26812
rect 4157 26803 4215 26809
rect 4516 26809 4528 26812
rect 4562 26840 4574 26843
rect 4890 26840 4896 26852
rect 4562 26812 4896 26840
rect 4562 26809 4574 26812
rect 4516 26803 4574 26809
rect 4890 26800 4896 26812
rect 4948 26800 4954 26852
rect 5810 26800 5816 26852
rect 5868 26840 5874 26852
rect 6546 26840 6552 26852
rect 5868 26812 6552 26840
rect 5868 26800 5874 26812
rect 6546 26800 6552 26812
rect 6604 26800 6610 26852
rect 7714 26843 7772 26849
rect 7714 26840 7726 26843
rect 7300 26812 7726 26840
rect 7300 26784 7328 26812
rect 7714 26809 7726 26812
rect 7760 26809 7772 26843
rect 7714 26803 7772 26809
rect 10686 26800 10692 26852
rect 10744 26840 10750 26852
rect 10781 26843 10839 26849
rect 10781 26840 10793 26843
rect 10744 26812 10793 26840
rect 10744 26800 10750 26812
rect 10781 26809 10793 26812
rect 10827 26809 10839 26843
rect 10781 26803 10839 26809
rect 7282 26772 7288 26784
rect 7243 26744 7288 26772
rect 7282 26732 7288 26744
rect 7340 26732 7346 26784
rect 8754 26732 8760 26784
rect 8812 26772 8818 26784
rect 8849 26775 8907 26781
rect 8849 26772 8861 26775
rect 8812 26744 8861 26772
rect 8812 26732 8818 26744
rect 8849 26741 8861 26744
rect 8895 26741 8907 26775
rect 8849 26735 8907 26741
rect 9677 26775 9735 26781
rect 9677 26741 9689 26775
rect 9723 26772 9735 26775
rect 9766 26772 9772 26784
rect 9723 26744 9772 26772
rect 9723 26741 9735 26744
rect 9677 26735 9735 26741
rect 9766 26732 9772 26744
rect 9824 26732 9830 26784
rect 10042 26772 10048 26784
rect 10003 26744 10048 26772
rect 10042 26732 10048 26744
rect 10100 26772 10106 26784
rect 10226 26772 10232 26784
rect 10100 26744 10232 26772
rect 10100 26732 10106 26744
rect 10226 26732 10232 26744
rect 10284 26732 10290 26784
rect 10410 26772 10416 26784
rect 10371 26744 10416 26772
rect 10410 26732 10416 26744
rect 10468 26732 10474 26784
rect 11422 26732 11428 26784
rect 11480 26772 11486 26784
rect 11885 26775 11943 26781
rect 11885 26772 11897 26775
rect 11480 26744 11897 26772
rect 11480 26732 11486 26744
rect 11885 26741 11897 26744
rect 11931 26741 11943 26775
rect 11885 26735 11943 26741
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 4062 26568 4068 26580
rect 4023 26540 4068 26568
rect 4062 26528 4068 26540
rect 4120 26528 4126 26580
rect 5350 26528 5356 26580
rect 5408 26568 5414 26580
rect 5537 26571 5595 26577
rect 5537 26568 5549 26571
rect 5408 26540 5549 26568
rect 5408 26528 5414 26540
rect 5537 26537 5549 26540
rect 5583 26568 5595 26571
rect 5626 26568 5632 26580
rect 5583 26540 5632 26568
rect 5583 26537 5595 26540
rect 5537 26531 5595 26537
rect 5626 26528 5632 26540
rect 5684 26528 5690 26580
rect 9674 26528 9680 26580
rect 9732 26568 9738 26580
rect 10137 26571 10195 26577
rect 10137 26568 10149 26571
rect 9732 26540 10149 26568
rect 9732 26528 9738 26540
rect 10137 26537 10149 26540
rect 10183 26537 10195 26571
rect 10137 26531 10195 26537
rect 10686 26528 10692 26580
rect 10744 26568 10750 26580
rect 11057 26571 11115 26577
rect 11057 26568 11069 26571
rect 10744 26540 11069 26568
rect 10744 26528 10750 26540
rect 11057 26537 11069 26540
rect 11103 26537 11115 26571
rect 11057 26531 11115 26537
rect 1670 26500 1676 26512
rect 1631 26472 1676 26500
rect 1670 26460 1676 26472
rect 1728 26460 1734 26512
rect 4433 26503 4491 26509
rect 4433 26469 4445 26503
rect 4479 26500 4491 26503
rect 4522 26500 4528 26512
rect 4479 26472 4528 26500
rect 4479 26469 4491 26472
rect 4433 26463 4491 26469
rect 4522 26460 4528 26472
rect 4580 26460 4586 26512
rect 6172 26503 6230 26509
rect 6172 26469 6184 26503
rect 6218 26500 6230 26503
rect 6270 26500 6276 26512
rect 6218 26472 6276 26500
rect 6218 26469 6230 26472
rect 6172 26463 6230 26469
rect 6270 26460 6276 26472
rect 6328 26500 6334 26512
rect 6730 26500 6736 26512
rect 6328 26472 6736 26500
rect 6328 26460 6334 26472
rect 6730 26460 6736 26472
rect 6788 26460 6794 26512
rect 10781 26503 10839 26509
rect 10781 26469 10793 26503
rect 10827 26500 10839 26503
rect 10962 26500 10968 26512
rect 10827 26472 10968 26500
rect 10827 26469 10839 26472
rect 10781 26463 10839 26469
rect 10962 26460 10968 26472
rect 11020 26460 11026 26512
rect 1397 26435 1455 26441
rect 1397 26401 1409 26435
rect 1443 26432 1455 26435
rect 1486 26432 1492 26444
rect 1443 26404 1492 26432
rect 1443 26401 1455 26404
rect 1397 26395 1455 26401
rect 1486 26392 1492 26404
rect 1544 26392 1550 26444
rect 7466 26432 7472 26444
rect 5920 26404 7472 26432
rect 5920 26376 5948 26404
rect 7466 26392 7472 26404
rect 7524 26432 7530 26444
rect 7929 26435 7987 26441
rect 7929 26432 7941 26435
rect 7524 26404 7941 26432
rect 7524 26392 7530 26404
rect 7929 26401 7941 26404
rect 7975 26401 7987 26435
rect 10042 26432 10048 26444
rect 10003 26404 10048 26432
rect 7929 26395 7987 26401
rect 10042 26392 10048 26404
rect 10100 26392 10106 26444
rect 4430 26324 4436 26376
rect 4488 26364 4494 26376
rect 4525 26367 4583 26373
rect 4525 26364 4537 26367
rect 4488 26336 4537 26364
rect 4488 26324 4494 26336
rect 4525 26333 4537 26336
rect 4571 26333 4583 26367
rect 4525 26327 4583 26333
rect 4709 26367 4767 26373
rect 4709 26333 4721 26367
rect 4755 26364 4767 26367
rect 4890 26364 4896 26376
rect 4755 26336 4896 26364
rect 4755 26333 4767 26336
rect 4709 26327 4767 26333
rect 4890 26324 4896 26336
rect 4948 26324 4954 26376
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26364 5319 26367
rect 5534 26364 5540 26376
rect 5307 26336 5540 26364
rect 5307 26333 5319 26336
rect 5261 26327 5319 26333
rect 5534 26324 5540 26336
rect 5592 26324 5598 26376
rect 5902 26364 5908 26376
rect 5863 26336 5908 26364
rect 5902 26324 5908 26336
rect 5960 26324 5966 26376
rect 9490 26324 9496 26376
rect 9548 26364 9554 26376
rect 10321 26367 10379 26373
rect 10321 26364 10333 26367
rect 9548 26336 10333 26364
rect 9548 26324 9554 26336
rect 10321 26333 10333 26336
rect 10367 26364 10379 26367
rect 10594 26364 10600 26376
rect 10367 26336 10600 26364
rect 10367 26333 10379 26336
rect 10321 26327 10379 26333
rect 10594 26324 10600 26336
rect 10652 26324 10658 26376
rect 5552 26296 5580 26324
rect 7282 26296 7288 26308
rect 5552 26268 5672 26296
rect 5644 26228 5672 26268
rect 6840 26268 7288 26296
rect 6840 26228 6868 26268
rect 7282 26256 7288 26268
rect 7340 26256 7346 26308
rect 9674 26296 9680 26308
rect 9635 26268 9680 26296
rect 9674 26256 9680 26268
rect 9732 26256 9738 26308
rect 5644 26200 6868 26228
rect 7190 26188 7196 26240
rect 7248 26228 7254 26240
rect 7561 26231 7619 26237
rect 7561 26228 7573 26231
rect 7248 26200 7573 26228
rect 7248 26188 7254 26200
rect 7561 26197 7573 26200
rect 7607 26197 7619 26231
rect 7561 26191 7619 26197
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 4157 26027 4215 26033
rect 4157 25993 4169 26027
rect 4203 26024 4215 26027
rect 4430 26024 4436 26036
rect 4203 25996 4436 26024
rect 4203 25993 4215 25996
rect 4157 25987 4215 25993
rect 4430 25984 4436 25996
rect 4488 25984 4494 26036
rect 6270 26024 6276 26036
rect 6231 25996 6276 26024
rect 6270 25984 6276 25996
rect 6328 25984 6334 26036
rect 6638 26024 6644 26036
rect 6599 25996 6644 26024
rect 6638 25984 6644 25996
rect 6696 25984 6702 26036
rect 7098 25984 7104 26036
rect 7156 26024 7162 26036
rect 7282 26024 7288 26036
rect 7156 25996 7288 26024
rect 7156 25984 7162 25996
rect 7282 25984 7288 25996
rect 7340 25984 7346 26036
rect 7469 26027 7527 26033
rect 7469 25993 7481 26027
rect 7515 26024 7527 26027
rect 7558 26024 7564 26036
rect 7515 25996 7564 26024
rect 7515 25993 7527 25996
rect 7469 25987 7527 25993
rect 7558 25984 7564 25996
rect 7616 25984 7622 26036
rect 9217 26027 9275 26033
rect 9217 25993 9229 26027
rect 9263 26024 9275 26027
rect 10226 26024 10232 26036
rect 9263 25996 10232 26024
rect 9263 25993 9275 25996
rect 9217 25987 9275 25993
rect 1486 25916 1492 25968
rect 1544 25956 1550 25968
rect 2225 25959 2283 25965
rect 2225 25956 2237 25959
rect 1544 25928 2237 25956
rect 1544 25916 1550 25928
rect 2225 25925 2237 25928
rect 2271 25956 2283 25959
rect 5169 25959 5227 25965
rect 5169 25956 5181 25959
rect 2271 25928 5181 25956
rect 2271 25925 2283 25928
rect 2225 25919 2283 25925
rect 5169 25925 5181 25928
rect 5215 25925 5227 25959
rect 5169 25919 5227 25925
rect 9033 25959 9091 25965
rect 9033 25925 9045 25959
rect 9079 25956 9091 25959
rect 9490 25956 9496 25968
rect 9079 25928 9496 25956
rect 9079 25925 9091 25928
rect 9033 25919 9091 25925
rect 9490 25916 9496 25928
rect 9548 25916 9554 25968
rect 9674 25916 9680 25968
rect 9732 25956 9738 25968
rect 10042 25956 10048 25968
rect 9732 25928 10048 25956
rect 9732 25916 9738 25928
rect 10042 25916 10048 25928
rect 10100 25916 10106 25968
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 5534 25848 5540 25900
rect 5592 25888 5598 25900
rect 5721 25891 5779 25897
rect 5721 25888 5733 25891
rect 5592 25860 5733 25888
rect 5592 25848 5598 25860
rect 5721 25857 5733 25860
rect 5767 25857 5779 25891
rect 10152 25888 10180 25996
rect 10226 25984 10232 25996
rect 10284 25984 10290 26036
rect 11241 26027 11299 26033
rect 11241 25993 11253 26027
rect 11287 26024 11299 26027
rect 11514 26024 11520 26036
rect 11287 25996 11520 26024
rect 11287 25993 11299 25996
rect 11241 25987 11299 25993
rect 5721 25851 5779 25857
rect 9968 25860 10180 25888
rect 10781 25891 10839 25897
rect 1397 25823 1455 25829
rect 1397 25789 1409 25823
rect 1443 25820 1455 25823
rect 5626 25820 5632 25832
rect 1443 25792 2544 25820
rect 5587 25792 5632 25820
rect 1443 25789 1455 25792
rect 1397 25783 1455 25789
rect 2516 25696 2544 25792
rect 5626 25780 5632 25792
rect 5684 25780 5690 25832
rect 4522 25752 4528 25764
rect 4483 25724 4528 25752
rect 4522 25712 4528 25724
rect 4580 25712 4586 25764
rect 5534 25752 5540 25764
rect 5495 25724 5540 25752
rect 5534 25712 5540 25724
rect 5592 25712 5598 25764
rect 9968 25752 9996 25860
rect 10781 25857 10793 25891
rect 10827 25888 10839 25891
rect 11256 25888 11284 25987
rect 11514 25984 11520 25996
rect 11572 25984 11578 26036
rect 10827 25860 11284 25888
rect 10827 25857 10839 25860
rect 10781 25851 10839 25857
rect 10045 25823 10103 25829
rect 10045 25789 10057 25823
rect 10091 25820 10103 25823
rect 10502 25820 10508 25832
rect 10091 25792 10508 25820
rect 10091 25789 10103 25792
rect 10045 25783 10103 25789
rect 10502 25780 10508 25792
rect 10560 25820 10566 25832
rect 11517 25823 11575 25829
rect 11517 25820 11529 25823
rect 10560 25792 11529 25820
rect 10560 25780 10566 25792
rect 11517 25789 11529 25792
rect 11563 25789 11575 25823
rect 11517 25783 11575 25789
rect 9968 25724 10548 25752
rect 2498 25684 2504 25696
rect 2459 25656 2504 25684
rect 2498 25644 2504 25656
rect 2556 25644 2562 25696
rect 4890 25684 4896 25696
rect 4851 25656 4896 25684
rect 4890 25644 4896 25656
rect 4948 25644 4954 25696
rect 5074 25644 5080 25696
rect 5132 25684 5138 25696
rect 5626 25684 5632 25696
rect 5132 25656 5632 25684
rect 5132 25644 5138 25656
rect 5626 25644 5632 25656
rect 5684 25644 5690 25696
rect 7650 25644 7656 25696
rect 7708 25684 7714 25696
rect 9217 25687 9275 25693
rect 9217 25684 9229 25687
rect 7708 25656 9229 25684
rect 7708 25644 7714 25656
rect 9217 25653 9229 25656
rect 9263 25684 9275 25687
rect 9309 25687 9367 25693
rect 9309 25684 9321 25687
rect 9263 25656 9321 25684
rect 9263 25653 9275 25656
rect 9217 25647 9275 25653
rect 9309 25653 9321 25656
rect 9355 25653 9367 25687
rect 9674 25684 9680 25696
rect 9635 25656 9680 25684
rect 9309 25647 9367 25653
rect 9674 25644 9680 25656
rect 9732 25644 9738 25696
rect 9858 25684 9864 25696
rect 9819 25656 9864 25684
rect 9858 25644 9864 25656
rect 9916 25644 9922 25696
rect 10134 25684 10140 25696
rect 10095 25656 10140 25684
rect 10134 25644 10140 25656
rect 10192 25644 10198 25696
rect 10520 25693 10548 25724
rect 10505 25687 10563 25693
rect 10505 25653 10517 25687
rect 10551 25653 10563 25687
rect 10505 25647 10563 25653
rect 10594 25644 10600 25696
rect 10652 25684 10658 25696
rect 10652 25656 10697 25684
rect 10652 25644 10658 25656
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 4890 25440 4896 25492
rect 4948 25480 4954 25492
rect 5445 25483 5503 25489
rect 5445 25480 5457 25483
rect 4948 25452 5457 25480
rect 4948 25440 4954 25452
rect 5445 25449 5457 25452
rect 5491 25449 5503 25483
rect 5445 25443 5503 25449
rect 5534 25440 5540 25492
rect 5592 25480 5598 25492
rect 5721 25483 5779 25489
rect 5721 25480 5733 25483
rect 5592 25452 5733 25480
rect 5592 25440 5598 25452
rect 5721 25449 5733 25452
rect 5767 25449 5779 25483
rect 5721 25443 5779 25449
rect 9493 25483 9551 25489
rect 9493 25449 9505 25483
rect 9539 25480 9551 25483
rect 9582 25480 9588 25492
rect 9539 25452 9588 25480
rect 9539 25449 9551 25452
rect 9493 25443 9551 25449
rect 9582 25440 9588 25452
rect 9640 25440 9646 25492
rect 10594 25480 10600 25492
rect 10152 25452 10600 25480
rect 10042 25372 10048 25424
rect 10100 25412 10106 25424
rect 10152 25421 10180 25452
rect 10594 25440 10600 25452
rect 10652 25440 10658 25492
rect 12618 25480 12624 25492
rect 12579 25452 12624 25480
rect 12618 25440 12624 25452
rect 12676 25440 12682 25492
rect 12894 25440 12900 25492
rect 12952 25480 12958 25492
rect 13173 25483 13231 25489
rect 13173 25480 13185 25483
rect 12952 25452 13185 25480
rect 12952 25440 12958 25452
rect 13173 25449 13185 25452
rect 13219 25449 13231 25483
rect 13173 25443 13231 25449
rect 10137 25415 10195 25421
rect 10137 25412 10149 25415
rect 10100 25384 10149 25412
rect 10100 25372 10106 25384
rect 10137 25381 10149 25384
rect 10183 25381 10195 25415
rect 10137 25375 10195 25381
rect 1394 25344 1400 25356
rect 1355 25316 1400 25344
rect 1394 25304 1400 25316
rect 1452 25304 1458 25356
rect 4154 25304 4160 25356
rect 4212 25344 4218 25356
rect 4321 25347 4379 25353
rect 4321 25344 4333 25347
rect 4212 25316 4333 25344
rect 4212 25304 4218 25316
rect 4321 25313 4333 25316
rect 4367 25313 4379 25347
rect 4321 25307 4379 25313
rect 6457 25347 6515 25353
rect 6457 25313 6469 25347
rect 6503 25344 6515 25347
rect 6638 25344 6644 25356
rect 6503 25316 6644 25344
rect 6503 25313 6515 25316
rect 6457 25307 6515 25313
rect 6638 25304 6644 25316
rect 6696 25304 6702 25356
rect 10594 25304 10600 25356
rect 10652 25344 10658 25356
rect 10965 25347 11023 25353
rect 10965 25344 10977 25347
rect 10652 25316 10977 25344
rect 10652 25304 10658 25316
rect 10965 25313 10977 25316
rect 11011 25344 11023 25347
rect 11609 25347 11667 25353
rect 11609 25344 11621 25347
rect 11011 25316 11621 25344
rect 11011 25313 11023 25316
rect 10965 25307 11023 25313
rect 11609 25313 11621 25316
rect 11655 25313 11667 25347
rect 12526 25344 12532 25356
rect 12487 25316 12532 25344
rect 11609 25307 11667 25313
rect 12526 25304 12532 25316
rect 12584 25304 12590 25356
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 4062 25276 4068 25288
rect 4023 25248 4068 25276
rect 4062 25236 4068 25248
rect 4120 25236 4126 25288
rect 10042 25236 10048 25288
rect 10100 25276 10106 25288
rect 10410 25276 10416 25288
rect 10100 25248 10416 25276
rect 10100 25236 10106 25248
rect 10410 25236 10416 25248
rect 10468 25276 10474 25288
rect 11057 25279 11115 25285
rect 11057 25276 11069 25279
rect 10468 25248 11069 25276
rect 10468 25236 10474 25248
rect 11057 25245 11069 25248
rect 11103 25245 11115 25279
rect 11057 25239 11115 25245
rect 11149 25279 11207 25285
rect 11149 25245 11161 25279
rect 11195 25245 11207 25279
rect 11149 25239 11207 25245
rect 12805 25279 12863 25285
rect 12805 25245 12817 25279
rect 12851 25276 12863 25279
rect 12894 25276 12900 25288
rect 12851 25248 12900 25276
rect 12851 25245 12863 25248
rect 12805 25239 12863 25245
rect 9490 25168 9496 25220
rect 9548 25208 9554 25220
rect 10597 25211 10655 25217
rect 10597 25208 10609 25211
rect 9548 25180 10609 25208
rect 9548 25168 9554 25180
rect 10597 25177 10609 25180
rect 10643 25177 10655 25211
rect 10597 25171 10655 25177
rect 10778 25168 10784 25220
rect 10836 25208 10842 25220
rect 11164 25208 11192 25239
rect 12894 25236 12900 25248
rect 12952 25236 12958 25288
rect 10836 25180 11192 25208
rect 10836 25168 10842 25180
rect 5902 25100 5908 25152
rect 5960 25140 5966 25152
rect 6181 25143 6239 25149
rect 6181 25140 6193 25143
rect 5960 25112 6193 25140
rect 5960 25100 5966 25112
rect 6181 25109 6193 25112
rect 6227 25140 6239 25143
rect 6273 25143 6331 25149
rect 6273 25140 6285 25143
rect 6227 25112 6285 25140
rect 6227 25109 6239 25112
rect 6181 25103 6239 25109
rect 6273 25109 6285 25112
rect 6319 25140 6331 25143
rect 6730 25140 6736 25152
rect 6319 25112 6736 25140
rect 6319 25109 6331 25112
rect 6273 25103 6331 25109
rect 6730 25100 6736 25112
rect 6788 25100 6794 25152
rect 7190 25140 7196 25152
rect 7151 25112 7196 25140
rect 7190 25100 7196 25112
rect 7248 25100 7254 25152
rect 7466 25140 7472 25152
rect 7427 25112 7472 25140
rect 7466 25100 7472 25112
rect 7524 25100 7530 25152
rect 9125 25143 9183 25149
rect 9125 25109 9137 25143
rect 9171 25140 9183 25143
rect 9582 25140 9588 25152
rect 9171 25112 9588 25140
rect 9171 25109 9183 25112
rect 9125 25103 9183 25109
rect 9582 25100 9588 25112
rect 9640 25100 9646 25152
rect 12161 25143 12219 25149
rect 12161 25109 12173 25143
rect 12207 25140 12219 25143
rect 12342 25140 12348 25152
rect 12207 25112 12348 25140
rect 12207 25109 12219 25112
rect 12161 25103 12219 25109
rect 12342 25100 12348 25112
rect 12400 25100 12406 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 1394 24896 1400 24948
rect 1452 24936 1458 24948
rect 1581 24939 1639 24945
rect 1581 24936 1593 24939
rect 1452 24908 1593 24936
rect 1452 24896 1458 24908
rect 1581 24905 1593 24908
rect 1627 24905 1639 24939
rect 1581 24899 1639 24905
rect 6273 24939 6331 24945
rect 6273 24905 6285 24939
rect 6319 24936 6331 24939
rect 6638 24936 6644 24948
rect 6319 24908 6644 24936
rect 6319 24905 6331 24908
rect 6273 24899 6331 24905
rect 6638 24896 6644 24908
rect 6696 24896 6702 24948
rect 10594 24936 10600 24948
rect 10555 24908 10600 24936
rect 10594 24896 10600 24908
rect 10652 24896 10658 24948
rect 12526 24896 12532 24948
rect 12584 24936 12590 24948
rect 13170 24936 13176 24948
rect 12584 24908 13176 24936
rect 12584 24896 12590 24908
rect 13170 24896 13176 24908
rect 13228 24936 13234 24948
rect 13449 24939 13507 24945
rect 13449 24936 13461 24939
rect 13228 24908 13461 24936
rect 13228 24896 13234 24908
rect 13449 24905 13461 24908
rect 13495 24905 13507 24939
rect 13449 24899 13507 24905
rect 7190 24828 7196 24880
rect 7248 24868 7254 24880
rect 7248 24840 7788 24868
rect 7248 24828 7254 24840
rect 4617 24803 4675 24809
rect 4617 24769 4629 24803
rect 4663 24800 4675 24803
rect 5721 24803 5779 24809
rect 5721 24800 5733 24803
rect 4663 24772 5733 24800
rect 4663 24769 4675 24772
rect 4617 24763 4675 24769
rect 5721 24769 5733 24772
rect 5767 24800 5779 24803
rect 5902 24800 5908 24812
rect 5767 24772 5908 24800
rect 5767 24769 5779 24772
rect 5721 24763 5779 24769
rect 5902 24760 5908 24772
rect 5960 24760 5966 24812
rect 7760 24809 7788 24840
rect 12894 24828 12900 24880
rect 12952 24868 12958 24880
rect 12952 24840 13032 24868
rect 12952 24828 12958 24840
rect 7745 24803 7803 24809
rect 7745 24769 7757 24803
rect 7791 24800 7803 24803
rect 8294 24800 8300 24812
rect 7791 24772 8300 24800
rect 7791 24769 7803 24772
rect 7745 24763 7803 24769
rect 8294 24760 8300 24772
rect 8352 24760 8358 24812
rect 9490 24800 9496 24812
rect 9451 24772 9496 24800
rect 9490 24760 9496 24772
rect 9548 24760 9554 24812
rect 9585 24803 9643 24809
rect 9585 24769 9597 24803
rect 9631 24769 9643 24803
rect 9585 24763 9643 24769
rect 4985 24735 5043 24741
rect 4985 24701 4997 24735
rect 5031 24732 5043 24735
rect 5258 24732 5264 24744
rect 5031 24704 5264 24732
rect 5031 24701 5043 24704
rect 4985 24695 5043 24701
rect 5258 24692 5264 24704
rect 5316 24732 5322 24744
rect 5442 24732 5448 24744
rect 5316 24704 5448 24732
rect 5316 24692 5322 24704
rect 5442 24692 5448 24704
rect 5500 24732 5506 24744
rect 5537 24735 5595 24741
rect 5537 24732 5549 24735
rect 5500 24704 5549 24732
rect 5500 24692 5506 24704
rect 5537 24701 5549 24704
rect 5583 24701 5595 24735
rect 5537 24695 5595 24701
rect 6914 24692 6920 24744
rect 6972 24732 6978 24744
rect 7466 24732 7472 24744
rect 6972 24704 7472 24732
rect 6972 24692 6978 24704
rect 7466 24692 7472 24704
rect 7524 24692 7530 24744
rect 8941 24735 8999 24741
rect 8941 24701 8953 24735
rect 8987 24732 8999 24735
rect 9306 24732 9312 24744
rect 8987 24704 9312 24732
rect 8987 24701 8999 24704
rect 8941 24695 8999 24701
rect 9306 24692 9312 24704
rect 9364 24732 9370 24744
rect 9600 24732 9628 24763
rect 10134 24760 10140 24812
rect 10192 24800 10198 24812
rect 13004 24809 13032 24840
rect 11057 24803 11115 24809
rect 11057 24800 11069 24803
rect 10192 24772 11069 24800
rect 10192 24760 10198 24772
rect 11057 24769 11069 24772
rect 11103 24769 11115 24803
rect 11057 24763 11115 24769
rect 11149 24803 11207 24809
rect 11149 24769 11161 24803
rect 11195 24800 11207 24803
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 11195 24772 13001 24800
rect 11195 24769 11207 24772
rect 11149 24763 11207 24769
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 9364 24704 9628 24732
rect 9364 24692 9370 24704
rect 10226 24692 10232 24744
rect 10284 24732 10290 24744
rect 10410 24732 10416 24744
rect 10284 24704 10416 24732
rect 10284 24692 10290 24704
rect 10410 24692 10416 24704
rect 10468 24732 10474 24744
rect 10468 24704 10916 24732
rect 10468 24692 10474 24704
rect 4062 24664 4068 24676
rect 3712 24636 4068 24664
rect 3142 24556 3148 24608
rect 3200 24596 3206 24608
rect 3712 24605 3740 24636
rect 4062 24624 4068 24636
rect 4120 24624 4126 24676
rect 6641 24667 6699 24673
rect 6641 24633 6653 24667
rect 6687 24664 6699 24667
rect 7006 24664 7012 24676
rect 6687 24636 7012 24664
rect 6687 24633 6699 24636
rect 6641 24627 6699 24633
rect 7006 24624 7012 24636
rect 7064 24664 7070 24676
rect 7561 24667 7619 24673
rect 7561 24664 7573 24667
rect 7064 24636 7573 24664
rect 7064 24624 7070 24636
rect 7561 24633 7573 24636
rect 7607 24633 7619 24667
rect 10778 24664 10784 24676
rect 7561 24627 7619 24633
rect 10060 24636 10784 24664
rect 3697 24599 3755 24605
rect 3697 24596 3709 24599
rect 3200 24568 3709 24596
rect 3200 24556 3206 24568
rect 3697 24565 3709 24568
rect 3743 24565 3755 24599
rect 4154 24596 4160 24608
rect 4115 24568 4160 24596
rect 3697 24559 3755 24565
rect 4154 24556 4160 24568
rect 4212 24556 4218 24608
rect 5074 24596 5080 24608
rect 5035 24568 5080 24596
rect 5074 24556 5080 24568
rect 5132 24556 5138 24608
rect 5166 24556 5172 24608
rect 5224 24596 5230 24608
rect 5445 24599 5503 24605
rect 5445 24596 5457 24599
rect 5224 24568 5457 24596
rect 5224 24556 5230 24568
rect 5445 24565 5457 24568
rect 5491 24565 5503 24599
rect 7098 24596 7104 24608
rect 7059 24568 7104 24596
rect 5445 24559 5503 24565
rect 7098 24556 7104 24568
rect 7156 24556 7162 24608
rect 9030 24596 9036 24608
rect 8991 24568 9036 24596
rect 9030 24556 9036 24568
rect 9088 24556 9094 24608
rect 9401 24599 9459 24605
rect 9401 24565 9413 24599
rect 9447 24596 9459 24599
rect 9582 24596 9588 24608
rect 9447 24568 9588 24596
rect 9447 24565 9459 24568
rect 9401 24559 9459 24565
rect 9582 24556 9588 24568
rect 9640 24556 9646 24608
rect 9858 24556 9864 24608
rect 9916 24596 9922 24608
rect 10060 24605 10088 24636
rect 10778 24624 10784 24636
rect 10836 24624 10842 24676
rect 10045 24599 10103 24605
rect 10045 24596 10057 24599
rect 9916 24568 10057 24596
rect 9916 24556 9922 24568
rect 10045 24565 10057 24568
rect 10091 24565 10103 24599
rect 10888 24596 10916 24704
rect 10962 24692 10968 24744
rect 11020 24732 11026 24744
rect 11164 24732 11192 24763
rect 12897 24735 12955 24741
rect 12897 24732 12909 24735
rect 11020 24704 11192 24732
rect 11992 24704 12909 24732
rect 11020 24692 11026 24704
rect 11992 24608 12020 24704
rect 12897 24701 12909 24704
rect 12943 24701 12955 24735
rect 12897 24695 12955 24701
rect 12158 24664 12164 24676
rect 12119 24636 12164 24664
rect 12158 24624 12164 24636
rect 12216 24664 12222 24676
rect 12216 24636 12848 24664
rect 12216 24624 12222 24636
rect 10965 24599 11023 24605
rect 10965 24596 10977 24599
rect 10888 24568 10977 24596
rect 10045 24559 10103 24565
rect 10965 24565 10977 24568
rect 11011 24565 11023 24599
rect 10965 24559 11023 24565
rect 11885 24599 11943 24605
rect 11885 24565 11897 24599
rect 11931 24596 11943 24599
rect 11974 24596 11980 24608
rect 11931 24568 11980 24596
rect 11931 24565 11943 24568
rect 11885 24559 11943 24565
rect 11974 24556 11980 24568
rect 12032 24556 12038 24608
rect 12437 24599 12495 24605
rect 12437 24565 12449 24599
rect 12483 24596 12495 24599
rect 12618 24596 12624 24608
rect 12483 24568 12624 24596
rect 12483 24565 12495 24568
rect 12437 24559 12495 24565
rect 12618 24556 12624 24568
rect 12676 24556 12682 24608
rect 12820 24605 12848 24636
rect 12805 24599 12863 24605
rect 12805 24565 12817 24599
rect 12851 24596 12863 24599
rect 12986 24596 12992 24608
rect 12851 24568 12992 24596
rect 12851 24565 12863 24568
rect 12805 24559 12863 24565
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 5166 24392 5172 24404
rect 5127 24364 5172 24392
rect 5166 24352 5172 24364
rect 5224 24352 5230 24404
rect 5721 24395 5779 24401
rect 5721 24361 5733 24395
rect 5767 24392 5779 24395
rect 5994 24392 6000 24404
rect 5767 24364 6000 24392
rect 5767 24361 5779 24364
rect 5721 24355 5779 24361
rect 5994 24352 6000 24364
rect 6052 24352 6058 24404
rect 8294 24392 8300 24404
rect 8255 24364 8300 24392
rect 8294 24352 8300 24364
rect 8352 24352 8358 24404
rect 9125 24395 9183 24401
rect 9125 24361 9137 24395
rect 9171 24392 9183 24395
rect 9490 24392 9496 24404
rect 9171 24364 9496 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 9490 24352 9496 24364
rect 9548 24352 9554 24404
rect 9953 24395 10011 24401
rect 9953 24361 9965 24395
rect 9999 24392 10011 24395
rect 10042 24392 10048 24404
rect 9999 24364 10048 24392
rect 9999 24361 10011 24364
rect 9953 24355 10011 24361
rect 10042 24352 10048 24364
rect 10100 24352 10106 24404
rect 10134 24352 10140 24404
rect 10192 24392 10198 24404
rect 10229 24395 10287 24401
rect 10229 24392 10241 24395
rect 10192 24364 10241 24392
rect 10192 24352 10198 24364
rect 10229 24361 10241 24364
rect 10275 24361 10287 24395
rect 10229 24355 10287 24361
rect 10689 24395 10747 24401
rect 10689 24361 10701 24395
rect 10735 24392 10747 24395
rect 10962 24392 10968 24404
rect 10735 24364 10968 24392
rect 10735 24361 10747 24364
rect 10689 24355 10747 24361
rect 10962 24352 10968 24364
rect 11020 24352 11026 24404
rect 12710 24392 12716 24404
rect 12671 24364 12716 24392
rect 12710 24352 12716 24364
rect 12768 24392 12774 24404
rect 12768 24364 12848 24392
rect 12768 24352 12774 24364
rect 10980 24324 11008 24352
rect 11210 24327 11268 24333
rect 11210 24324 11222 24327
rect 10980 24296 11222 24324
rect 11210 24293 11222 24296
rect 11256 24293 11268 24327
rect 11210 24287 11268 24293
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6086 24256 6092 24268
rect 5859 24228 6092 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 6086 24216 6092 24228
rect 6144 24216 6150 24268
rect 7190 24265 7196 24268
rect 7184 24256 7196 24265
rect 7151 24228 7196 24256
rect 7184 24219 7196 24228
rect 7190 24216 7196 24219
rect 7248 24216 7254 24268
rect 10686 24216 10692 24268
rect 10744 24256 10750 24268
rect 10965 24259 11023 24265
rect 10965 24256 10977 24259
rect 10744 24228 10977 24256
rect 10744 24216 10750 24228
rect 10965 24225 10977 24228
rect 11011 24225 11023 24259
rect 12820 24256 12848 24364
rect 12894 24352 12900 24404
rect 12952 24392 12958 24404
rect 12989 24395 13047 24401
rect 12989 24392 13001 24395
rect 12952 24364 13001 24392
rect 12952 24352 12958 24364
rect 12989 24361 13001 24364
rect 13035 24361 13047 24395
rect 13170 24392 13176 24404
rect 13131 24364 13176 24392
rect 12989 24355 13047 24361
rect 13170 24352 13176 24364
rect 13228 24352 13234 24404
rect 13170 24256 13176 24268
rect 12820 24228 13176 24256
rect 10965 24219 11023 24225
rect 13170 24216 13176 24228
rect 13228 24216 13234 24268
rect 5902 24188 5908 24200
rect 5863 24160 5908 24188
rect 5902 24148 5908 24160
rect 5960 24148 5966 24200
rect 6917 24191 6975 24197
rect 6917 24188 6929 24191
rect 6748 24160 6929 24188
rect 6748 24064 6776 24160
rect 6917 24157 6929 24160
rect 6963 24157 6975 24191
rect 6917 24151 6975 24157
rect 3142 24052 3148 24064
rect 3103 24024 3148 24052
rect 3142 24012 3148 24024
rect 3200 24012 3206 24064
rect 5350 24052 5356 24064
rect 5311 24024 5356 24052
rect 5350 24012 5356 24024
rect 5408 24012 5414 24064
rect 6457 24055 6515 24061
rect 6457 24021 6469 24055
rect 6503 24052 6515 24055
rect 6730 24052 6736 24064
rect 6503 24024 6736 24052
rect 6503 24021 6515 24024
rect 6457 24015 6515 24021
rect 6730 24012 6736 24024
rect 6788 24012 6794 24064
rect 6825 24055 6883 24061
rect 6825 24021 6837 24055
rect 6871 24052 6883 24055
rect 6914 24052 6920 24064
rect 6871 24024 6920 24052
rect 6871 24021 6883 24024
rect 6825 24015 6883 24021
rect 6914 24012 6920 24024
rect 6972 24012 6978 24064
rect 8662 24052 8668 24064
rect 8623 24024 8668 24052
rect 8662 24012 8668 24024
rect 8720 24012 8726 24064
rect 12342 24052 12348 24064
rect 12303 24024 12348 24052
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 12434 24012 12440 24064
rect 12492 24052 12498 24064
rect 12710 24052 12716 24064
rect 12492 24024 12716 24052
rect 12492 24012 12498 24024
rect 12710 24012 12716 24024
rect 12768 24012 12774 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 4430 23808 4436 23860
rect 4488 23848 4494 23860
rect 5169 23851 5227 23857
rect 5169 23848 5181 23851
rect 4488 23820 5181 23848
rect 4488 23808 4494 23820
rect 5169 23817 5181 23820
rect 5215 23848 5227 23851
rect 5902 23848 5908 23860
rect 5215 23820 5908 23848
rect 5215 23817 5227 23820
rect 5169 23811 5227 23817
rect 5902 23808 5908 23820
rect 5960 23808 5966 23860
rect 7006 23848 7012 23860
rect 6967 23820 7012 23848
rect 7006 23808 7012 23820
rect 7064 23808 7070 23860
rect 9858 23808 9864 23860
rect 9916 23848 9922 23860
rect 9953 23851 10011 23857
rect 9953 23848 9965 23851
rect 9916 23820 9965 23848
rect 9916 23808 9922 23820
rect 9953 23817 9965 23820
rect 9999 23817 10011 23851
rect 11514 23848 11520 23860
rect 11475 23820 11520 23848
rect 9953 23811 10011 23817
rect 5813 23783 5871 23789
rect 5813 23749 5825 23783
rect 5859 23780 5871 23783
rect 5994 23780 6000 23792
rect 5859 23752 6000 23780
rect 5859 23749 5871 23752
rect 5813 23743 5871 23749
rect 5994 23740 6000 23752
rect 6052 23740 6058 23792
rect 7926 23780 7932 23792
rect 7484 23752 7932 23780
rect 5166 23672 5172 23724
rect 5224 23712 5230 23724
rect 7484 23721 7512 23752
rect 7926 23740 7932 23752
rect 7984 23780 7990 23792
rect 8573 23783 8631 23789
rect 8573 23780 8585 23783
rect 7984 23752 8585 23780
rect 7984 23740 7990 23752
rect 8573 23749 8585 23752
rect 8619 23749 8631 23783
rect 8573 23743 8631 23749
rect 5261 23715 5319 23721
rect 5261 23712 5273 23715
rect 5224 23684 5273 23712
rect 5224 23672 5230 23684
rect 5261 23681 5273 23684
rect 5307 23681 5319 23715
rect 5261 23675 5319 23681
rect 7469 23715 7527 23721
rect 7469 23681 7481 23715
rect 7515 23681 7527 23715
rect 7469 23675 7527 23681
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23712 7619 23715
rect 8202 23712 8208 23724
rect 7607 23684 8208 23712
rect 7607 23681 7619 23684
rect 7561 23675 7619 23681
rect 3053 23647 3111 23653
rect 3053 23613 3065 23647
rect 3099 23644 3111 23647
rect 3142 23644 3148 23656
rect 3099 23616 3148 23644
rect 3099 23613 3111 23616
rect 3053 23607 3111 23613
rect 3142 23604 3148 23616
rect 3200 23644 3206 23656
rect 3878 23644 3884 23656
rect 3200 23616 3884 23644
rect 3200 23604 3206 23616
rect 3878 23604 3884 23616
rect 3936 23604 3942 23656
rect 5626 23604 5632 23656
rect 5684 23644 5690 23656
rect 5994 23644 6000 23656
rect 5684 23616 6000 23644
rect 5684 23604 5690 23616
rect 5994 23604 6000 23616
rect 6052 23604 6058 23656
rect 6273 23647 6331 23653
rect 6273 23613 6285 23647
rect 6319 23644 6331 23647
rect 6638 23644 6644 23656
rect 6319 23616 6644 23644
rect 6319 23613 6331 23616
rect 6273 23607 6331 23613
rect 6638 23604 6644 23616
rect 6696 23644 6702 23656
rect 7190 23644 7196 23656
rect 6696 23616 7196 23644
rect 6696 23604 6702 23616
rect 7190 23604 7196 23616
rect 7248 23644 7254 23656
rect 7576 23644 7604 23675
rect 8202 23672 8208 23684
rect 8260 23672 8266 23724
rect 8662 23672 8668 23724
rect 8720 23712 8726 23724
rect 9033 23715 9091 23721
rect 9033 23712 9045 23715
rect 8720 23684 9045 23712
rect 8720 23672 8726 23684
rect 9033 23681 9045 23684
rect 9079 23681 9091 23715
rect 9214 23712 9220 23724
rect 9175 23684 9220 23712
rect 9033 23675 9091 23681
rect 9214 23672 9220 23684
rect 9272 23672 9278 23724
rect 9968 23712 9996 23811
rect 11514 23808 11520 23820
rect 11572 23848 11578 23860
rect 12526 23848 12532 23860
rect 11572 23820 12532 23848
rect 11572 23808 11578 23820
rect 12526 23808 12532 23820
rect 12584 23808 12590 23860
rect 11885 23783 11943 23789
rect 11885 23749 11897 23783
rect 11931 23780 11943 23783
rect 12894 23780 12900 23792
rect 11931 23752 12900 23780
rect 11931 23749 11943 23752
rect 11885 23743 11943 23749
rect 12894 23740 12900 23752
rect 12952 23740 12958 23792
rect 9968 23684 10272 23712
rect 8386 23644 8392 23656
rect 7248 23616 7604 23644
rect 7659 23616 8392 23644
rect 7248 23604 7254 23616
rect 2961 23579 3019 23585
rect 2961 23545 2973 23579
rect 3007 23576 3019 23579
rect 3298 23579 3356 23585
rect 3298 23576 3310 23579
rect 3007 23548 3310 23576
rect 3007 23545 3019 23548
rect 2961 23539 3019 23545
rect 3298 23545 3310 23548
rect 3344 23576 3356 23579
rect 3510 23576 3516 23588
rect 3344 23548 3516 23576
rect 3344 23545 3356 23548
rect 3298 23539 3356 23545
rect 3510 23536 3516 23548
rect 3568 23536 3574 23588
rect 4801 23579 4859 23585
rect 4801 23545 4813 23579
rect 4847 23576 4859 23579
rect 6086 23576 6092 23588
rect 4847 23548 6092 23576
rect 4847 23545 4859 23548
rect 4801 23539 4859 23545
rect 6086 23536 6092 23548
rect 6144 23536 6150 23588
rect 6914 23536 6920 23588
rect 6972 23576 6978 23588
rect 7377 23579 7435 23585
rect 7377 23576 7389 23579
rect 6972 23548 7389 23576
rect 6972 23536 6978 23548
rect 7377 23545 7389 23548
rect 7423 23576 7435 23579
rect 7659 23576 7687 23616
rect 8386 23604 8392 23616
rect 8444 23604 8450 23656
rect 8481 23647 8539 23653
rect 8481 23613 8493 23647
rect 8527 23644 8539 23647
rect 9232 23644 9260 23672
rect 8527 23616 9260 23644
rect 10137 23647 10195 23653
rect 8527 23613 8539 23616
rect 8481 23607 8539 23613
rect 10137 23613 10149 23647
rect 10183 23613 10195 23647
rect 10244 23644 10272 23684
rect 12434 23672 12440 23724
rect 12492 23672 12498 23724
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23712 13139 23715
rect 13262 23712 13268 23724
rect 13127 23684 13268 23712
rect 13127 23681 13139 23684
rect 13081 23675 13139 23681
rect 13262 23672 13268 23684
rect 13320 23672 13326 23724
rect 10393 23647 10451 23653
rect 10393 23644 10405 23647
rect 10244 23616 10405 23644
rect 10137 23607 10195 23613
rect 10393 23613 10405 23616
rect 10439 23644 10451 23647
rect 12161 23647 12219 23653
rect 12161 23644 12173 23647
rect 10439 23616 12173 23644
rect 10439 23613 10451 23616
rect 10393 23607 10451 23613
rect 12161 23613 12173 23616
rect 12207 23613 12219 23647
rect 12161 23607 12219 23613
rect 7423 23548 7687 23576
rect 7423 23545 7435 23548
rect 7377 23539 7435 23545
rect 8018 23536 8024 23588
rect 8076 23576 8082 23588
rect 8113 23579 8171 23585
rect 8113 23576 8125 23579
rect 8076 23548 8125 23576
rect 8076 23536 8082 23548
rect 8113 23545 8125 23548
rect 8159 23576 8171 23579
rect 8941 23579 8999 23585
rect 8941 23576 8953 23579
rect 8159 23548 8953 23576
rect 8159 23545 8171 23548
rect 8113 23539 8171 23545
rect 8941 23545 8953 23548
rect 8987 23545 8999 23579
rect 9674 23576 9680 23588
rect 9587 23548 9680 23576
rect 8941 23539 8999 23545
rect 9674 23536 9680 23548
rect 9732 23576 9738 23588
rect 10152 23576 10180 23607
rect 10686 23576 10692 23588
rect 9732 23548 10692 23576
rect 9732 23536 9738 23548
rect 10686 23536 10692 23548
rect 10744 23536 10750 23588
rect 12176 23576 12204 23607
rect 12342 23576 12348 23588
rect 12176 23548 12348 23576
rect 12342 23536 12348 23548
rect 12400 23576 12406 23588
rect 12452 23576 12480 23672
rect 12618 23604 12624 23656
rect 12676 23644 12682 23656
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12676 23616 12909 23644
rect 12676 23604 12682 23616
rect 12897 23613 12909 23616
rect 12943 23644 12955 23647
rect 13449 23647 13507 23653
rect 13449 23644 13461 23647
rect 12943 23616 13461 23644
rect 12943 23613 12955 23616
rect 12897 23607 12955 23613
rect 13449 23613 13461 23616
rect 13495 23613 13507 23647
rect 13449 23607 13507 23613
rect 12400 23548 12480 23576
rect 12400 23536 12406 23548
rect 12710 23536 12716 23588
rect 12768 23576 12774 23588
rect 12805 23579 12863 23585
rect 12805 23576 12817 23579
rect 12768 23548 12817 23576
rect 12768 23536 12774 23548
rect 12805 23545 12817 23548
rect 12851 23576 12863 23579
rect 13817 23579 13875 23585
rect 13817 23576 13829 23579
rect 12851 23548 13829 23576
rect 12851 23545 12863 23548
rect 12805 23539 12863 23545
rect 13817 23545 13829 23548
rect 13863 23545 13875 23579
rect 13817 23539 13875 23545
rect 4154 23468 4160 23520
rect 4212 23508 4218 23520
rect 4433 23511 4491 23517
rect 4433 23508 4445 23511
rect 4212 23480 4445 23508
rect 4212 23468 4218 23480
rect 4433 23477 4445 23480
rect 4479 23477 4491 23511
rect 4433 23471 4491 23477
rect 4614 23468 4620 23520
rect 4672 23508 4678 23520
rect 5166 23508 5172 23520
rect 4672 23480 5172 23508
rect 4672 23468 4678 23480
rect 5166 23468 5172 23480
rect 5224 23468 5230 23520
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 12492 23480 12537 23508
rect 12492 23468 12498 23480
rect 12618 23468 12624 23520
rect 12676 23508 12682 23520
rect 13170 23508 13176 23520
rect 12676 23480 13176 23508
rect 12676 23468 12682 23480
rect 13170 23468 13176 23480
rect 13228 23468 13234 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 3050 23264 3056 23316
rect 3108 23304 3114 23316
rect 4798 23304 4804 23316
rect 3108 23276 4804 23304
rect 3108 23264 3114 23276
rect 4798 23264 4804 23276
rect 4856 23264 4862 23316
rect 6457 23307 6515 23313
rect 6457 23273 6469 23307
rect 6503 23304 6515 23307
rect 6822 23304 6828 23316
rect 6503 23276 6828 23304
rect 6503 23273 6515 23276
rect 6457 23267 6515 23273
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 7558 23304 7564 23316
rect 7519 23276 7564 23304
rect 7558 23264 7564 23276
rect 7616 23264 7622 23316
rect 8018 23304 8024 23316
rect 7979 23276 8024 23304
rect 8018 23264 8024 23276
rect 8076 23264 8082 23316
rect 11054 23304 11060 23316
rect 11015 23276 11060 23304
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 12250 23264 12256 23316
rect 12308 23304 12314 23316
rect 12894 23304 12900 23316
rect 12308 23276 12900 23304
rect 12308 23264 12314 23276
rect 12894 23264 12900 23276
rect 12952 23264 12958 23316
rect 2317 23239 2375 23245
rect 2317 23205 2329 23239
rect 2363 23236 2375 23239
rect 2774 23236 2780 23248
rect 2363 23208 2780 23236
rect 2363 23205 2375 23208
rect 2317 23199 2375 23205
rect 2774 23196 2780 23208
rect 2832 23196 2838 23248
rect 4430 23245 4436 23248
rect 4424 23236 4436 23245
rect 4391 23208 4436 23236
rect 4424 23199 4436 23208
rect 4430 23196 4436 23199
rect 4488 23196 4494 23248
rect 7926 23236 7932 23248
rect 7887 23208 7932 23236
rect 7926 23196 7932 23208
rect 7984 23196 7990 23248
rect 10686 23196 10692 23248
rect 10744 23236 10750 23248
rect 11333 23239 11391 23245
rect 11333 23236 11345 23239
rect 10744 23208 11345 23236
rect 10744 23196 10750 23208
rect 11333 23205 11345 23208
rect 11379 23236 11391 23239
rect 11422 23236 11428 23248
rect 11379 23208 11428 23236
rect 11379 23205 11391 23208
rect 11333 23199 11391 23205
rect 11422 23196 11428 23208
rect 11480 23196 11486 23248
rect 12526 23196 12532 23248
rect 12584 23245 12590 23248
rect 12584 23239 12648 23245
rect 12584 23205 12602 23239
rect 12636 23205 12648 23239
rect 12584 23199 12648 23205
rect 12584 23196 12590 23199
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 3878 23168 3884 23180
rect 2924 23140 2969 23168
rect 3791 23140 3884 23168
rect 2924 23128 2930 23140
rect 3878 23128 3884 23140
rect 3936 23168 3942 23180
rect 6822 23168 6828 23180
rect 3936 23140 4200 23168
rect 6783 23140 6828 23168
rect 3936 23128 3942 23140
rect 4172 23112 4200 23140
rect 6822 23128 6828 23140
rect 6880 23128 6886 23180
rect 8202 23128 8208 23180
rect 8260 23168 8266 23180
rect 8389 23171 8447 23177
rect 8389 23168 8401 23171
rect 8260 23140 8401 23168
rect 8260 23128 8266 23140
rect 8389 23137 8401 23140
rect 8435 23137 8447 23171
rect 9933 23171 9991 23177
rect 9933 23168 9945 23171
rect 8389 23131 8447 23137
rect 8772 23140 9945 23168
rect 8772 23112 8800 23140
rect 9933 23137 9945 23140
rect 9979 23168 9991 23171
rect 10226 23168 10232 23180
rect 9979 23140 10232 23168
rect 9979 23137 9991 23140
rect 9933 23131 9991 23137
rect 10226 23128 10232 23140
rect 10284 23128 10290 23180
rect 11440 23168 11468 23196
rect 12345 23171 12403 23177
rect 12345 23168 12357 23171
rect 11440 23140 12357 23168
rect 12345 23137 12357 23140
rect 12391 23168 12403 23171
rect 12434 23168 12440 23180
rect 12391 23140 12440 23168
rect 12391 23137 12403 23140
rect 12345 23131 12403 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 2958 23100 2964 23112
rect 2919 23072 2964 23100
rect 2958 23060 2964 23072
rect 3016 23100 3022 23112
rect 4062 23100 4068 23112
rect 3016 23072 4068 23100
rect 3016 23060 3022 23072
rect 4062 23060 4068 23072
rect 4120 23060 4126 23112
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 4212 23072 4257 23100
rect 4212 23060 4218 23072
rect 6178 23060 6184 23112
rect 6236 23100 6242 23112
rect 6914 23100 6920 23112
rect 6236 23072 6920 23100
rect 6236 23060 6242 23072
rect 6914 23060 6920 23072
rect 6972 23060 6978 23112
rect 7009 23103 7067 23109
rect 7009 23069 7021 23103
rect 7055 23069 7067 23103
rect 7009 23063 7067 23069
rect 6638 22992 6644 23044
rect 6696 23032 6702 23044
rect 7024 23032 7052 23063
rect 7190 23060 7196 23112
rect 7248 23100 7254 23112
rect 8481 23103 8539 23109
rect 8481 23100 8493 23103
rect 7248 23072 8493 23100
rect 7248 23060 7254 23072
rect 8481 23069 8493 23072
rect 8527 23069 8539 23103
rect 8481 23063 8539 23069
rect 8665 23103 8723 23109
rect 8665 23069 8677 23103
rect 8711 23100 8723 23103
rect 8754 23100 8760 23112
rect 8711 23072 8760 23100
rect 8711 23069 8723 23072
rect 8665 23063 8723 23069
rect 8754 23060 8760 23072
rect 8812 23060 8818 23112
rect 9674 23100 9680 23112
rect 9635 23072 9680 23100
rect 9674 23060 9680 23072
rect 9732 23060 9738 23112
rect 6696 23004 7052 23032
rect 6696 22992 6702 23004
rect 2406 22964 2412 22976
rect 2367 22936 2412 22964
rect 2406 22924 2412 22936
rect 2464 22924 2470 22976
rect 4890 22924 4896 22976
rect 4948 22964 4954 22976
rect 5537 22967 5595 22973
rect 5537 22964 5549 22967
rect 4948 22936 5549 22964
rect 4948 22924 4954 22936
rect 5537 22933 5549 22936
rect 5583 22933 5595 22967
rect 5537 22927 5595 22933
rect 9674 22924 9680 22976
rect 9732 22964 9738 22976
rect 9858 22964 9864 22976
rect 9732 22936 9864 22964
rect 9732 22924 9738 22936
rect 9858 22924 9864 22936
rect 9916 22924 9922 22976
rect 13446 22924 13452 22976
rect 13504 22964 13510 22976
rect 13725 22967 13783 22973
rect 13725 22964 13737 22967
rect 13504 22936 13737 22964
rect 13504 22924 13510 22936
rect 13725 22933 13737 22936
rect 13771 22933 13783 22967
rect 13725 22927 13783 22933
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 2866 22720 2872 22772
rect 2924 22760 2930 22772
rect 4341 22763 4399 22769
rect 4341 22760 4353 22763
rect 2924 22732 4353 22760
rect 2924 22720 2930 22732
rect 4341 22729 4353 22732
rect 4387 22729 4399 22763
rect 5350 22760 5356 22772
rect 4341 22723 4399 22729
rect 4816 22732 5356 22760
rect 2777 22695 2835 22701
rect 2777 22661 2789 22695
rect 2823 22692 2835 22695
rect 4430 22692 4436 22704
rect 2823 22664 4436 22692
rect 2823 22661 2835 22664
rect 2777 22655 2835 22661
rect 4430 22652 4436 22664
rect 4488 22652 4494 22704
rect 1578 22624 1584 22636
rect 1539 22596 1584 22624
rect 1578 22584 1584 22596
rect 1636 22584 1642 22636
rect 2317 22627 2375 22633
rect 2317 22593 2329 22627
rect 2363 22624 2375 22627
rect 2958 22624 2964 22636
rect 2363 22596 2964 22624
rect 2363 22593 2375 22596
rect 2317 22587 2375 22593
rect 2958 22584 2964 22596
rect 3016 22584 3022 22636
rect 3421 22627 3479 22633
rect 3421 22593 3433 22627
rect 3467 22593 3479 22627
rect 3421 22587 3479 22593
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 1670 22556 1676 22568
rect 1443 22528 1676 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 1670 22516 1676 22528
rect 1728 22556 1734 22568
rect 2406 22556 2412 22568
rect 1728 22528 2412 22556
rect 1728 22516 1734 22528
rect 2406 22516 2412 22528
rect 2464 22516 2470 22568
rect 2685 22559 2743 22565
rect 2685 22525 2697 22559
rect 2731 22556 2743 22559
rect 3050 22556 3056 22568
rect 2731 22528 3056 22556
rect 2731 22525 2743 22528
rect 2685 22519 2743 22525
rect 3050 22516 3056 22528
rect 3108 22556 3114 22568
rect 3145 22559 3203 22565
rect 3145 22556 3157 22559
rect 3108 22528 3157 22556
rect 3108 22516 3114 22528
rect 3145 22525 3157 22528
rect 3191 22525 3203 22559
rect 3145 22519 3203 22525
rect 3234 22516 3240 22568
rect 3292 22556 3298 22568
rect 3436 22556 3464 22587
rect 3510 22584 3516 22636
rect 3568 22624 3574 22636
rect 3789 22627 3847 22633
rect 3789 22624 3801 22627
rect 3568 22596 3801 22624
rect 3568 22584 3574 22596
rect 3789 22593 3801 22596
rect 3835 22593 3847 22627
rect 3789 22587 3847 22593
rect 4249 22627 4307 22633
rect 4249 22593 4261 22627
rect 4295 22624 4307 22627
rect 4338 22624 4344 22636
rect 4295 22596 4344 22624
rect 4295 22593 4307 22596
rect 4249 22587 4307 22593
rect 4338 22584 4344 22596
rect 4396 22584 4402 22636
rect 4816 22633 4844 22732
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 6178 22760 6184 22772
rect 6139 22732 6184 22760
rect 6178 22720 6184 22732
rect 6236 22720 6242 22772
rect 6549 22763 6607 22769
rect 6549 22729 6561 22763
rect 6595 22760 6607 22763
rect 6638 22760 6644 22772
rect 6595 22732 6644 22760
rect 6595 22729 6607 22732
rect 6549 22723 6607 22729
rect 6638 22720 6644 22732
rect 6696 22720 6702 22772
rect 8294 22720 8300 22772
rect 8352 22720 8358 22772
rect 8662 22720 8668 22772
rect 8720 22760 8726 22772
rect 9585 22763 9643 22769
rect 9585 22760 9597 22763
rect 8720 22732 9597 22760
rect 8720 22720 8726 22732
rect 9585 22729 9597 22732
rect 9631 22729 9643 22763
rect 9585 22723 9643 22729
rect 10962 22720 10968 22772
rect 11020 22760 11026 22772
rect 11422 22760 11428 22772
rect 11020 22732 11428 22760
rect 11020 22720 11026 22732
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 12989 22763 13047 22769
rect 12989 22760 13001 22763
rect 12492 22732 13001 22760
rect 12492 22720 12498 22732
rect 12989 22729 13001 22732
rect 13035 22729 13047 22763
rect 12989 22723 13047 22729
rect 7190 22692 7196 22704
rect 7151 22664 7196 22692
rect 7190 22652 7196 22664
rect 7248 22652 7254 22704
rect 8312 22692 8340 22720
rect 8757 22695 8815 22701
rect 8757 22692 8769 22695
rect 8312 22664 8769 22692
rect 8757 22661 8769 22664
rect 8803 22661 8815 22695
rect 8757 22655 8815 22661
rect 12526 22652 12532 22704
rect 12584 22692 12590 22704
rect 12621 22695 12679 22701
rect 12621 22692 12633 22695
rect 12584 22664 12633 22692
rect 12584 22652 12590 22664
rect 12621 22661 12633 22664
rect 12667 22661 12679 22695
rect 12621 22655 12679 22661
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22593 4859 22627
rect 4801 22587 4859 22593
rect 4890 22584 4896 22636
rect 4948 22624 4954 22636
rect 4985 22627 5043 22633
rect 4985 22624 4997 22627
rect 4948 22596 4997 22624
rect 4948 22584 4954 22596
rect 4985 22593 4997 22596
rect 5031 22593 5043 22627
rect 10226 22624 10232 22636
rect 10187 22596 10232 22624
rect 4985 22587 5043 22593
rect 10226 22584 10232 22596
rect 10284 22624 10290 22636
rect 10597 22627 10655 22633
rect 10597 22624 10609 22627
rect 10284 22596 10609 22624
rect 10284 22584 10290 22596
rect 10597 22593 10609 22596
rect 10643 22624 10655 22627
rect 10965 22627 11023 22633
rect 10965 22624 10977 22627
rect 10643 22596 10977 22624
rect 10643 22593 10655 22596
rect 10597 22587 10655 22593
rect 10965 22593 10977 22596
rect 11011 22593 11023 22627
rect 10965 22587 11023 22593
rect 5813 22559 5871 22565
rect 3292 22528 3556 22556
rect 3292 22516 3298 22528
rect 3528 22488 3556 22528
rect 5813 22525 5825 22559
rect 5859 22556 5871 22559
rect 6822 22556 6828 22568
rect 5859 22528 6828 22556
rect 5859 22525 5871 22528
rect 5813 22519 5871 22525
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 7374 22556 7380 22568
rect 7335 22528 7380 22556
rect 7374 22516 7380 22528
rect 7432 22516 7438 22568
rect 8018 22516 8024 22568
rect 8076 22556 8082 22568
rect 9401 22559 9459 22565
rect 9401 22556 9413 22559
rect 8076 22528 9413 22556
rect 8076 22516 8082 22528
rect 9401 22525 9413 22528
rect 9447 22556 9459 22559
rect 10045 22559 10103 22565
rect 10045 22556 10057 22559
rect 9447 22528 10057 22556
rect 9447 22525 9459 22528
rect 9401 22519 9459 22525
rect 10045 22525 10057 22528
rect 10091 22525 10103 22559
rect 10045 22519 10103 22525
rect 4338 22488 4344 22500
rect 3528 22460 4344 22488
rect 4338 22448 4344 22460
rect 4396 22448 4402 22500
rect 4982 22488 4988 22500
rect 4439 22460 4988 22488
rect 2958 22380 2964 22432
rect 3016 22420 3022 22432
rect 3237 22423 3295 22429
rect 3237 22420 3249 22423
rect 3016 22392 3249 22420
rect 3016 22380 3022 22392
rect 3237 22389 3249 22392
rect 3283 22420 3295 22423
rect 3418 22420 3424 22432
rect 3283 22392 3424 22420
rect 3283 22389 3295 22392
rect 3237 22383 3295 22389
rect 3418 22380 3424 22392
rect 3476 22420 3482 22432
rect 4439 22420 4467 22460
rect 4982 22448 4988 22460
rect 5040 22448 5046 22500
rect 7558 22448 7564 22500
rect 7616 22497 7622 22500
rect 7616 22491 7680 22497
rect 7616 22457 7634 22491
rect 7668 22457 7680 22491
rect 7616 22451 7680 22457
rect 7616 22448 7622 22451
rect 8294 22448 8300 22500
rect 8352 22488 8358 22500
rect 8478 22488 8484 22500
rect 8352 22460 8484 22488
rect 8352 22448 8358 22460
rect 8478 22448 8484 22460
rect 8536 22488 8542 22500
rect 9033 22491 9091 22497
rect 9033 22488 9045 22491
rect 8536 22460 9045 22488
rect 8536 22448 8542 22460
rect 9033 22457 9045 22460
rect 9079 22488 9091 22491
rect 9953 22491 10011 22497
rect 9953 22488 9965 22491
rect 9079 22460 9965 22488
rect 9079 22457 9091 22460
rect 9033 22451 9091 22457
rect 9953 22457 9965 22460
rect 9999 22457 10011 22491
rect 9953 22451 10011 22457
rect 3476 22392 4467 22420
rect 3476 22380 3482 22392
rect 4614 22380 4620 22432
rect 4672 22420 4678 22432
rect 4709 22423 4767 22429
rect 4709 22420 4721 22423
rect 4672 22392 4721 22420
rect 4672 22380 4678 22392
rect 4709 22389 4721 22392
rect 4755 22389 4767 22423
rect 4709 22383 4767 22389
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 1670 22216 1676 22228
rect 1631 22188 1676 22216
rect 1670 22176 1676 22188
rect 1728 22176 1734 22228
rect 2777 22219 2835 22225
rect 2777 22185 2789 22219
rect 2823 22216 2835 22219
rect 2958 22216 2964 22228
rect 2823 22188 2964 22216
rect 2823 22185 2835 22188
rect 2777 22179 2835 22185
rect 2958 22176 2964 22188
rect 3016 22176 3022 22228
rect 3234 22216 3240 22228
rect 3195 22188 3240 22216
rect 3234 22176 3240 22188
rect 3292 22176 3298 22228
rect 4062 22176 4068 22228
rect 4120 22216 4126 22228
rect 4709 22219 4767 22225
rect 4709 22216 4721 22219
rect 4120 22188 4721 22216
rect 4120 22176 4126 22188
rect 4709 22185 4721 22188
rect 4755 22216 4767 22219
rect 5074 22216 5080 22228
rect 4755 22188 5080 22216
rect 4755 22185 4767 22188
rect 4709 22179 4767 22185
rect 5074 22176 5080 22188
rect 5132 22176 5138 22228
rect 8754 22216 8760 22228
rect 8312 22188 8760 22216
rect 2866 22148 2872 22160
rect 2792 22120 2872 22148
rect 2501 22083 2559 22089
rect 2501 22049 2513 22083
rect 2547 22080 2559 22083
rect 2792 22080 2820 22120
rect 2866 22108 2872 22120
rect 2924 22108 2930 22160
rect 3510 22108 3516 22160
rect 3568 22148 3574 22160
rect 4890 22148 4896 22160
rect 3568 22120 4896 22148
rect 3568 22108 3574 22120
rect 4890 22108 4896 22120
rect 4948 22148 4954 22160
rect 6730 22148 6736 22160
rect 4948 22120 5028 22148
rect 4948 22108 4954 22120
rect 2547 22052 2820 22080
rect 2547 22049 2559 22052
rect 2501 22043 2559 22049
rect 4430 21972 4436 22024
rect 4488 22012 4494 22024
rect 5000 22021 5028 22120
rect 5736 22120 6736 22148
rect 5736 22024 5764 22120
rect 6730 22108 6736 22120
rect 6788 22148 6794 22160
rect 7374 22148 7380 22160
rect 6788 22120 7380 22148
rect 6788 22108 6794 22120
rect 7374 22108 7380 22120
rect 7432 22148 7438 22160
rect 7561 22151 7619 22157
rect 7561 22148 7573 22151
rect 7432 22120 7573 22148
rect 7432 22108 7438 22120
rect 7561 22117 7573 22120
rect 7607 22117 7619 22151
rect 7561 22111 7619 22117
rect 5810 22040 5816 22092
rect 5868 22080 5874 22092
rect 6161 22083 6219 22089
rect 6161 22080 6173 22083
rect 5868 22052 6173 22080
rect 5868 22040 5874 22052
rect 6161 22049 6173 22052
rect 6207 22049 6219 22083
rect 6161 22043 6219 22049
rect 8021 22083 8079 22089
rect 8021 22049 8033 22083
rect 8067 22080 8079 22083
rect 8312 22080 8340 22188
rect 8754 22176 8760 22188
rect 8812 22176 8818 22228
rect 11146 22176 11152 22228
rect 11204 22176 11210 22228
rect 11164 22092 11192 22176
rect 10042 22080 10048 22092
rect 8067 22052 8340 22080
rect 10003 22052 10048 22080
rect 8067 22049 8079 22052
rect 8021 22043 8079 22049
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 11146 22040 11152 22092
rect 11204 22040 11210 22092
rect 13446 22080 13452 22092
rect 13407 22052 13452 22080
rect 13446 22040 13452 22052
rect 13504 22040 13510 22092
rect 4801 22015 4859 22021
rect 4801 22012 4813 22015
rect 4488 21984 4813 22012
rect 4488 21972 4494 21984
rect 4801 21981 4813 21984
rect 4847 21981 4859 22015
rect 4801 21975 4859 21981
rect 4985 22015 5043 22021
rect 4985 21981 4997 22015
rect 5031 21981 5043 22015
rect 4985 21975 5043 21981
rect 5718 21972 5724 22024
rect 5776 22012 5782 22024
rect 5905 22015 5963 22021
rect 5905 22012 5917 22015
rect 5776 21984 5917 22012
rect 5776 21972 5782 21984
rect 5905 21981 5917 21984
rect 5951 21981 5963 22015
rect 8110 22012 8116 22024
rect 8071 21984 8116 22012
rect 5905 21975 5963 21981
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 9858 21972 9864 22024
rect 9916 22012 9922 22024
rect 10137 22015 10195 22021
rect 10137 22012 10149 22015
rect 9916 21984 10149 22012
rect 9916 21972 9922 21984
rect 10137 21981 10149 21984
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 10226 21972 10232 22024
rect 10284 22012 10290 22024
rect 10284 21984 10329 22012
rect 10284 21972 10290 21984
rect 2774 21904 2780 21956
rect 2832 21944 2838 21956
rect 4341 21947 4399 21953
rect 4341 21944 4353 21947
rect 2832 21916 4353 21944
rect 2832 21904 2838 21916
rect 4341 21913 4353 21916
rect 4387 21913 4399 21947
rect 13630 21944 13636 21956
rect 13591 21916 13636 21944
rect 4341 21907 4399 21913
rect 13630 21904 13636 21916
rect 13688 21904 13694 21956
rect 3881 21879 3939 21885
rect 3881 21845 3893 21879
rect 3927 21876 3939 21879
rect 4614 21876 4620 21888
rect 3927 21848 4620 21876
rect 3927 21845 3939 21848
rect 3881 21839 3939 21845
rect 4614 21836 4620 21848
rect 4672 21876 4678 21888
rect 4798 21876 4804 21888
rect 4672 21848 4804 21876
rect 4672 21836 4678 21848
rect 4798 21836 4804 21848
rect 4856 21836 4862 21888
rect 7098 21836 7104 21888
rect 7156 21876 7162 21888
rect 7285 21879 7343 21885
rect 7285 21876 7297 21879
rect 7156 21848 7297 21876
rect 7156 21836 7162 21848
rect 7285 21845 7297 21848
rect 7331 21845 7343 21879
rect 7285 21839 7343 21845
rect 8202 21836 8208 21888
rect 8260 21876 8266 21888
rect 8478 21876 8484 21888
rect 8260 21848 8484 21876
rect 8260 21836 8266 21848
rect 8478 21836 8484 21848
rect 8536 21876 8542 21888
rect 8573 21879 8631 21885
rect 8573 21876 8585 21879
rect 8536 21848 8585 21876
rect 8536 21836 8542 21848
rect 8573 21845 8585 21848
rect 8619 21845 8631 21879
rect 8573 21839 8631 21845
rect 9306 21836 9312 21888
rect 9364 21876 9370 21888
rect 9677 21879 9735 21885
rect 9677 21876 9689 21879
rect 9364 21848 9689 21876
rect 9364 21836 9370 21848
rect 9677 21845 9689 21848
rect 9723 21845 9735 21879
rect 9677 21839 9735 21845
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 3510 21632 3516 21684
rect 3568 21672 3574 21684
rect 3881 21675 3939 21681
rect 3881 21672 3893 21675
rect 3568 21644 3893 21672
rect 3568 21632 3574 21644
rect 3881 21641 3893 21644
rect 3927 21641 3939 21675
rect 4798 21672 4804 21684
rect 4759 21644 4804 21672
rect 3881 21635 3939 21641
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 6914 21632 6920 21684
rect 6972 21672 6978 21684
rect 7285 21675 7343 21681
rect 7285 21672 7297 21675
rect 6972 21644 7297 21672
rect 6972 21632 6978 21644
rect 7285 21641 7297 21644
rect 7331 21641 7343 21675
rect 7285 21635 7343 21641
rect 8386 21632 8392 21684
rect 8444 21672 8450 21684
rect 8849 21675 8907 21681
rect 8849 21672 8861 21675
rect 8444 21644 8861 21672
rect 8444 21632 8450 21644
rect 8849 21641 8861 21644
rect 8895 21641 8907 21675
rect 8849 21635 8907 21641
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 10229 21675 10287 21681
rect 10229 21672 10241 21675
rect 10100 21644 10241 21672
rect 10100 21632 10106 21644
rect 10229 21641 10241 21644
rect 10275 21641 10287 21675
rect 10229 21635 10287 21641
rect 3605 21607 3663 21613
rect 3605 21573 3617 21607
rect 3651 21604 3663 21607
rect 4062 21604 4068 21616
rect 3651 21576 4068 21604
rect 3651 21573 3663 21576
rect 3605 21567 3663 21573
rect 4062 21564 4068 21576
rect 4120 21564 4126 21616
rect 4338 21536 4344 21548
rect 4251 21508 4344 21536
rect 4338 21496 4344 21508
rect 4396 21536 4402 21548
rect 5442 21536 5448 21548
rect 4396 21508 5448 21536
rect 4396 21496 4402 21508
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21536 6699 21539
rect 7558 21536 7564 21548
rect 6687 21508 7564 21536
rect 6687 21505 6699 21508
rect 6641 21499 6699 21505
rect 7558 21496 7564 21508
rect 7616 21536 7622 21548
rect 7837 21539 7895 21545
rect 7837 21536 7849 21539
rect 7616 21508 7849 21536
rect 7616 21496 7622 21508
rect 7837 21505 7849 21508
rect 7883 21505 7895 21539
rect 7837 21499 7895 21505
rect 8389 21539 8447 21545
rect 8389 21505 8401 21539
rect 8435 21536 8447 21539
rect 9306 21536 9312 21548
rect 8435 21508 9312 21536
rect 8435 21505 8447 21508
rect 8389 21499 8447 21505
rect 9306 21496 9312 21508
rect 9364 21496 9370 21548
rect 9490 21536 9496 21548
rect 9451 21508 9496 21536
rect 9490 21496 9496 21508
rect 9548 21496 9554 21548
rect 5534 21428 5540 21480
rect 5592 21468 5598 21480
rect 5902 21468 5908 21480
rect 5592 21440 5908 21468
rect 5592 21428 5598 21440
rect 5902 21428 5908 21440
rect 5960 21428 5966 21480
rect 7374 21428 7380 21480
rect 7432 21468 7438 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7432 21440 7665 21468
rect 7432 21428 7438 21440
rect 7653 21437 7665 21440
rect 7699 21468 7711 21471
rect 8110 21468 8116 21480
rect 7699 21440 8116 21468
rect 7699 21437 7711 21440
rect 7653 21431 7711 21437
rect 8110 21428 8116 21440
rect 8168 21428 8174 21480
rect 4709 21403 4767 21409
rect 4709 21369 4721 21403
rect 4755 21400 4767 21403
rect 5166 21400 5172 21412
rect 4755 21372 5172 21400
rect 4755 21369 4767 21372
rect 4709 21363 4767 21369
rect 5166 21360 5172 21372
rect 5224 21360 5230 21412
rect 4614 21292 4620 21344
rect 4672 21332 4678 21344
rect 5261 21335 5319 21341
rect 5261 21332 5273 21335
rect 4672 21304 5273 21332
rect 4672 21292 4678 21304
rect 5261 21301 5273 21304
rect 5307 21301 5319 21335
rect 5902 21332 5908 21344
rect 5863 21304 5908 21332
rect 5261 21295 5319 21301
rect 5902 21292 5908 21304
rect 5960 21292 5966 21344
rect 7193 21335 7251 21341
rect 7193 21301 7205 21335
rect 7239 21332 7251 21335
rect 7742 21332 7748 21344
rect 7239 21304 7748 21332
rect 7239 21301 7251 21304
rect 7193 21295 7251 21301
rect 7742 21292 7748 21304
rect 7800 21292 7806 21344
rect 8570 21292 8576 21344
rect 8628 21332 8634 21344
rect 8665 21335 8723 21341
rect 8665 21332 8677 21335
rect 8628 21304 8677 21332
rect 8628 21292 8634 21304
rect 8665 21301 8677 21304
rect 8711 21332 8723 21335
rect 9217 21335 9275 21341
rect 9217 21332 9229 21335
rect 8711 21304 9229 21332
rect 8711 21301 8723 21304
rect 8665 21295 8723 21301
rect 9217 21301 9229 21304
rect 9263 21301 9275 21335
rect 9858 21332 9864 21344
rect 9819 21304 9864 21332
rect 9217 21295 9275 21301
rect 9858 21292 9864 21304
rect 9916 21292 9922 21344
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 13446 21332 13452 21344
rect 12492 21304 13452 21332
rect 12492 21292 12498 21304
rect 13446 21292 13452 21304
rect 13504 21292 13510 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 4430 21128 4436 21140
rect 4391 21100 4436 21128
rect 4430 21088 4436 21100
rect 4488 21088 4494 21140
rect 6086 21128 6092 21140
rect 6047 21100 6092 21128
rect 6086 21088 6092 21100
rect 6144 21088 6150 21140
rect 7374 21128 7380 21140
rect 7335 21100 7380 21128
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 7834 21128 7840 21140
rect 7484 21100 7840 21128
rect 7484 21060 7512 21100
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 8202 21128 8208 21140
rect 8163 21100 8208 21128
rect 8202 21088 8208 21100
rect 8260 21088 8266 21140
rect 8478 21088 8484 21140
rect 8536 21128 8542 21140
rect 8938 21128 8944 21140
rect 8536 21100 8944 21128
rect 8536 21088 8542 21100
rect 8938 21088 8944 21100
rect 8996 21088 9002 21140
rect 9953 21131 10011 21137
rect 9953 21097 9965 21131
rect 9999 21128 10011 21131
rect 10226 21128 10232 21140
rect 9999 21100 10232 21128
rect 9999 21097 10011 21100
rect 9953 21091 10011 21097
rect 10226 21088 10232 21100
rect 10284 21088 10290 21140
rect 6472 21032 7512 21060
rect 6472 21004 6500 21032
rect 7558 21020 7564 21072
rect 7616 21060 7622 21072
rect 8849 21063 8907 21069
rect 8849 21060 8861 21063
rect 7616 21032 8861 21060
rect 7616 21020 7622 21032
rect 6454 20992 6460 21004
rect 6415 20964 6460 20992
rect 6454 20952 6460 20964
rect 6512 20952 6518 21004
rect 8404 20936 8432 21032
rect 8849 21029 8861 21032
rect 8895 21060 8907 21063
rect 9490 21060 9496 21072
rect 8895 21032 9496 21060
rect 8895 21029 8907 21032
rect 8849 21023 8907 21029
rect 9490 21020 9496 21032
rect 9548 21020 9554 21072
rect 10502 21001 10508 21004
rect 10496 20955 10508 21001
rect 10560 20992 10566 21004
rect 10560 20964 10596 20992
rect 10502 20952 10508 20955
rect 10560 20952 10566 20964
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 6086 20924 6092 20936
rect 5592 20896 6092 20924
rect 5592 20884 5598 20896
rect 6086 20884 6092 20896
rect 6144 20924 6150 20936
rect 6549 20927 6607 20933
rect 6549 20924 6561 20927
rect 6144 20896 6561 20924
rect 6144 20884 6150 20896
rect 6549 20893 6561 20896
rect 6595 20893 6607 20927
rect 6730 20924 6736 20936
rect 6691 20896 6736 20924
rect 6549 20887 6607 20893
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 8110 20884 8116 20936
rect 8168 20924 8174 20936
rect 8297 20927 8355 20933
rect 8297 20924 8309 20927
rect 8168 20896 8309 20924
rect 8168 20884 8174 20896
rect 8297 20893 8309 20896
rect 8343 20893 8355 20927
rect 8297 20887 8355 20893
rect 8386 20884 8392 20936
rect 8444 20924 8450 20936
rect 8444 20896 8537 20924
rect 8444 20884 8450 20896
rect 10134 20884 10140 20936
rect 10192 20924 10198 20936
rect 10229 20927 10287 20933
rect 10229 20924 10241 20927
rect 10192 20896 10241 20924
rect 10192 20884 10198 20896
rect 10229 20893 10241 20896
rect 10275 20893 10287 20927
rect 10229 20887 10287 20893
rect 2774 20816 2780 20868
rect 2832 20856 2838 20868
rect 4154 20856 4160 20868
rect 2832 20828 4160 20856
rect 2832 20816 2838 20828
rect 4154 20816 4160 20828
rect 4212 20856 4218 20868
rect 5718 20856 5724 20868
rect 4212 20828 5724 20856
rect 4212 20816 4218 20828
rect 5718 20816 5724 20828
rect 5776 20856 5782 20868
rect 5905 20859 5963 20865
rect 5905 20856 5917 20859
rect 5776 20828 5917 20856
rect 5776 20816 5782 20828
rect 5905 20825 5917 20828
rect 5951 20856 5963 20859
rect 6822 20856 6828 20868
rect 5951 20828 6828 20856
rect 5951 20825 5963 20828
rect 5905 20819 5963 20825
rect 6822 20816 6828 20828
rect 6880 20816 6886 20868
rect 7006 20816 7012 20868
rect 7064 20856 7070 20868
rect 7837 20859 7895 20865
rect 7837 20856 7849 20859
rect 7064 20828 7849 20856
rect 7064 20816 7070 20828
rect 7837 20825 7849 20828
rect 7883 20825 7895 20859
rect 7837 20819 7895 20825
rect 4614 20748 4620 20800
rect 4672 20788 4678 20800
rect 4801 20791 4859 20797
rect 4801 20788 4813 20791
rect 4672 20760 4813 20788
rect 4672 20748 4678 20760
rect 4801 20757 4813 20760
rect 4847 20757 4859 20791
rect 4801 20751 4859 20757
rect 10042 20748 10048 20800
rect 10100 20788 10106 20800
rect 11609 20791 11667 20797
rect 11609 20788 11621 20791
rect 10100 20760 11621 20788
rect 10100 20748 10106 20760
rect 11609 20757 11621 20760
rect 11655 20757 11667 20791
rect 12526 20788 12532 20800
rect 12487 20760 12532 20788
rect 11609 20751 11667 20757
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 5813 20587 5871 20593
rect 5813 20553 5825 20587
rect 5859 20584 5871 20587
rect 5902 20584 5908 20596
rect 5859 20556 5908 20584
rect 5859 20553 5871 20556
rect 5813 20547 5871 20553
rect 5902 20544 5908 20556
rect 5960 20584 5966 20596
rect 6730 20584 6736 20596
rect 5960 20556 6736 20584
rect 5960 20544 5966 20556
rect 6730 20544 6736 20556
rect 6788 20584 6794 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 6788 20556 8217 20584
rect 6788 20544 6794 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 8205 20547 8263 20553
rect 8294 20544 8300 20596
rect 8352 20584 8358 20596
rect 8481 20587 8539 20593
rect 8481 20584 8493 20587
rect 8352 20556 8493 20584
rect 8352 20544 8358 20556
rect 8481 20553 8493 20556
rect 8527 20584 8539 20587
rect 9490 20584 9496 20596
rect 8527 20556 9496 20584
rect 8527 20553 8539 20556
rect 8481 20547 8539 20553
rect 9490 20544 9496 20556
rect 9548 20544 9554 20596
rect 10134 20584 10140 20596
rect 9784 20556 10140 20584
rect 6822 20448 6828 20460
rect 6783 20420 6828 20448
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 9784 20457 9812 20556
rect 10134 20544 10140 20556
rect 10192 20584 10198 20596
rect 10962 20584 10968 20596
rect 10192 20556 10968 20584
rect 10192 20544 10198 20556
rect 10962 20544 10968 20556
rect 11020 20584 11026 20596
rect 11146 20584 11152 20596
rect 11020 20556 11152 20584
rect 11020 20544 11026 20556
rect 11146 20544 11152 20556
rect 11204 20544 11210 20596
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20448 9367 20451
rect 9769 20451 9827 20457
rect 9769 20448 9781 20451
rect 9355 20420 9781 20448
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 9769 20417 9781 20420
rect 9815 20417 9827 20451
rect 9769 20411 9827 20417
rect 12526 20408 12532 20460
rect 12584 20448 12590 20460
rect 12897 20451 12955 20457
rect 12897 20448 12909 20451
rect 12584 20420 12909 20448
rect 12584 20408 12590 20420
rect 12897 20417 12909 20420
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20417 13047 20451
rect 12989 20411 13047 20417
rect 10042 20389 10048 20392
rect 9677 20383 9735 20389
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 10036 20380 10048 20389
rect 9723 20352 10048 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 10036 20343 10048 20352
rect 10042 20340 10048 20343
rect 10100 20340 10106 20392
rect 11146 20340 11152 20392
rect 11204 20380 11210 20392
rect 11425 20383 11483 20389
rect 11425 20380 11437 20383
rect 11204 20352 11437 20380
rect 11204 20340 11210 20352
rect 11425 20349 11437 20352
rect 11471 20349 11483 20383
rect 11425 20343 11483 20349
rect 12342 20340 12348 20392
rect 12400 20380 12406 20392
rect 13004 20380 13032 20411
rect 12400 20352 13032 20380
rect 12400 20340 12406 20352
rect 5810 20272 5816 20324
rect 5868 20312 5874 20324
rect 6454 20312 6460 20324
rect 5868 20284 6460 20312
rect 5868 20272 5874 20284
rect 6454 20272 6460 20284
rect 6512 20272 6518 20324
rect 6914 20272 6920 20324
rect 6972 20312 6978 20324
rect 7070 20315 7128 20321
rect 7070 20312 7082 20315
rect 6972 20284 7082 20312
rect 6972 20272 6978 20284
rect 7070 20281 7082 20284
rect 7116 20281 7128 20315
rect 7070 20275 7128 20281
rect 11885 20315 11943 20321
rect 11885 20281 11897 20315
rect 11931 20312 11943 20315
rect 12066 20312 12072 20324
rect 11931 20284 12072 20312
rect 11931 20281 11943 20284
rect 11885 20275 11943 20281
rect 12066 20272 12072 20284
rect 12124 20312 12130 20324
rect 12805 20315 12863 20321
rect 12805 20312 12817 20315
rect 12124 20284 12817 20312
rect 12124 20272 12130 20284
rect 12805 20281 12817 20284
rect 12851 20281 12863 20315
rect 12805 20275 12863 20281
rect 5902 20204 5908 20256
rect 5960 20244 5966 20256
rect 6086 20244 6092 20256
rect 5960 20216 6092 20244
rect 5960 20204 5966 20216
rect 6086 20204 6092 20216
rect 6144 20204 6150 20256
rect 10962 20204 10968 20256
rect 11020 20244 11026 20256
rect 11149 20247 11207 20253
rect 11149 20244 11161 20247
rect 11020 20216 11161 20244
rect 11020 20204 11026 20216
rect 11149 20213 11161 20216
rect 11195 20213 11207 20247
rect 11149 20207 11207 20213
rect 12253 20247 12311 20253
rect 12253 20213 12265 20247
rect 12299 20244 12311 20247
rect 12342 20244 12348 20256
rect 12299 20216 12348 20244
rect 12299 20213 12311 20216
rect 12253 20207 12311 20213
rect 12342 20204 12348 20216
rect 12400 20204 12406 20256
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 12492 20216 12537 20244
rect 12492 20204 12498 20216
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 6822 20000 6828 20052
rect 6880 20040 6886 20052
rect 7193 20043 7251 20049
rect 7193 20040 7205 20043
rect 6880 20012 7205 20040
rect 6880 20000 6886 20012
rect 7193 20009 7205 20012
rect 7239 20009 7251 20043
rect 7193 20003 7251 20009
rect 8297 20043 8355 20049
rect 8297 20009 8309 20043
rect 8343 20040 8355 20043
rect 8386 20040 8392 20052
rect 8343 20012 8392 20040
rect 8343 20009 8355 20012
rect 8297 20003 8355 20009
rect 8386 20000 8392 20012
rect 8444 20000 8450 20052
rect 10321 20043 10379 20049
rect 10321 20009 10333 20043
rect 10367 20040 10379 20043
rect 10502 20040 10508 20052
rect 10367 20012 10508 20040
rect 10367 20009 10379 20012
rect 10321 20003 10379 20009
rect 10502 20000 10508 20012
rect 10560 20040 10566 20052
rect 12342 20040 12348 20052
rect 10560 20012 12348 20040
rect 10560 20000 10566 20012
rect 12342 20000 12348 20012
rect 12400 20040 12406 20052
rect 12529 20043 12587 20049
rect 12529 20040 12541 20043
rect 12400 20012 12541 20040
rect 12400 20000 12406 20012
rect 12529 20009 12541 20012
rect 12575 20009 12587 20043
rect 12529 20003 12587 20009
rect 9950 19904 9956 19916
rect 9911 19876 9956 19904
rect 9950 19864 9956 19876
rect 10008 19864 10014 19916
rect 11238 19864 11244 19916
rect 11296 19904 11302 19916
rect 11405 19907 11463 19913
rect 11405 19904 11417 19907
rect 11296 19876 11417 19904
rect 11296 19864 11302 19876
rect 11405 19873 11417 19876
rect 11451 19873 11463 19907
rect 11405 19867 11463 19873
rect 11146 19836 11152 19848
rect 11107 19808 11152 19836
rect 11146 19796 11152 19808
rect 11204 19796 11210 19848
rect 2774 19700 2780 19712
rect 2735 19672 2780 19700
rect 2774 19660 2780 19672
rect 2832 19660 2838 19712
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 5258 19700 5264 19712
rect 5123 19672 5264 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 6914 19700 6920 19712
rect 6875 19672 6920 19700
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 7929 19703 7987 19709
rect 7929 19669 7941 19703
rect 7975 19700 7987 19703
rect 8202 19700 8208 19712
rect 7975 19672 8208 19700
rect 7975 19669 7987 19672
rect 7929 19663 7987 19669
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 10502 19660 10508 19712
rect 10560 19700 10566 19712
rect 10597 19703 10655 19709
rect 10597 19700 10609 19703
rect 10560 19672 10609 19700
rect 10560 19660 10566 19672
rect 10597 19669 10609 19672
rect 10643 19669 10655 19703
rect 10597 19663 10655 19669
rect 12897 19703 12955 19709
rect 12897 19669 12909 19703
rect 12943 19700 12955 19703
rect 12986 19700 12992 19712
rect 12943 19672 12992 19700
rect 12943 19669 12955 19672
rect 12897 19663 12955 19669
rect 12986 19660 12992 19672
rect 13044 19660 13050 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 9953 19499 10011 19505
rect 9953 19465 9965 19499
rect 9999 19496 10011 19499
rect 10042 19496 10048 19508
rect 9999 19468 10048 19496
rect 9999 19465 10011 19468
rect 9953 19459 10011 19465
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 12437 19499 12495 19505
rect 12437 19465 12449 19499
rect 12483 19496 12495 19499
rect 12526 19496 12532 19508
rect 12483 19468 12532 19496
rect 12483 19465 12495 19468
rect 12437 19459 12495 19465
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 4246 19388 4252 19440
rect 4304 19428 4310 19440
rect 4798 19428 4804 19440
rect 4304 19400 4804 19428
rect 4304 19388 4310 19400
rect 4798 19388 4804 19400
rect 4856 19388 4862 19440
rect 10060 19428 10088 19456
rect 10060 19400 10640 19428
rect 2774 19360 2780 19372
rect 2735 19332 2780 19360
rect 2774 19320 2780 19332
rect 2832 19320 2838 19372
rect 5537 19363 5595 19369
rect 5537 19360 5549 19363
rect 4540 19332 5549 19360
rect 2685 19227 2743 19233
rect 2685 19193 2697 19227
rect 2731 19224 2743 19227
rect 3044 19227 3102 19233
rect 3044 19224 3056 19227
rect 2731 19196 3056 19224
rect 2731 19193 2743 19196
rect 2685 19187 2743 19193
rect 3044 19193 3056 19196
rect 3090 19224 3102 19227
rect 4540 19224 4568 19332
rect 5537 19329 5549 19332
rect 5583 19329 5595 19363
rect 10502 19360 10508 19372
rect 10463 19332 10508 19360
rect 5537 19323 5595 19329
rect 10502 19320 10508 19332
rect 10560 19320 10566 19372
rect 10612 19369 10640 19400
rect 10597 19363 10655 19369
rect 10597 19329 10609 19363
rect 10643 19329 10655 19363
rect 10597 19323 10655 19329
rect 11238 19320 11244 19372
rect 11296 19360 11302 19372
rect 12526 19360 12532 19372
rect 11296 19332 12532 19360
rect 11296 19320 11302 19332
rect 12526 19320 12532 19332
rect 12584 19360 12590 19372
rect 12986 19360 12992 19372
rect 12584 19332 12992 19360
rect 12584 19320 12590 19332
rect 12986 19320 12992 19332
rect 13044 19320 13050 19372
rect 9950 19252 9956 19304
rect 10008 19292 10014 19304
rect 10413 19295 10471 19301
rect 10413 19292 10425 19295
rect 10008 19264 10425 19292
rect 10008 19252 10014 19264
rect 10413 19261 10425 19264
rect 10459 19261 10471 19295
rect 10413 19255 10471 19261
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 11112 19264 12173 19292
rect 11112 19252 11118 19264
rect 12161 19261 12173 19264
rect 12207 19292 12219 19295
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12207 19264 12817 19292
rect 12207 19261 12219 19264
rect 12161 19255 12219 19261
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 3090 19196 4568 19224
rect 3090 19193 3102 19196
rect 3044 19187 3102 19193
rect 4540 19168 4568 19196
rect 4893 19227 4951 19233
rect 4893 19193 4905 19227
rect 4939 19224 4951 19227
rect 5166 19224 5172 19236
rect 4939 19196 5172 19224
rect 4939 19193 4951 19196
rect 4893 19187 4951 19193
rect 5166 19184 5172 19196
rect 5224 19224 5230 19236
rect 5445 19227 5503 19233
rect 5445 19224 5457 19227
rect 5224 19196 5457 19224
rect 5224 19184 5230 19196
rect 5445 19193 5457 19196
rect 5491 19193 5503 19227
rect 5445 19187 5503 19193
rect 7469 19227 7527 19233
rect 7469 19193 7481 19227
rect 7515 19224 7527 19227
rect 7558 19224 7564 19236
rect 7515 19196 7564 19224
rect 7515 19193 7527 19196
rect 7469 19187 7527 19193
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 11790 19224 11796 19236
rect 11751 19196 11796 19224
rect 11790 19184 11796 19196
rect 11848 19184 11854 19236
rect 12618 19184 12624 19236
rect 12676 19224 12682 19236
rect 12897 19227 12955 19233
rect 12897 19224 12909 19227
rect 12676 19196 12909 19224
rect 12676 19184 12682 19196
rect 12897 19193 12909 19196
rect 12943 19193 12955 19227
rect 12897 19187 12955 19193
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 4157 19159 4215 19165
rect 4157 19156 4169 19159
rect 4120 19128 4169 19156
rect 4120 19116 4126 19128
rect 4157 19125 4169 19128
rect 4203 19125 4215 19159
rect 4522 19156 4528 19168
rect 4483 19128 4528 19156
rect 4157 19119 4215 19125
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 4982 19156 4988 19168
rect 4943 19128 4988 19156
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 5353 19159 5411 19165
rect 5353 19156 5365 19159
rect 5316 19128 5365 19156
rect 5316 19116 5322 19128
rect 5353 19125 5365 19128
rect 5399 19125 5411 19159
rect 5353 19119 5411 19125
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 7009 19159 7067 19165
rect 7009 19156 7021 19159
rect 6880 19128 7021 19156
rect 6880 19116 6886 19128
rect 7009 19125 7021 19128
rect 7055 19125 7067 19159
rect 7009 19119 7067 19125
rect 8754 19116 8760 19168
rect 8812 19156 8818 19168
rect 8849 19159 8907 19165
rect 8849 19156 8861 19159
rect 8812 19128 8861 19156
rect 8812 19116 8818 19128
rect 8849 19125 8861 19128
rect 8895 19125 8907 19159
rect 10042 19156 10048 19168
rect 10003 19128 10048 19156
rect 8849 19119 8907 19125
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 11238 19156 11244 19168
rect 11199 19128 11244 19156
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 4982 18912 4988 18964
rect 5040 18952 5046 18964
rect 5442 18952 5448 18964
rect 5040 18924 5448 18952
rect 5040 18912 5046 18924
rect 5442 18912 5448 18924
rect 5500 18952 5506 18964
rect 5905 18955 5963 18961
rect 5905 18952 5917 18955
rect 5500 18924 5917 18952
rect 5500 18912 5506 18924
rect 5905 18921 5917 18924
rect 5951 18921 5963 18955
rect 6730 18952 6736 18964
rect 6691 18924 6736 18952
rect 5905 18915 5963 18921
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 10318 18912 10324 18964
rect 10376 18952 10382 18964
rect 10594 18952 10600 18964
rect 10376 18924 10600 18952
rect 10376 18912 10382 18924
rect 10594 18912 10600 18924
rect 10652 18952 10658 18964
rect 10689 18955 10747 18961
rect 10689 18952 10701 18955
rect 10652 18924 10701 18952
rect 10652 18912 10658 18924
rect 10689 18921 10701 18924
rect 10735 18921 10747 18955
rect 10689 18915 10747 18921
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11425 18955 11483 18961
rect 11425 18952 11437 18955
rect 11204 18924 11437 18952
rect 11204 18912 11210 18924
rect 11425 18921 11437 18924
rect 11471 18921 11483 18955
rect 11425 18915 11483 18921
rect 11977 18955 12035 18961
rect 11977 18921 11989 18955
rect 12023 18952 12035 18955
rect 12066 18952 12072 18964
rect 12023 18924 12072 18952
rect 12023 18921 12035 18924
rect 11977 18915 12035 18921
rect 12066 18912 12072 18924
rect 12124 18912 12130 18964
rect 1670 18884 1676 18896
rect 1631 18856 1676 18884
rect 1670 18844 1676 18856
rect 1728 18844 1734 18896
rect 4246 18844 4252 18896
rect 4304 18884 4310 18896
rect 4494 18887 4552 18893
rect 4494 18884 4506 18887
rect 4304 18856 4506 18884
rect 4304 18844 4310 18856
rect 4494 18853 4506 18856
rect 4540 18853 4552 18887
rect 4494 18847 4552 18853
rect 4798 18844 4804 18896
rect 4856 18884 4862 18896
rect 10134 18884 10140 18896
rect 4856 18856 10140 18884
rect 4856 18844 4862 18856
rect 10134 18844 10140 18856
rect 10192 18844 10198 18896
rect 11330 18844 11336 18896
rect 11388 18884 11394 18896
rect 11882 18884 11888 18896
rect 11388 18856 11888 18884
rect 11388 18844 11394 18856
rect 11882 18844 11888 18856
rect 11940 18884 11946 18896
rect 12437 18887 12495 18893
rect 12437 18884 12449 18887
rect 11940 18856 12449 18884
rect 11940 18844 11946 18856
rect 12437 18853 12449 18856
rect 12483 18853 12495 18887
rect 12437 18847 12495 18853
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 6641 18819 6699 18825
rect 6641 18785 6653 18819
rect 6687 18816 6699 18819
rect 7098 18816 7104 18828
rect 6687 18788 7104 18816
rect 6687 18785 6699 18788
rect 6641 18779 6699 18785
rect 7098 18776 7104 18788
rect 7156 18776 7162 18828
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 10594 18816 10600 18828
rect 10091 18788 10600 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 10594 18776 10600 18788
rect 10652 18816 10658 18828
rect 11514 18816 11520 18828
rect 10652 18788 11520 18816
rect 10652 18776 10658 18788
rect 11514 18776 11520 18788
rect 11572 18776 11578 18828
rect 12342 18816 12348 18828
rect 12303 18788 12348 18816
rect 12342 18776 12348 18788
rect 12400 18776 12406 18828
rect 3970 18708 3976 18760
rect 4028 18748 4034 18760
rect 4249 18751 4307 18757
rect 4249 18748 4261 18751
rect 4028 18720 4261 18748
rect 4028 18708 4034 18720
rect 4249 18717 4261 18720
rect 4295 18717 4307 18751
rect 7190 18748 7196 18760
rect 7151 18720 7196 18748
rect 4249 18711 4307 18717
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 7377 18751 7435 18757
rect 7377 18717 7389 18751
rect 7423 18748 7435 18751
rect 8202 18748 8208 18760
rect 7423 18720 8208 18748
rect 7423 18717 7435 18720
rect 7377 18711 7435 18717
rect 6638 18640 6644 18692
rect 6696 18680 6702 18692
rect 6914 18680 6920 18692
rect 6696 18652 6920 18680
rect 6696 18640 6702 18652
rect 6914 18640 6920 18652
rect 6972 18680 6978 18692
rect 7392 18680 7420 18711
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 9858 18748 9864 18760
rect 9732 18720 9864 18748
rect 9732 18708 9738 18720
rect 9858 18708 9864 18720
rect 9916 18708 9922 18760
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 10962 18748 10968 18760
rect 10367 18720 10968 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 6972 18652 7420 18680
rect 9125 18683 9183 18689
rect 6972 18640 6978 18652
rect 9125 18649 9137 18683
rect 9171 18680 9183 18683
rect 9582 18680 9588 18692
rect 9171 18652 9588 18680
rect 9171 18649 9183 18652
rect 9125 18643 9183 18649
rect 9582 18640 9588 18652
rect 9640 18640 9646 18692
rect 9950 18640 9956 18692
rect 10008 18680 10014 18692
rect 10336 18680 10364 18711
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 12526 18748 12532 18760
rect 12487 18720 12532 18748
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 10008 18652 10364 18680
rect 10008 18640 10014 18652
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 5629 18615 5687 18621
rect 5629 18612 5641 18615
rect 5592 18584 5641 18612
rect 5592 18572 5598 18584
rect 5629 18581 5641 18584
rect 5675 18581 5687 18615
rect 9674 18612 9680 18624
rect 9635 18584 9680 18612
rect 5629 18575 5687 18581
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 11054 18612 11060 18624
rect 11015 18584 11060 18612
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 6638 18408 6644 18420
rect 6599 18380 6644 18408
rect 6638 18368 6644 18380
rect 6696 18368 6702 18420
rect 7190 18368 7196 18420
rect 7248 18408 7254 18420
rect 7834 18408 7840 18420
rect 7248 18380 7840 18408
rect 7248 18368 7254 18380
rect 7834 18368 7840 18380
rect 7892 18408 7898 18420
rect 8481 18411 8539 18417
rect 8481 18408 8493 18411
rect 7892 18380 8493 18408
rect 7892 18368 7898 18380
rect 8481 18377 8493 18380
rect 8527 18377 8539 18411
rect 10134 18408 10140 18420
rect 10095 18380 10140 18408
rect 8481 18371 8539 18377
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 10502 18368 10508 18420
rect 10560 18408 10566 18420
rect 10597 18411 10655 18417
rect 10597 18408 10609 18411
rect 10560 18380 10609 18408
rect 10560 18368 10566 18380
rect 10597 18377 10609 18380
rect 10643 18377 10655 18411
rect 10597 18371 10655 18377
rect 4154 18300 4160 18352
rect 4212 18340 4218 18352
rect 5077 18343 5135 18349
rect 5077 18340 5089 18343
rect 4212 18312 5089 18340
rect 4212 18300 4218 18312
rect 5077 18309 5089 18312
rect 5123 18309 5135 18343
rect 8202 18340 8208 18352
rect 8163 18312 8208 18340
rect 5077 18303 5135 18309
rect 8202 18300 8208 18312
rect 8260 18300 8266 18352
rect 10152 18340 10180 18368
rect 10686 18340 10692 18352
rect 10152 18312 10692 18340
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 1578 18272 1584 18284
rect 1539 18244 1584 18272
rect 1578 18232 1584 18244
rect 1636 18232 1642 18284
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 4908 18244 5641 18272
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18173 1455 18207
rect 1397 18167 1455 18173
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 2958 18204 2964 18216
rect 2915 18176 2964 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 1412 18136 1440 18167
rect 2958 18164 2964 18176
rect 3016 18204 3022 18216
rect 3970 18204 3976 18216
rect 3016 18176 3976 18204
rect 3016 18164 3022 18176
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 2222 18136 2228 18148
rect 1412 18108 2228 18136
rect 2222 18096 2228 18108
rect 2280 18096 2286 18148
rect 2777 18139 2835 18145
rect 2777 18105 2789 18139
rect 2823 18136 2835 18139
rect 3050 18136 3056 18148
rect 2823 18108 3056 18136
rect 2823 18105 2835 18108
rect 2777 18099 2835 18105
rect 3050 18096 3056 18108
rect 3108 18145 3114 18148
rect 3108 18139 3172 18145
rect 3108 18105 3126 18139
rect 3160 18136 3172 18139
rect 4062 18136 4068 18148
rect 3160 18108 4068 18136
rect 3160 18105 3172 18108
rect 3108 18099 3172 18105
rect 3108 18096 3114 18099
rect 4062 18096 4068 18108
rect 4120 18136 4126 18148
rect 4908 18145 4936 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 9582 18272 9588 18284
rect 9543 18244 9588 18272
rect 5629 18235 5687 18241
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 11149 18275 11207 18281
rect 11149 18272 11161 18275
rect 10376 18244 11161 18272
rect 10376 18232 10382 18244
rect 11149 18241 11161 18244
rect 11195 18241 11207 18275
rect 11149 18235 11207 18241
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18272 11759 18275
rect 12342 18272 12348 18284
rect 11747 18244 12348 18272
rect 11747 18241 11759 18244
rect 11701 18235 11759 18241
rect 12342 18232 12348 18244
rect 12400 18272 12406 18284
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 12400 18244 12449 18272
rect 12400 18232 12406 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 5442 18204 5448 18216
rect 5403 18176 5448 18204
rect 5442 18164 5448 18176
rect 5500 18164 5506 18216
rect 6822 18204 6828 18216
rect 6783 18176 6828 18204
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 8294 18164 8300 18216
rect 8352 18204 8358 18216
rect 8570 18204 8576 18216
rect 8352 18176 8576 18204
rect 8352 18164 8358 18176
rect 8570 18164 8576 18176
rect 8628 18204 8634 18216
rect 9493 18207 9551 18213
rect 9493 18204 9505 18207
rect 8628 18176 9505 18204
rect 8628 18164 8634 18176
rect 9493 18173 9505 18176
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 12250 18164 12256 18216
rect 12308 18204 12314 18216
rect 13906 18204 13912 18216
rect 12308 18176 13912 18204
rect 12308 18164 12314 18176
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 4893 18139 4951 18145
rect 4893 18136 4905 18139
rect 4120 18108 4905 18136
rect 4120 18096 4126 18108
rect 4893 18105 4905 18108
rect 4939 18105 4951 18139
rect 4893 18099 4951 18105
rect 6273 18139 6331 18145
rect 6273 18105 6285 18139
rect 6319 18136 6331 18139
rect 7070 18139 7128 18145
rect 7070 18136 7082 18139
rect 6319 18108 7082 18136
rect 6319 18105 6331 18108
rect 6273 18099 6331 18105
rect 7070 18105 7082 18108
rect 7116 18136 7128 18139
rect 8110 18136 8116 18148
rect 7116 18108 8116 18136
rect 7116 18105 7128 18108
rect 7070 18099 7128 18105
rect 8110 18096 8116 18108
rect 8168 18096 8174 18148
rect 8849 18139 8907 18145
rect 8849 18105 8861 18139
rect 8895 18136 8907 18139
rect 8895 18108 9352 18136
rect 8895 18105 8907 18108
rect 8849 18099 8907 18105
rect 9324 18080 9352 18108
rect 10226 18096 10232 18148
rect 10284 18136 10290 18148
rect 11054 18136 11060 18148
rect 10284 18108 11060 18136
rect 10284 18096 10290 18108
rect 11054 18096 11060 18108
rect 11112 18096 11118 18148
rect 11882 18096 11888 18148
rect 11940 18096 11946 18148
rect 4246 18068 4252 18080
rect 4207 18040 4252 18068
rect 4246 18028 4252 18040
rect 4304 18068 4310 18080
rect 4525 18071 4583 18077
rect 4525 18068 4537 18071
rect 4304 18040 4537 18068
rect 4304 18028 4310 18040
rect 4525 18037 4537 18040
rect 4571 18037 4583 18071
rect 4525 18031 4583 18037
rect 5442 18028 5448 18080
rect 5500 18068 5506 18080
rect 5537 18071 5595 18077
rect 5537 18068 5549 18071
rect 5500 18040 5549 18068
rect 5500 18028 5506 18040
rect 5537 18037 5549 18040
rect 5583 18037 5595 18071
rect 5537 18031 5595 18037
rect 8938 18028 8944 18080
rect 8996 18068 9002 18080
rect 9033 18071 9091 18077
rect 9033 18068 9045 18071
rect 8996 18040 9045 18068
rect 8996 18028 9002 18040
rect 9033 18037 9045 18040
rect 9079 18037 9091 18071
rect 9033 18031 9091 18037
rect 9306 18028 9312 18080
rect 9364 18068 9370 18080
rect 9401 18071 9459 18077
rect 9401 18068 9413 18071
rect 9364 18040 9413 18068
rect 9364 18028 9370 18040
rect 9401 18037 9413 18040
rect 9447 18037 9459 18071
rect 9401 18031 9459 18037
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 10042 18068 10048 18080
rect 9916 18040 10048 18068
rect 9916 18028 9922 18040
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 10502 18068 10508 18080
rect 10463 18040 10508 18068
rect 10502 18028 10508 18040
rect 10560 18028 10566 18080
rect 10962 18068 10968 18080
rect 10923 18040 10968 18068
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 11422 18028 11428 18080
rect 11480 18068 11486 18080
rect 11900 18068 11928 18096
rect 11977 18071 12035 18077
rect 11977 18068 11989 18071
rect 11480 18040 11989 18068
rect 11480 18028 11486 18040
rect 11977 18037 11989 18040
rect 12023 18037 12035 18071
rect 11977 18031 12035 18037
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 1394 17824 1400 17876
rect 1452 17864 1458 17876
rect 1581 17867 1639 17873
rect 1581 17864 1593 17867
rect 1452 17836 1593 17864
rect 1452 17824 1458 17836
rect 1581 17833 1593 17836
rect 1627 17833 1639 17867
rect 1581 17827 1639 17833
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2777 17867 2835 17873
rect 2777 17864 2789 17867
rect 1820 17836 2789 17864
rect 1820 17824 1826 17836
rect 2777 17833 2789 17836
rect 2823 17864 2835 17867
rect 4062 17864 4068 17876
rect 2823 17836 4068 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 4341 17867 4399 17873
rect 4341 17833 4353 17867
rect 4387 17864 4399 17867
rect 5258 17864 5264 17876
rect 4387 17836 5264 17864
rect 4387 17833 4399 17836
rect 4341 17827 4399 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 7561 17867 7619 17873
rect 7561 17864 7573 17867
rect 7156 17836 7573 17864
rect 7156 17824 7162 17836
rect 7561 17833 7573 17836
rect 7607 17833 7619 17867
rect 11054 17864 11060 17876
rect 11015 17836 11060 17864
rect 7561 17827 7619 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 5534 17756 5540 17808
rect 5592 17805 5598 17808
rect 9950 17805 9956 17808
rect 5592 17799 5656 17805
rect 5592 17765 5610 17799
rect 5644 17765 5656 17799
rect 5592 17759 5656 17765
rect 9493 17799 9551 17805
rect 9493 17765 9505 17799
rect 9539 17796 9551 17799
rect 9944 17796 9956 17805
rect 9539 17768 9956 17796
rect 9539 17765 9551 17768
rect 9493 17759 9551 17765
rect 9944 17759 9956 17768
rect 5592 17756 5598 17759
rect 9950 17756 9956 17759
rect 10008 17756 10014 17808
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 4614 17728 4620 17740
rect 2832 17700 4620 17728
rect 2832 17688 2838 17700
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 5261 17731 5319 17737
rect 5261 17697 5273 17731
rect 5307 17728 5319 17731
rect 5442 17728 5448 17740
rect 5307 17700 5448 17728
rect 5307 17697 5319 17700
rect 5261 17691 5319 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 7926 17728 7932 17740
rect 7887 17700 7932 17728
rect 7926 17688 7932 17700
rect 7984 17688 7990 17740
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17728 8079 17731
rect 8938 17728 8944 17740
rect 8067 17700 8944 17728
rect 8067 17697 8079 17700
rect 8021 17691 8079 17697
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17728 9735 17731
rect 9766 17728 9772 17740
rect 9723 17700 9772 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 2866 17660 2872 17672
rect 2827 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 2958 17620 2964 17672
rect 3016 17660 3022 17672
rect 4246 17660 4252 17672
rect 3016 17632 4252 17660
rect 3016 17620 3022 17632
rect 4246 17620 4252 17632
rect 4304 17620 4310 17672
rect 4890 17620 4896 17672
rect 4948 17660 4954 17672
rect 5166 17660 5172 17672
rect 4948 17632 5172 17660
rect 4948 17620 4954 17632
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 5353 17663 5411 17669
rect 5353 17629 5365 17663
rect 5399 17629 5411 17663
rect 8110 17660 8116 17672
rect 8071 17632 8116 17660
rect 5353 17623 5411 17629
rect 5368 17592 5396 17623
rect 8110 17620 8116 17632
rect 8168 17620 8174 17672
rect 8846 17620 8852 17672
rect 8904 17620 8910 17672
rect 4080 17564 5396 17592
rect 4080 17536 4108 17564
rect 7098 17552 7104 17604
rect 7156 17592 7162 17604
rect 8864 17592 8892 17620
rect 7156 17564 8892 17592
rect 7156 17552 7162 17564
rect 2406 17524 2412 17536
rect 2367 17496 2412 17524
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 3881 17527 3939 17533
rect 3881 17493 3893 17527
rect 3927 17524 3939 17527
rect 4062 17524 4068 17536
rect 3927 17496 4068 17524
rect 3927 17493 3939 17496
rect 3881 17487 3939 17493
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 4522 17484 4528 17536
rect 4580 17524 4586 17536
rect 4893 17527 4951 17533
rect 4893 17524 4905 17527
rect 4580 17496 4905 17524
rect 4580 17484 4586 17496
rect 4893 17493 4905 17496
rect 4939 17524 4951 17527
rect 4982 17524 4988 17536
rect 4939 17496 4988 17524
rect 4939 17493 4951 17496
rect 4893 17487 4951 17493
rect 4982 17484 4988 17496
rect 5040 17484 5046 17536
rect 6730 17524 6736 17536
rect 6691 17496 6736 17524
rect 6730 17484 6736 17496
rect 6788 17484 6794 17536
rect 7190 17524 7196 17536
rect 7151 17496 7196 17524
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 9033 17527 9091 17533
rect 9033 17524 9045 17527
rect 8628 17496 9045 17524
rect 8628 17484 8634 17496
rect 9033 17493 9045 17496
rect 9079 17493 9091 17527
rect 11330 17524 11336 17536
rect 11291 17496 11336 17524
rect 9033 17487 9091 17493
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 11882 17484 11888 17536
rect 11940 17524 11946 17536
rect 11977 17527 12035 17533
rect 11977 17524 11989 17527
rect 11940 17496 11989 17524
rect 11940 17484 11946 17496
rect 11977 17493 11989 17496
rect 12023 17493 12035 17527
rect 11977 17487 12035 17493
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 1762 17320 1768 17332
rect 1723 17292 1768 17320
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 2866 17320 2872 17332
rect 2827 17292 2872 17320
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 5442 17320 5448 17332
rect 4479 17292 5448 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 8110 17280 8116 17332
rect 8168 17320 8174 17332
rect 8481 17323 8539 17329
rect 8481 17320 8493 17323
rect 8168 17292 8493 17320
rect 8168 17280 8174 17292
rect 8481 17289 8493 17292
rect 8527 17289 8539 17323
rect 8846 17320 8852 17332
rect 8807 17292 8852 17320
rect 8481 17283 8539 17289
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9861 17323 9919 17329
rect 9861 17289 9873 17323
rect 9907 17320 9919 17323
rect 9950 17320 9956 17332
rect 9907 17292 9956 17320
rect 9907 17289 9919 17292
rect 9861 17283 9919 17289
rect 9950 17280 9956 17292
rect 10008 17280 10014 17332
rect 10594 17320 10600 17332
rect 10555 17292 10600 17320
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 10781 17323 10839 17329
rect 10781 17289 10793 17323
rect 10827 17320 10839 17323
rect 10962 17320 10968 17332
rect 10827 17292 10968 17320
rect 10827 17289 10839 17292
rect 10781 17283 10839 17289
rect 10962 17280 10968 17292
rect 11020 17320 11026 17332
rect 11330 17320 11336 17332
rect 11020 17292 11336 17320
rect 11020 17280 11026 17292
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 2501 17255 2559 17261
rect 2501 17221 2513 17255
rect 2547 17252 2559 17255
rect 2958 17252 2964 17264
rect 2547 17224 2964 17252
rect 2547 17221 2559 17224
rect 2501 17215 2559 17221
rect 2958 17212 2964 17224
rect 3016 17212 3022 17264
rect 9766 17212 9772 17264
rect 9824 17252 9830 17264
rect 11514 17252 11520 17264
rect 9824 17224 11520 17252
rect 9824 17212 9830 17224
rect 11514 17212 11520 17224
rect 11572 17252 11578 17264
rect 11793 17255 11851 17261
rect 11793 17252 11805 17255
rect 11572 17224 11805 17252
rect 11572 17212 11578 17224
rect 11793 17221 11805 17224
rect 11839 17221 11851 17255
rect 11793 17215 11851 17221
rect 3050 17144 3056 17196
rect 3108 17184 3114 17196
rect 3421 17187 3479 17193
rect 3421 17184 3433 17187
rect 3108 17156 3433 17184
rect 3108 17144 3114 17156
rect 3421 17153 3433 17156
rect 3467 17153 3479 17187
rect 4982 17184 4988 17196
rect 4943 17156 4988 17184
rect 3421 17147 3479 17153
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 10318 17144 10324 17196
rect 10376 17184 10382 17196
rect 11238 17184 11244 17196
rect 10376 17156 11244 17184
rect 10376 17144 10382 17156
rect 11238 17144 11244 17156
rect 11296 17184 11302 17196
rect 11333 17187 11391 17193
rect 11333 17184 11345 17187
rect 11296 17156 11345 17184
rect 11296 17144 11302 17156
rect 11333 17153 11345 17156
rect 11379 17184 11391 17187
rect 11882 17184 11888 17196
rect 11379 17156 11888 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 11882 17144 11888 17156
rect 11940 17184 11946 17196
rect 12066 17184 12072 17196
rect 11940 17156 12072 17184
rect 11940 17144 11946 17156
rect 12066 17144 12072 17156
rect 12124 17144 12130 17196
rect 2958 17076 2964 17128
rect 3016 17116 3022 17128
rect 4338 17116 4344 17128
rect 3016 17088 4016 17116
rect 4299 17088 4344 17116
rect 3016 17076 3022 17088
rect 2133 17051 2191 17057
rect 2133 17017 2145 17051
rect 2179 17048 2191 17051
rect 2498 17048 2504 17060
rect 2179 17020 2504 17048
rect 2179 17017 2191 17020
rect 2133 17011 2191 17017
rect 2498 17008 2504 17020
rect 2556 17048 2562 17060
rect 3988 17057 4016 17088
rect 4338 17076 4344 17088
rect 4396 17116 4402 17128
rect 4706 17116 4712 17128
rect 4396 17088 4712 17116
rect 4396 17076 4402 17088
rect 4706 17076 4712 17088
rect 4764 17116 4770 17128
rect 4801 17119 4859 17125
rect 4801 17116 4813 17119
rect 4764 17088 4813 17116
rect 4764 17076 4770 17088
rect 4801 17085 4813 17088
rect 4847 17085 4859 17119
rect 4801 17079 4859 17085
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17116 4951 17119
rect 5166 17116 5172 17128
rect 4939 17088 5172 17116
rect 4939 17085 4951 17088
rect 4893 17079 4951 17085
rect 3329 17051 3387 17057
rect 3329 17048 3341 17051
rect 2556 17020 3341 17048
rect 2556 17008 2562 17020
rect 3329 17017 3341 17020
rect 3375 17017 3387 17051
rect 3329 17011 3387 17017
rect 3973 17051 4031 17057
rect 3973 17017 3985 17051
rect 4019 17048 4031 17051
rect 4908 17048 4936 17079
rect 5166 17076 5172 17088
rect 5224 17076 5230 17128
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 7006 17116 7012 17128
rect 6687 17088 7012 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 7006 17076 7012 17088
rect 7064 17116 7070 17128
rect 7101 17119 7159 17125
rect 7101 17116 7113 17119
rect 7064 17088 7113 17116
rect 7064 17076 7070 17088
rect 7101 17085 7113 17088
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 9309 17119 9367 17125
rect 9309 17116 9321 17119
rect 8352 17088 9321 17116
rect 8352 17076 8358 17088
rect 9309 17085 9321 17088
rect 9355 17085 9367 17119
rect 9309 17079 9367 17085
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 10410 17116 10416 17128
rect 9824 17088 10416 17116
rect 9824 17076 9830 17088
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 10594 17076 10600 17128
rect 10652 17116 10658 17128
rect 11149 17119 11207 17125
rect 11149 17116 11161 17119
rect 10652 17088 11161 17116
rect 10652 17076 10658 17088
rect 11149 17085 11161 17088
rect 11195 17116 11207 17119
rect 12158 17116 12164 17128
rect 11195 17088 12164 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 12158 17076 12164 17088
rect 12216 17076 12222 17128
rect 5813 17051 5871 17057
rect 5813 17048 5825 17051
rect 4019 17020 4936 17048
rect 5000 17020 5825 17048
rect 4019 17017 4031 17020
rect 3973 17011 4031 17017
rect 3237 16983 3295 16989
rect 3237 16949 3249 16983
rect 3283 16980 3295 16983
rect 3602 16980 3608 16992
rect 3283 16952 3608 16980
rect 3283 16949 3295 16952
rect 3237 16943 3295 16949
rect 3602 16940 3608 16952
rect 3660 16940 3666 16992
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 5000 16980 5028 17020
rect 5813 17017 5825 17020
rect 5859 17048 5871 17051
rect 6822 17048 6828 17060
rect 5859 17020 6828 17048
rect 5859 17017 5871 17020
rect 5813 17011 5871 17017
rect 6822 17008 6828 17020
rect 6880 17008 6886 17060
rect 7190 17008 7196 17060
rect 7248 17048 7254 17060
rect 7368 17051 7426 17057
rect 7368 17048 7380 17051
rect 7248 17020 7380 17048
rect 7248 17008 7254 17020
rect 7368 17017 7380 17020
rect 7414 17048 7426 17051
rect 7742 17048 7748 17060
rect 7414 17020 7748 17048
rect 7414 17017 7426 17020
rect 7368 17011 7426 17017
rect 7742 17008 7748 17020
rect 7800 17008 7806 17060
rect 7926 17008 7932 17060
rect 7984 17048 7990 17060
rect 9125 17051 9183 17057
rect 9125 17048 9137 17051
rect 7984 17020 9137 17048
rect 7984 17008 7990 17020
rect 9125 17017 9137 17020
rect 9171 17017 9183 17051
rect 9125 17011 9183 17017
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 12618 17048 12624 17060
rect 10836 17020 12624 17048
rect 10836 17008 10842 17020
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 5534 16980 5540 16992
rect 4120 16952 5028 16980
rect 5495 16952 5540 16980
rect 4120 16940 4126 16952
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 10318 16980 10324 16992
rect 10279 16952 10324 16980
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 11238 16940 11244 16992
rect 11296 16980 11302 16992
rect 11296 16952 11341 16980
rect 11296 16940 11302 16952
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16776 2559 16779
rect 2866 16776 2872 16788
rect 2547 16748 2872 16776
rect 2547 16745 2559 16748
rect 2501 16739 2559 16745
rect 2866 16736 2872 16748
rect 2924 16736 2930 16788
rect 2961 16779 3019 16785
rect 2961 16745 2973 16779
rect 3007 16776 3019 16779
rect 3050 16776 3056 16788
rect 3007 16748 3056 16776
rect 3007 16745 3019 16748
rect 2961 16739 3019 16745
rect 3050 16736 3056 16748
rect 3108 16736 3114 16788
rect 3237 16779 3295 16785
rect 3237 16745 3249 16779
rect 3283 16776 3295 16779
rect 3602 16776 3608 16788
rect 3283 16748 3608 16776
rect 3283 16745 3295 16748
rect 3237 16739 3295 16745
rect 3602 16736 3608 16748
rect 3660 16776 3666 16788
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 3660 16748 4077 16776
rect 3660 16736 3666 16748
rect 4065 16745 4077 16748
rect 4111 16745 4123 16779
rect 4065 16739 4123 16745
rect 4154 16736 4160 16788
rect 4212 16776 4218 16788
rect 4433 16779 4491 16785
rect 4433 16776 4445 16779
rect 4212 16748 4445 16776
rect 4212 16736 4218 16748
rect 4433 16745 4445 16748
rect 4479 16776 4491 16779
rect 4614 16776 4620 16788
rect 4479 16748 4620 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 5261 16779 5319 16785
rect 5261 16745 5273 16779
rect 5307 16776 5319 16779
rect 5718 16776 5724 16788
rect 5307 16748 5724 16776
rect 5307 16745 5319 16748
rect 5261 16739 5319 16745
rect 5718 16736 5724 16748
rect 5776 16776 5782 16788
rect 6730 16776 6736 16788
rect 5776 16748 6736 16776
rect 5776 16736 5782 16748
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 7834 16776 7840 16788
rect 7795 16748 7840 16776
rect 7834 16736 7840 16748
rect 7892 16736 7898 16788
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 8846 16776 8852 16788
rect 8720 16748 8852 16776
rect 8720 16736 8726 16748
rect 8846 16736 8852 16748
rect 8904 16736 8910 16788
rect 8941 16779 8999 16785
rect 8941 16745 8953 16779
rect 8987 16776 8999 16779
rect 9582 16776 9588 16788
rect 8987 16748 9588 16776
rect 8987 16745 8999 16748
rect 8941 16739 8999 16745
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 10226 16776 10232 16788
rect 10187 16748 10232 16776
rect 10226 16736 10232 16748
rect 10284 16736 10290 16788
rect 11238 16776 11244 16788
rect 11199 16748 11244 16776
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 13173 16779 13231 16785
rect 13173 16776 13185 16779
rect 12124 16748 13185 16776
rect 12124 16736 12130 16748
rect 13173 16745 13185 16748
rect 13219 16745 13231 16779
rect 13173 16739 13231 16745
rect 3970 16668 3976 16720
rect 4028 16708 4034 16720
rect 4525 16711 4583 16717
rect 4525 16708 4537 16711
rect 4028 16680 4537 16708
rect 4028 16668 4034 16680
rect 4525 16677 4537 16680
rect 4571 16677 4583 16711
rect 4525 16671 4583 16677
rect 6178 16668 6184 16720
rect 6236 16708 6242 16720
rect 6365 16711 6423 16717
rect 6365 16708 6377 16711
rect 6236 16680 6377 16708
rect 6236 16668 6242 16680
rect 6365 16677 6377 16680
rect 6411 16677 6423 16711
rect 6365 16671 6423 16677
rect 7653 16711 7711 16717
rect 7653 16677 7665 16711
rect 7699 16708 7711 16711
rect 8110 16708 8116 16720
rect 7699 16680 8116 16708
rect 7699 16677 7711 16680
rect 7653 16671 7711 16677
rect 6270 16640 6276 16652
rect 6231 16612 6276 16640
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 4154 16532 4160 16584
rect 4212 16572 4218 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4212 16544 4629 16572
rect 4212 16532 4218 16544
rect 4617 16541 4629 16544
rect 4663 16572 4675 16575
rect 4982 16572 4988 16584
rect 4663 16544 4988 16572
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 4982 16532 4988 16544
rect 5040 16532 5046 16584
rect 5902 16532 5908 16584
rect 5960 16532 5966 16584
rect 6549 16575 6607 16581
rect 6549 16541 6561 16575
rect 6595 16572 6607 16575
rect 6638 16572 6644 16584
rect 6595 16544 6644 16572
rect 6595 16541 6607 16544
rect 6549 16535 6607 16541
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 8036 16572 8064 16680
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 10137 16711 10195 16717
rect 10137 16677 10149 16711
rect 10183 16708 10195 16711
rect 10183 16680 10732 16708
rect 10183 16677 10195 16680
rect 10137 16671 10195 16677
rect 10704 16652 10732 16680
rect 8202 16640 8208 16652
rect 8163 16612 8208 16640
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16640 8355 16643
rect 8662 16640 8668 16652
rect 8343 16612 8668 16640
rect 8343 16609 8355 16612
rect 8297 16603 8355 16609
rect 8662 16600 8668 16612
rect 8720 16640 8726 16652
rect 9217 16643 9275 16649
rect 9217 16640 9229 16643
rect 8720 16612 9229 16640
rect 8720 16600 8726 16612
rect 9217 16609 9229 16612
rect 9263 16609 9275 16643
rect 10594 16640 10600 16652
rect 10555 16612 10600 16640
rect 9217 16603 9275 16609
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 10744 16612 10789 16640
rect 10744 16600 10750 16612
rect 11514 16600 11520 16652
rect 11572 16640 11578 16652
rect 11793 16643 11851 16649
rect 11793 16640 11805 16643
rect 11572 16612 11805 16640
rect 11572 16600 11578 16612
rect 11793 16609 11805 16612
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 12049 16643 12107 16649
rect 12049 16640 12061 16643
rect 11940 16612 12061 16640
rect 11940 16600 11946 16612
rect 12049 16609 12061 16612
rect 12095 16609 12107 16643
rect 12049 16603 12107 16609
rect 8386 16572 8392 16584
rect 8036 16544 8392 16572
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 10318 16532 10324 16584
rect 10376 16572 10382 16584
rect 10781 16575 10839 16581
rect 10781 16572 10793 16575
rect 10376 16544 10793 16572
rect 10376 16532 10382 16544
rect 10781 16541 10793 16544
rect 10827 16541 10839 16575
rect 10781 16535 10839 16541
rect 4522 16464 4528 16516
rect 4580 16504 4586 16516
rect 5920 16504 5948 16532
rect 4580 16476 5948 16504
rect 7193 16507 7251 16513
rect 4580 16464 4586 16476
rect 7193 16473 7205 16507
rect 7239 16504 7251 16507
rect 7466 16504 7472 16516
rect 7239 16476 7472 16504
rect 7239 16473 7251 16476
rect 7193 16467 7251 16473
rect 7466 16464 7472 16476
rect 7524 16504 7530 16516
rect 8478 16504 8484 16516
rect 7524 16476 8484 16504
rect 7524 16464 7530 16476
rect 8478 16464 8484 16476
rect 8536 16464 8542 16516
rect 5626 16436 5632 16448
rect 5587 16408 5632 16436
rect 5626 16396 5632 16408
rect 5684 16396 5690 16448
rect 5902 16436 5908 16448
rect 5863 16408 5908 16436
rect 5902 16396 5908 16408
rect 5960 16396 5966 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 3789 16235 3847 16241
rect 3789 16201 3801 16235
rect 3835 16232 3847 16235
rect 3970 16232 3976 16244
rect 3835 16204 3976 16232
rect 3835 16201 3847 16204
rect 3789 16195 3847 16201
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 4157 16235 4215 16241
rect 4157 16201 4169 16235
rect 4203 16232 4215 16235
rect 4614 16232 4620 16244
rect 4203 16204 4620 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 6178 16232 6184 16244
rect 6139 16204 6184 16232
rect 6178 16192 6184 16204
rect 6236 16232 6242 16244
rect 6730 16232 6736 16244
rect 6236 16204 6736 16232
rect 6236 16192 6242 16204
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 10781 16235 10839 16241
rect 10781 16201 10793 16235
rect 10827 16232 10839 16235
rect 11238 16232 11244 16244
rect 10827 16204 11244 16232
rect 10827 16201 10839 16204
rect 10781 16195 10839 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 11572 16204 12173 16232
rect 11572 16192 11578 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 5718 16096 5724 16108
rect 5679 16068 5724 16096
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 7650 16096 7656 16108
rect 7611 16068 7656 16096
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 8205 16099 8263 16105
rect 8205 16096 8217 16099
rect 7800 16068 8217 16096
rect 7800 16056 7806 16068
rect 8205 16065 8217 16068
rect 8251 16096 8263 16099
rect 8478 16096 8484 16108
rect 8251 16068 8484 16096
rect 8251 16065 8263 16068
rect 8205 16059 8263 16065
rect 8478 16056 8484 16068
rect 8536 16096 8542 16108
rect 9306 16096 9312 16108
rect 8536 16068 9312 16096
rect 8536 16056 8542 16068
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16096 10011 16099
rect 11146 16096 11152 16108
rect 9999 16068 11152 16096
rect 9999 16065 10011 16068
rect 9953 16059 10011 16065
rect 11146 16056 11152 16068
rect 11204 16096 11210 16108
rect 11333 16099 11391 16105
rect 11333 16096 11345 16099
rect 11204 16068 11345 16096
rect 11204 16056 11210 16068
rect 11333 16065 11345 16068
rect 11379 16096 11391 16099
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 11379 16068 11805 16096
rect 11379 16065 11391 16068
rect 11333 16059 11391 16065
rect 11793 16065 11805 16068
rect 11839 16096 11851 16099
rect 11882 16096 11888 16108
rect 11839 16068 11888 16096
rect 11839 16065 11851 16068
rect 11793 16059 11851 16065
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 5166 15988 5172 16040
rect 5224 16028 5230 16040
rect 5537 16031 5595 16037
rect 5537 16028 5549 16031
rect 5224 16000 5549 16028
rect 5224 15988 5230 16000
rect 5537 15997 5549 16000
rect 5583 16028 5595 16031
rect 5902 16028 5908 16040
rect 5583 16000 5908 16028
rect 5583 15997 5595 16000
rect 5537 15991 5595 15997
rect 5902 15988 5908 16000
rect 5960 15988 5966 16040
rect 7466 16028 7472 16040
rect 7427 16000 7472 16028
rect 7466 15988 7472 16000
rect 7524 15988 7530 16040
rect 7558 15988 7564 16040
rect 7616 16028 7622 16040
rect 8018 16028 8024 16040
rect 7616 16000 8024 16028
rect 7616 15988 7622 16000
rect 8018 15988 8024 16000
rect 8076 15988 8082 16040
rect 9125 16031 9183 16037
rect 9125 15997 9137 16031
rect 9171 16028 9183 16031
rect 9582 16028 9588 16040
rect 9171 16000 9588 16028
rect 9171 15997 9183 16000
rect 9125 15991 9183 15997
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 5077 15963 5135 15969
rect 5077 15929 5089 15963
rect 5123 15960 5135 15963
rect 5350 15960 5356 15972
rect 5123 15932 5356 15960
rect 5123 15929 5135 15932
rect 5077 15923 5135 15929
rect 5350 15920 5356 15932
rect 5408 15920 5414 15972
rect 6270 15920 6276 15972
rect 6328 15960 6334 15972
rect 6641 15963 6699 15969
rect 6641 15960 6653 15963
rect 6328 15932 6653 15960
rect 6328 15920 6334 15932
rect 6641 15929 6653 15932
rect 6687 15960 6699 15963
rect 7190 15960 7196 15972
rect 6687 15932 7196 15960
rect 6687 15929 6699 15932
rect 6641 15923 6699 15929
rect 7190 15920 7196 15932
rect 7248 15920 7254 15972
rect 8573 15963 8631 15969
rect 8573 15960 8585 15963
rect 8036 15932 8585 15960
rect 8036 15904 8064 15932
rect 8573 15929 8585 15932
rect 8619 15960 8631 15963
rect 8846 15960 8852 15972
rect 8619 15932 8852 15960
rect 8619 15929 8631 15932
rect 8573 15923 8631 15929
rect 8846 15920 8852 15932
rect 8904 15960 8910 15972
rect 9033 15963 9091 15969
rect 9033 15960 9045 15963
rect 8904 15932 9045 15960
rect 8904 15920 8910 15932
rect 9033 15929 9045 15932
rect 9079 15929 9091 15963
rect 9033 15923 9091 15929
rect 10321 15963 10379 15969
rect 10321 15929 10333 15963
rect 10367 15960 10379 15963
rect 11149 15963 11207 15969
rect 11149 15960 11161 15963
rect 10367 15932 11161 15960
rect 10367 15929 10379 15932
rect 10321 15923 10379 15929
rect 11149 15929 11161 15932
rect 11195 15960 11207 15963
rect 11330 15960 11336 15972
rect 11195 15932 11336 15960
rect 11195 15929 11207 15932
rect 11149 15923 11207 15929
rect 11330 15920 11336 15932
rect 11388 15920 11394 15972
rect 4154 15852 4160 15904
rect 4212 15892 4218 15904
rect 4433 15895 4491 15901
rect 4433 15892 4445 15895
rect 4212 15864 4445 15892
rect 4212 15852 4218 15864
rect 4433 15861 4445 15864
rect 4479 15861 4491 15895
rect 4433 15855 4491 15861
rect 5169 15895 5227 15901
rect 5169 15861 5181 15895
rect 5215 15892 5227 15895
rect 5442 15892 5448 15904
rect 5215 15864 5448 15892
rect 5215 15861 5227 15864
rect 5169 15855 5227 15861
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 5626 15892 5632 15904
rect 5539 15864 5632 15892
rect 5626 15852 5632 15864
rect 5684 15892 5690 15904
rect 5994 15892 6000 15904
rect 5684 15864 6000 15892
rect 5684 15852 5690 15864
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 8018 15852 8024 15904
rect 8076 15852 8082 15904
rect 8202 15852 8208 15904
rect 8260 15892 8266 15904
rect 8665 15895 8723 15901
rect 8665 15892 8677 15895
rect 8260 15864 8677 15892
rect 8260 15852 8266 15864
rect 8665 15861 8677 15864
rect 8711 15861 8723 15895
rect 8665 15855 8723 15861
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 10689 15895 10747 15901
rect 10689 15892 10701 15895
rect 10468 15864 10701 15892
rect 10468 15852 10474 15864
rect 10689 15861 10701 15864
rect 10735 15892 10747 15895
rect 11241 15895 11299 15901
rect 11241 15892 11253 15895
rect 10735 15864 11253 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 11241 15861 11253 15864
rect 11287 15892 11299 15895
rect 12250 15892 12256 15904
rect 11287 15864 12256 15892
rect 11287 15861 11299 15864
rect 11241 15855 11299 15861
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 3970 15648 3976 15700
rect 4028 15688 4034 15700
rect 4065 15691 4123 15697
rect 4065 15688 4077 15691
rect 4028 15660 4077 15688
rect 4028 15648 4034 15660
rect 4065 15657 4077 15660
rect 4111 15657 4123 15691
rect 5166 15688 5172 15700
rect 5127 15660 5172 15688
rect 4065 15651 4123 15657
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5810 15648 5816 15700
rect 5868 15688 5874 15700
rect 5997 15691 6055 15697
rect 5997 15688 6009 15691
rect 5868 15660 6009 15688
rect 5868 15648 5874 15660
rect 5997 15657 6009 15660
rect 6043 15688 6055 15691
rect 6178 15688 6184 15700
rect 6043 15660 6184 15688
rect 6043 15657 6055 15660
rect 5997 15651 6055 15657
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 6822 15688 6828 15700
rect 6783 15660 6828 15688
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 7561 15691 7619 15697
rect 7561 15657 7573 15691
rect 7607 15688 7619 15691
rect 7650 15688 7656 15700
rect 7607 15660 7656 15688
rect 7607 15657 7619 15660
rect 7561 15651 7619 15657
rect 7650 15648 7656 15660
rect 7708 15648 7714 15700
rect 7837 15691 7895 15697
rect 7837 15657 7849 15691
rect 7883 15688 7895 15691
rect 7926 15688 7932 15700
rect 7883 15660 7932 15688
rect 7883 15657 7895 15660
rect 7837 15651 7895 15657
rect 7926 15648 7932 15660
rect 7984 15648 7990 15700
rect 8202 15688 8208 15700
rect 8163 15660 8208 15688
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8386 15648 8392 15700
rect 8444 15688 8450 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 8444 15660 8953 15688
rect 8444 15648 8450 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 8941 15651 8999 15657
rect 9953 15691 10011 15697
rect 9953 15657 9965 15691
rect 9999 15688 10011 15691
rect 10505 15691 10563 15697
rect 10505 15688 10517 15691
rect 9999 15660 10517 15688
rect 9999 15657 10011 15660
rect 9953 15651 10011 15657
rect 10505 15657 10517 15660
rect 10551 15688 10563 15691
rect 10594 15688 10600 15700
rect 10551 15660 10600 15688
rect 10551 15657 10563 15660
rect 10505 15651 10563 15657
rect 10594 15648 10600 15660
rect 10652 15648 10658 15700
rect 4430 15620 4436 15632
rect 4343 15592 4436 15620
rect 4430 15580 4436 15592
rect 4488 15620 4494 15632
rect 4706 15620 4712 15632
rect 4488 15592 4712 15620
rect 4488 15580 4494 15592
rect 4706 15580 4712 15592
rect 4764 15580 4770 15632
rect 5902 15580 5908 15632
rect 5960 15620 5966 15632
rect 6089 15623 6147 15629
rect 6089 15620 6101 15623
rect 5960 15592 6101 15620
rect 5960 15580 5966 15592
rect 6089 15589 6101 15592
rect 6135 15589 6147 15623
rect 6089 15583 6147 15589
rect 7098 15580 7104 15632
rect 7156 15620 7162 15632
rect 8846 15620 8852 15632
rect 7156 15592 8852 15620
rect 7156 15580 7162 15592
rect 8846 15580 8852 15592
rect 8904 15620 8910 15632
rect 9217 15623 9275 15629
rect 9217 15620 9229 15623
rect 8904 15592 9229 15620
rect 8904 15580 8910 15592
rect 9217 15589 9229 15592
rect 9263 15589 9275 15623
rect 10318 15620 10324 15632
rect 10279 15592 10324 15620
rect 9217 15583 9275 15589
rect 10318 15580 10324 15592
rect 10376 15580 10382 15632
rect 10873 15623 10931 15629
rect 10873 15589 10885 15623
rect 10919 15620 10931 15623
rect 10962 15620 10968 15632
rect 10919 15592 10968 15620
rect 10919 15589 10931 15592
rect 10873 15583 10931 15589
rect 10962 15580 10968 15592
rect 11020 15580 11026 15632
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 4525 15555 4583 15561
rect 4525 15552 4537 15555
rect 4304 15524 4537 15552
rect 4304 15512 4310 15524
rect 4525 15521 4537 15524
rect 4571 15521 4583 15555
rect 4525 15515 4583 15521
rect 7193 15555 7251 15561
rect 7193 15521 7205 15555
rect 7239 15552 7251 15555
rect 7558 15552 7564 15564
rect 7239 15524 7564 15552
rect 7239 15521 7251 15524
rect 7193 15515 7251 15521
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 8202 15512 8208 15564
rect 8260 15552 8266 15564
rect 8297 15555 8355 15561
rect 8297 15552 8309 15555
rect 8260 15524 8309 15552
rect 8260 15512 8266 15524
rect 8297 15521 8309 15524
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 8386 15512 8392 15564
rect 8444 15552 8450 15564
rect 8570 15552 8576 15564
rect 8444 15524 8576 15552
rect 8444 15512 8450 15524
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 4614 15484 4620 15496
rect 4575 15456 4620 15484
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15484 6331 15487
rect 6638 15484 6644 15496
rect 6319 15456 6644 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 5350 15376 5356 15428
rect 5408 15416 5414 15428
rect 5537 15419 5595 15425
rect 5537 15416 5549 15419
rect 5408 15388 5549 15416
rect 5408 15376 5414 15388
rect 5537 15385 5549 15388
rect 5583 15416 5595 15419
rect 6288 15416 6316 15447
rect 6638 15444 6644 15456
rect 6696 15484 6702 15496
rect 6822 15484 6828 15496
rect 6696 15456 6828 15484
rect 6696 15444 6702 15456
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 7282 15444 7288 15496
rect 7340 15484 7346 15496
rect 7926 15484 7932 15496
rect 7340 15456 7932 15484
rect 7340 15444 7346 15456
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 8478 15484 8484 15496
rect 8439 15456 8484 15484
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 10042 15444 10048 15496
rect 10100 15484 10106 15496
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10100 15456 10977 15484
rect 10100 15444 10106 15456
rect 10965 15453 10977 15456
rect 11011 15453 11023 15487
rect 11146 15484 11152 15496
rect 11107 15456 11152 15484
rect 10965 15447 11023 15453
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 5583 15388 6316 15416
rect 5583 15385 5595 15388
rect 5537 15379 5595 15385
rect 3237 15351 3295 15357
rect 3237 15317 3249 15351
rect 3283 15348 3295 15351
rect 3510 15348 3516 15360
rect 3283 15320 3516 15348
rect 3283 15317 3295 15320
rect 3237 15311 3295 15317
rect 3510 15308 3516 15320
rect 3568 15308 3574 15360
rect 5626 15348 5632 15360
rect 5587 15320 5632 15348
rect 5626 15308 5632 15320
rect 5684 15308 5690 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 2498 15104 2504 15156
rect 2556 15144 2562 15156
rect 3145 15147 3203 15153
rect 3145 15144 3157 15147
rect 2556 15116 3157 15144
rect 2556 15104 2562 15116
rect 3145 15113 3157 15116
rect 3191 15113 3203 15147
rect 3145 15107 3203 15113
rect 5994 15104 6000 15156
rect 6052 15144 6058 15156
rect 6825 15147 6883 15153
rect 6825 15144 6837 15147
rect 6052 15116 6837 15144
rect 6052 15104 6058 15116
rect 6825 15113 6837 15116
rect 6871 15113 6883 15147
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 6825 15107 6883 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 8662 15144 8668 15156
rect 8623 15116 8668 15144
rect 8662 15104 8668 15116
rect 8720 15104 8726 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 10042 15144 10048 15156
rect 9732 15116 10048 15144
rect 9732 15104 9738 15116
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 10505 15147 10563 15153
rect 10505 15113 10517 15147
rect 10551 15144 10563 15147
rect 10686 15144 10692 15156
rect 10551 15116 10692 15144
rect 10551 15113 10563 15116
rect 10505 15107 10563 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 11146 15104 11152 15156
rect 11204 15144 11210 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11204 15116 11897 15144
rect 11204 15104 11210 15116
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 5902 15036 5908 15088
rect 5960 15076 5966 15088
rect 6181 15079 6239 15085
rect 6181 15076 6193 15079
rect 5960 15048 6193 15076
rect 5960 15036 5966 15048
rect 6181 15045 6193 15048
rect 6227 15045 6239 15079
rect 6181 15039 6239 15045
rect 7929 15079 7987 15085
rect 7929 15045 7941 15079
rect 7975 15076 7987 15079
rect 8202 15076 8208 15088
rect 7975 15048 8208 15076
rect 7975 15045 7987 15048
rect 7929 15039 7987 15045
rect 1578 15008 1584 15020
rect 1539 14980 1584 15008
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 15008 3111 15011
rect 3789 15011 3847 15017
rect 3789 15008 3801 15011
rect 3099 14980 3801 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 3789 14977 3801 14980
rect 3835 15008 3847 15011
rect 4062 15008 4068 15020
rect 3835 14980 4068 15008
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 4798 14968 4804 15020
rect 4856 15008 4862 15020
rect 4985 15011 5043 15017
rect 4985 15008 4997 15011
rect 4856 14980 4997 15008
rect 4856 14968 4862 14980
rect 4985 14977 4997 14980
rect 5031 15008 5043 15011
rect 5718 15008 5724 15020
rect 5031 14980 5580 15008
rect 5679 14980 5724 15008
rect 5031 14977 5043 14980
rect 4985 14971 5043 14977
rect 5552 14949 5580 14980
rect 5718 14968 5724 14980
rect 5776 14968 5782 15020
rect 6196 15008 6224 15039
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 6822 15008 6828 15020
rect 6196 14980 6828 15008
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7282 15008 7288 15020
rect 6972 14980 7288 15008
rect 6972 14968 6978 14980
rect 7282 14968 7288 14980
rect 7340 15008 7346 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 7340 14980 7389 15008
rect 7340 14968 7346 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 9125 15011 9183 15017
rect 9125 15008 9137 15011
rect 8904 14980 9137 15008
rect 8904 14968 8910 14980
rect 9125 14977 9137 14980
rect 9171 14977 9183 15011
rect 9306 15008 9312 15020
rect 9267 14980 9312 15008
rect 9125 14971 9183 14977
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 10962 14968 10968 15020
rect 11020 14968 11026 15020
rect 11164 15017 11192 15104
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 14977 11207 15011
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 11149 14971 11207 14977
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14909 1455 14943
rect 1397 14903 1455 14909
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14909 5595 14943
rect 5537 14903 5595 14909
rect 7193 14943 7251 14949
rect 7193 14909 7205 14943
rect 7239 14940 7251 14943
rect 7466 14940 7472 14952
rect 7239 14912 7472 14940
rect 7239 14909 7251 14912
rect 7193 14903 7251 14909
rect 1412 14872 1440 14903
rect 7466 14900 7472 14912
rect 7524 14900 7530 14952
rect 8662 14900 8668 14952
rect 8720 14940 8726 14952
rect 9398 14940 9404 14952
rect 8720 14912 9404 14940
rect 8720 14900 8726 14912
rect 9398 14900 9404 14912
rect 9456 14900 9462 14952
rect 10318 14900 10324 14952
rect 10376 14940 10382 14952
rect 10980 14940 11008 14968
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 10376 14912 11529 14940
rect 10376 14900 10382 14912
rect 11517 14909 11529 14912
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 13265 14943 13323 14949
rect 13265 14909 13277 14943
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 2222 14872 2228 14884
rect 1412 14844 2228 14872
rect 2222 14832 2228 14844
rect 2280 14832 2286 14884
rect 5902 14832 5908 14884
rect 5960 14872 5966 14884
rect 6641 14875 6699 14881
rect 6641 14872 6653 14875
rect 5960 14844 6653 14872
rect 5960 14832 5966 14844
rect 6641 14841 6653 14844
rect 6687 14872 6699 14875
rect 7285 14875 7343 14881
rect 7285 14872 7297 14875
rect 6687 14844 7297 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7285 14841 7297 14844
rect 7331 14872 7343 14875
rect 7558 14872 7564 14884
rect 7331 14844 7564 14872
rect 7331 14841 7343 14844
rect 7285 14835 7343 14841
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 10965 14875 11023 14881
rect 10965 14872 10977 14875
rect 10336 14844 10977 14872
rect 3510 14804 3516 14816
rect 3471 14776 3516 14804
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 3602 14764 3608 14816
rect 3660 14804 3666 14816
rect 4246 14804 4252 14816
rect 3660 14776 3705 14804
rect 4207 14776 4252 14804
rect 3660 14764 3666 14776
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4617 14807 4675 14813
rect 4617 14773 4629 14807
rect 4663 14804 4675 14807
rect 4706 14804 4712 14816
rect 4663 14776 4712 14804
rect 4663 14773 4675 14776
rect 4617 14767 4675 14773
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 5166 14804 5172 14816
rect 5127 14776 5172 14804
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 5994 14804 6000 14816
rect 5684 14776 6000 14804
rect 5684 14764 5690 14776
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 9033 14807 9091 14813
rect 9033 14804 9045 14807
rect 8904 14776 9045 14804
rect 8904 14764 8910 14776
rect 9033 14773 9045 14776
rect 9079 14773 9091 14807
rect 9033 14767 9091 14773
rect 10226 14764 10232 14816
rect 10284 14804 10290 14816
rect 10336 14813 10364 14844
rect 10965 14841 10977 14844
rect 11011 14841 11023 14875
rect 10965 14835 11023 14841
rect 11238 14832 11244 14884
rect 11296 14872 11302 14884
rect 13280 14872 13308 14903
rect 14001 14875 14059 14881
rect 14001 14872 14013 14875
rect 11296 14844 14013 14872
rect 11296 14832 11302 14844
rect 14001 14841 14013 14844
rect 14047 14841 14059 14875
rect 14001 14835 14059 14841
rect 10321 14807 10379 14813
rect 10321 14804 10333 14807
rect 10284 14776 10333 14804
rect 10284 14764 10290 14776
rect 10321 14773 10333 14776
rect 10367 14773 10379 14807
rect 10321 14767 10379 14773
rect 10778 14764 10784 14816
rect 10836 14804 10842 14816
rect 10873 14807 10931 14813
rect 10873 14804 10885 14807
rect 10836 14776 10885 14804
rect 10836 14764 10842 14776
rect 10873 14773 10885 14776
rect 10919 14773 10931 14807
rect 10873 14767 10931 14773
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 3602 14600 3608 14612
rect 3283 14572 3608 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 3602 14560 3608 14572
rect 3660 14600 3666 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 3660 14572 4077 14600
rect 3660 14560 3666 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 5166 14560 5172 14612
rect 5224 14600 5230 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5224 14572 6009 14600
rect 5224 14560 5230 14572
rect 5997 14569 6009 14572
rect 6043 14600 6055 14603
rect 7006 14600 7012 14612
rect 6043 14572 7012 14600
rect 6043 14569 6055 14572
rect 5997 14563 6055 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7282 14600 7288 14612
rect 7243 14572 7288 14600
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 7524 14572 8493 14600
rect 7524 14560 7530 14572
rect 8481 14569 8493 14572
rect 8527 14600 8539 14603
rect 8754 14600 8760 14612
rect 8527 14572 8760 14600
rect 8527 14569 8539 14572
rect 8481 14563 8539 14569
rect 8754 14560 8760 14572
rect 8812 14560 8818 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 8904 14572 9689 14600
rect 8904 14560 8910 14572
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 9677 14563 9735 14569
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10045 14603 10103 14609
rect 10045 14600 10057 14603
rect 9916 14572 10057 14600
rect 9916 14560 9922 14572
rect 10045 14569 10057 14572
rect 10091 14600 10103 14603
rect 10962 14600 10968 14612
rect 10091 14572 10968 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11146 14600 11152 14612
rect 11107 14572 11152 14600
rect 11146 14560 11152 14572
rect 11204 14600 11210 14612
rect 12897 14603 12955 14609
rect 12897 14600 12909 14603
rect 11204 14572 12909 14600
rect 11204 14560 11210 14572
rect 12897 14569 12909 14572
rect 12943 14569 12955 14603
rect 12897 14563 12955 14569
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 6089 14535 6147 14541
rect 6089 14532 6101 14535
rect 5592 14504 6101 14532
rect 5592 14492 5598 14504
rect 6089 14501 6101 14504
rect 6135 14532 6147 14535
rect 6362 14532 6368 14544
rect 6135 14504 6368 14532
rect 6135 14501 6147 14504
rect 6089 14495 6147 14501
rect 6362 14492 6368 14504
rect 6420 14492 6426 14544
rect 6917 14535 6975 14541
rect 6917 14501 6929 14535
rect 6963 14532 6975 14535
rect 7484 14532 7512 14560
rect 6963 14504 7512 14532
rect 6963 14501 6975 14504
rect 6917 14495 6975 14501
rect 9582 14492 9588 14544
rect 9640 14532 9646 14544
rect 9950 14532 9956 14544
rect 9640 14504 9956 14532
rect 9640 14492 9646 14504
rect 9950 14492 9956 14504
rect 10008 14532 10014 14544
rect 10008 14504 10272 14532
rect 10008 14492 10014 14504
rect 4430 14464 4436 14476
rect 4391 14436 4436 14464
rect 4430 14424 4436 14436
rect 4488 14424 4494 14476
rect 4522 14424 4528 14476
rect 4580 14464 4586 14476
rect 5166 14464 5172 14476
rect 4580 14436 4625 14464
rect 5079 14436 5172 14464
rect 4580 14424 4586 14436
rect 5166 14424 5172 14436
rect 5224 14464 5230 14476
rect 5718 14464 5724 14476
rect 5224 14436 5724 14464
rect 5224 14424 5230 14436
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14464 7987 14467
rect 8478 14464 8484 14476
rect 7975 14436 8484 14464
rect 7975 14433 7987 14436
rect 7929 14427 7987 14433
rect 8478 14424 8484 14436
rect 8536 14464 8542 14476
rect 8849 14467 8907 14473
rect 8849 14464 8861 14467
rect 8536 14436 8861 14464
rect 8536 14424 8542 14436
rect 8849 14433 8861 14436
rect 8895 14433 8907 14467
rect 8849 14427 8907 14433
rect 4614 14396 4620 14408
rect 4575 14368 4620 14396
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 5537 14399 5595 14405
rect 5537 14365 5549 14399
rect 5583 14396 5595 14399
rect 5810 14396 5816 14408
rect 5583 14368 5816 14396
rect 5583 14365 5595 14368
rect 5537 14359 5595 14365
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 6178 14396 6184 14408
rect 6139 14368 6184 14396
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 9674 14396 9680 14408
rect 6788 14368 9680 14396
rect 6788 14356 6794 14368
rect 9674 14356 9680 14368
rect 9732 14396 9738 14408
rect 10244 14405 10272 14504
rect 11514 14464 11520 14476
rect 11475 14436 11520 14464
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 11790 14473 11796 14476
rect 11784 14464 11796 14473
rect 11751 14436 11796 14464
rect 11784 14427 11796 14436
rect 11790 14424 11796 14427
rect 11848 14424 11854 14476
rect 10137 14399 10195 14405
rect 10137 14396 10149 14399
rect 9732 14368 10149 14396
rect 9732 14356 9738 14368
rect 10137 14365 10149 14368
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 2409 14331 2467 14337
rect 2409 14297 2421 14331
rect 2455 14328 2467 14331
rect 3881 14331 3939 14337
rect 3881 14328 3893 14331
rect 2455 14300 3893 14328
rect 2455 14297 2467 14300
rect 2409 14291 2467 14297
rect 3881 14297 3893 14300
rect 3927 14328 3939 14331
rect 4154 14328 4160 14340
rect 3927 14300 4160 14328
rect 3927 14297 3939 14300
rect 3881 14291 3939 14297
rect 4154 14288 4160 14300
rect 4212 14328 4218 14340
rect 4632 14328 4660 14356
rect 4212 14300 4660 14328
rect 4212 14288 4218 14300
rect 5626 14260 5632 14272
rect 5587 14232 5632 14260
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 9490 14260 9496 14272
rect 9451 14232 9496 14260
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 10134 14220 10140 14272
rect 10192 14260 10198 14272
rect 10689 14263 10747 14269
rect 10689 14260 10701 14263
rect 10192 14232 10701 14260
rect 10192 14220 10198 14232
rect 10689 14229 10701 14232
rect 10735 14260 10747 14263
rect 10778 14260 10784 14272
rect 10735 14232 10784 14260
rect 10735 14229 10747 14232
rect 10689 14223 10747 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 2317 14059 2375 14065
rect 2317 14025 2329 14059
rect 2363 14056 2375 14059
rect 3510 14056 3516 14068
rect 2363 14028 3516 14056
rect 2363 14025 2375 14028
rect 2317 14019 2375 14025
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 4062 14016 4068 14068
rect 4120 14056 4126 14068
rect 5261 14059 5319 14065
rect 5261 14056 5273 14059
rect 4120 14028 5273 14056
rect 4120 14016 4126 14028
rect 5261 14025 5273 14028
rect 5307 14025 5319 14059
rect 5994 14056 6000 14068
rect 5955 14028 6000 14056
rect 5261 14019 5319 14025
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 6362 14056 6368 14068
rect 6323 14028 6368 14056
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 7006 14056 7012 14068
rect 6967 14028 7012 14056
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7558 14016 7564 14068
rect 7616 14056 7622 14068
rect 8297 14059 8355 14065
rect 8297 14056 8309 14059
rect 7616 14028 8309 14056
rect 7616 14016 7622 14028
rect 8297 14025 8309 14028
rect 8343 14025 8355 14059
rect 9674 14056 9680 14068
rect 9635 14028 9680 14056
rect 8297 14019 8355 14025
rect 8312 13988 8340 14019
rect 9674 14016 9680 14028
rect 9732 14056 9738 14068
rect 9858 14056 9864 14068
rect 9732 14028 9864 14056
rect 9732 14016 9738 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 11020 14028 11069 14056
rect 11020 14016 11026 14028
rect 11057 14025 11069 14028
rect 11103 14025 11115 14059
rect 11057 14019 11115 14025
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11572 14028 12173 14056
rect 11572 14016 11578 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 8938 13988 8944 14000
rect 8312 13960 8944 13988
rect 8938 13948 8944 13960
rect 8996 13948 9002 14000
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13920 3019 13923
rect 3421 13923 3479 13929
rect 3421 13920 3433 13923
rect 3007 13892 3433 13920
rect 3007 13889 3019 13892
rect 2961 13883 3019 13889
rect 3421 13889 3433 13892
rect 3467 13920 3479 13923
rect 8021 13923 8079 13929
rect 3467 13892 4016 13920
rect 3467 13889 3479 13892
rect 3421 13883 3479 13889
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13852 2743 13855
rect 2774 13852 2780 13864
rect 2731 13824 2780 13852
rect 2731 13821 2743 13824
rect 2685 13815 2743 13821
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 3878 13852 3884 13864
rect 3839 13824 3884 13852
rect 3878 13812 3884 13824
rect 3936 13812 3942 13864
rect 3988 13852 4016 13892
rect 8021 13889 8033 13923
rect 8067 13920 8079 13923
rect 9125 13923 9183 13929
rect 9125 13920 9137 13923
rect 8067 13892 9137 13920
rect 8067 13889 8079 13892
rect 8021 13883 8079 13889
rect 9125 13889 9137 13892
rect 9171 13889 9183 13923
rect 9125 13883 9183 13889
rect 4154 13861 4160 13864
rect 4148 13852 4160 13861
rect 3988 13824 4160 13852
rect 4148 13815 4160 13824
rect 4154 13812 4160 13815
rect 4212 13812 4218 13864
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 8754 13852 8760 13864
rect 8444 13824 8760 13852
rect 8444 13812 8450 13824
rect 8754 13812 8760 13824
rect 8812 13852 8818 13864
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8812 13824 8861 13852
rect 8812 13812 8818 13824
rect 8849 13821 8861 13824
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 8938 13812 8944 13864
rect 8996 13852 9002 13864
rect 9140 13852 9168 13883
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 10042 13920 10048 13932
rect 9548 13892 10048 13920
rect 9548 13880 9554 13892
rect 10042 13880 10048 13892
rect 10100 13920 10106 13932
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 10100 13892 10517 13920
rect 10100 13880 10106 13892
rect 10505 13889 10517 13892
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 9674 13852 9680 13864
rect 8996 13824 9041 13852
rect 9140 13824 9680 13852
rect 8996 13812 9002 13824
rect 9674 13812 9680 13824
rect 9732 13812 9738 13864
rect 10704 13852 10732 13883
rect 11517 13855 11575 13861
rect 11517 13852 11529 13855
rect 10704 13824 11529 13852
rect 11517 13821 11529 13824
rect 11563 13852 11575 13855
rect 11790 13852 11796 13864
rect 11563 13824 11796 13852
rect 11563 13821 11575 13824
rect 11517 13815 11575 13821
rect 11790 13812 11796 13824
rect 11848 13852 11854 13864
rect 11885 13855 11943 13861
rect 11885 13852 11897 13855
rect 11848 13824 11897 13852
rect 11848 13812 11854 13824
rect 11885 13821 11897 13824
rect 11931 13852 11943 13855
rect 12342 13852 12348 13864
rect 11931 13824 12348 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 2225 13787 2283 13793
rect 2225 13753 2237 13787
rect 2271 13784 2283 13787
rect 3789 13787 3847 13793
rect 2271 13756 2820 13784
rect 2271 13753 2283 13756
rect 2225 13747 2283 13753
rect 2792 13725 2820 13756
rect 3789 13753 3801 13787
rect 3835 13784 3847 13787
rect 4522 13784 4528 13796
rect 3835 13756 4528 13784
rect 3835 13753 3847 13756
rect 3789 13747 3847 13753
rect 4522 13744 4528 13756
rect 4580 13744 4586 13796
rect 7190 13784 7196 13796
rect 5644 13756 7196 13784
rect 2777 13719 2835 13725
rect 2777 13685 2789 13719
rect 2823 13716 2835 13719
rect 5644 13716 5672 13756
rect 7190 13744 7196 13756
rect 7248 13744 7254 13796
rect 2823 13688 5672 13716
rect 5721 13719 5779 13725
rect 2823 13685 2835 13688
rect 2777 13679 2835 13685
rect 5721 13685 5733 13719
rect 5767 13716 5779 13719
rect 5810 13716 5816 13728
rect 5767 13688 5816 13716
rect 5767 13685 5779 13688
rect 5721 13679 5779 13685
rect 5810 13676 5816 13688
rect 5868 13716 5874 13728
rect 6178 13716 6184 13728
rect 5868 13688 6184 13716
rect 5868 13676 5874 13688
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 8478 13716 8484 13728
rect 8439 13688 8484 13716
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 10410 13716 10416 13728
rect 10371 13688 10416 13716
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 2774 13512 2780 13524
rect 2455 13484 2780 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4617 13515 4675 13521
rect 4617 13512 4629 13515
rect 4212 13484 4629 13512
rect 4212 13472 4218 13484
rect 4617 13481 4629 13484
rect 4663 13481 4675 13515
rect 8846 13512 8852 13524
rect 8807 13484 8852 13512
rect 4617 13475 4675 13481
rect 8846 13472 8852 13484
rect 8904 13472 8910 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 9582 13512 9588 13524
rect 9539 13484 9588 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 1670 13444 1676 13456
rect 1631 13416 1676 13444
rect 1670 13404 1676 13416
rect 1728 13404 1734 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2792 13376 2820 13472
rect 4341 13447 4399 13453
rect 4341 13413 4353 13447
rect 4387 13444 4399 13447
rect 4430 13444 4436 13456
rect 4387 13416 4436 13444
rect 4387 13413 4399 13416
rect 4341 13407 4399 13413
rect 4430 13404 4436 13416
rect 4488 13404 4494 13456
rect 5166 13453 5172 13456
rect 5160 13444 5172 13453
rect 5127 13416 5172 13444
rect 5160 13407 5172 13416
rect 5166 13404 5172 13407
rect 5224 13404 5230 13456
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 8754 13444 8760 13456
rect 8352 13416 8760 13444
rect 8352 13404 8358 13416
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 9674 13404 9680 13456
rect 9732 13444 9738 13456
rect 9922 13447 9980 13453
rect 9922 13444 9934 13447
rect 9732 13416 9934 13444
rect 9732 13404 9738 13416
rect 9922 13413 9934 13416
rect 9968 13413 9980 13447
rect 9922 13407 9980 13413
rect 6730 13376 6736 13388
rect 1443 13348 1716 13376
rect 2792 13348 6736 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1688 13320 1716 13348
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 7098 13376 7104 13388
rect 7059 13348 7104 13376
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 7368 13379 7426 13385
rect 7368 13345 7380 13379
rect 7414 13376 7426 13379
rect 8202 13376 8208 13388
rect 7414 13348 8208 13376
rect 7414 13345 7426 13348
rect 7368 13339 7426 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 1670 13268 1676 13320
rect 1728 13268 1734 13320
rect 4614 13308 4620 13320
rect 3896 13280 4620 13308
rect 3896 13252 3924 13280
rect 4614 13268 4620 13280
rect 4672 13308 4678 13320
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4672 13280 4905 13308
rect 4672 13268 4678 13280
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9640 13280 9689 13308
rect 9640 13268 9646 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 3878 13200 3884 13252
rect 3936 13200 3942 13252
rect 6730 13200 6736 13252
rect 6788 13240 6794 13252
rect 6917 13243 6975 13249
rect 6917 13240 6929 13243
rect 6788 13212 6929 13240
rect 6788 13200 6794 13212
rect 6917 13209 6929 13212
rect 6963 13209 6975 13243
rect 6917 13203 6975 13209
rect 2498 13132 2504 13184
rect 2556 13172 2562 13184
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 2556 13144 3801 13172
rect 2556 13132 2562 13144
rect 3789 13141 3801 13144
rect 3835 13172 3847 13175
rect 3896 13172 3924 13200
rect 3835 13144 3924 13172
rect 3835 13141 3847 13144
rect 3789 13135 3847 13141
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 6086 13172 6092 13184
rect 5868 13144 6092 13172
rect 5868 13132 5874 13144
rect 6086 13132 6092 13144
rect 6144 13172 6150 13184
rect 6273 13175 6331 13181
rect 6273 13172 6285 13175
rect 6144 13144 6285 13172
rect 6144 13132 6150 13144
rect 6273 13141 6285 13144
rect 6319 13141 6331 13175
rect 6273 13135 6331 13141
rect 6641 13175 6699 13181
rect 6641 13141 6653 13175
rect 6687 13172 6699 13175
rect 6822 13172 6828 13184
rect 6687 13144 6828 13172
rect 6687 13141 6699 13144
rect 6641 13135 6699 13141
rect 6822 13132 6828 13144
rect 6880 13132 6886 13184
rect 8481 13175 8539 13181
rect 8481 13141 8493 13175
rect 8527 13172 8539 13175
rect 8846 13172 8852 13184
rect 8527 13144 8852 13172
rect 8527 13141 8539 13144
rect 8481 13135 8539 13141
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 9950 13172 9956 13184
rect 9456 13144 9956 13172
rect 9456 13132 9462 13144
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10836 13144 11069 13172
rect 10836 13132 10842 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 3881 12971 3939 12977
rect 3881 12937 3893 12971
rect 3927 12968 3939 12971
rect 4154 12968 4160 12980
rect 3927 12940 4160 12968
rect 3927 12937 3939 12940
rect 3881 12931 3939 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4985 12971 5043 12977
rect 4985 12937 4997 12971
rect 5031 12968 5043 12971
rect 5166 12968 5172 12980
rect 5031 12940 5172 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 7098 12968 7104 12980
rect 5951 12940 7104 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 5261 12903 5319 12909
rect 5261 12900 5273 12903
rect 4672 12872 5273 12900
rect 4672 12860 4678 12872
rect 5261 12869 5273 12872
rect 5307 12869 5319 12903
rect 5261 12863 5319 12869
rect 2498 12764 2504 12776
rect 2459 12736 2504 12764
rect 2498 12724 2504 12736
rect 2556 12724 2562 12776
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3970 12764 3976 12776
rect 3200 12736 3976 12764
rect 3200 12724 3206 12736
rect 3970 12724 3976 12736
rect 4028 12724 4034 12776
rect 5276 12764 5304 12863
rect 6840 12832 6868 12940
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 8202 12968 8208 12980
rect 7616 12940 8208 12968
rect 7616 12928 7622 12940
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 8478 12968 8484 12980
rect 8439 12940 8484 12968
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 10042 12928 10048 12980
rect 10100 12928 10106 12980
rect 10410 12928 10416 12980
rect 10468 12968 10474 12980
rect 10689 12971 10747 12977
rect 10689 12968 10701 12971
rect 10468 12940 10701 12968
rect 10468 12928 10474 12940
rect 10689 12937 10701 12940
rect 10735 12937 10747 12971
rect 10689 12931 10747 12937
rect 11149 12971 11207 12977
rect 11149 12937 11161 12971
rect 11195 12968 11207 12971
rect 11514 12968 11520 12980
rect 11195 12940 11520 12968
rect 11195 12937 11207 12940
rect 11149 12931 11207 12937
rect 6840 12804 6960 12832
rect 6730 12764 6736 12776
rect 5276 12736 6736 12764
rect 6730 12724 6736 12736
rect 6788 12764 6794 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6788 12736 6837 12764
rect 6788 12724 6794 12736
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 6932 12764 6960 12804
rect 10060 12776 10088 12928
rect 10502 12860 10508 12912
rect 10560 12900 10566 12912
rect 11164 12900 11192 12931
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 10560 12872 11192 12900
rect 10560 12860 10566 12872
rect 9030 12764 9036 12776
rect 6932 12736 9036 12764
rect 6825 12727 6883 12733
rect 9030 12724 9036 12736
rect 9088 12764 9094 12776
rect 9582 12764 9588 12776
rect 9088 12736 9588 12764
rect 9088 12724 9094 12736
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 10042 12724 10048 12776
rect 10100 12724 10106 12776
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 2682 12696 2688 12708
rect 2455 12668 2688 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 2682 12656 2688 12668
rect 2740 12705 2746 12708
rect 2740 12699 2804 12705
rect 2740 12665 2758 12699
rect 2792 12665 2804 12699
rect 2740 12659 2804 12665
rect 6273 12699 6331 12705
rect 6273 12665 6285 12699
rect 6319 12696 6331 12699
rect 6638 12696 6644 12708
rect 6319 12668 6644 12696
rect 6319 12665 6331 12668
rect 6273 12659 6331 12665
rect 2740 12656 2746 12659
rect 6638 12656 6644 12668
rect 6696 12656 6702 12708
rect 7092 12699 7150 12705
rect 7092 12696 7104 12699
rect 7024 12668 7104 12696
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12628 6607 12631
rect 7024 12628 7052 12668
rect 7092 12665 7104 12668
rect 7138 12696 7150 12699
rect 7834 12696 7840 12708
rect 7138 12668 7840 12696
rect 7138 12665 7150 12668
rect 7092 12659 7150 12665
rect 7834 12656 7840 12668
rect 7892 12656 7898 12708
rect 9278 12699 9336 12705
rect 9278 12696 9290 12699
rect 8864 12668 9290 12696
rect 8864 12640 8892 12668
rect 9278 12665 9290 12668
rect 9324 12665 9336 12699
rect 9278 12659 9336 12665
rect 8846 12628 8852 12640
rect 6595 12600 7052 12628
rect 8807 12600 8852 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10134 12628 10140 12640
rect 9732 12600 10140 12628
rect 9732 12588 9738 12600
rect 10134 12588 10140 12600
rect 10192 12628 10198 12640
rect 10413 12631 10471 12637
rect 10413 12628 10425 12631
rect 10192 12600 10425 12628
rect 10192 12588 10198 12600
rect 10413 12597 10425 12600
rect 10459 12597 10471 12631
rect 10413 12591 10471 12597
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 4614 12384 4620 12436
rect 4672 12424 4678 12436
rect 4893 12427 4951 12433
rect 4893 12424 4905 12427
rect 4672 12396 4905 12424
rect 4672 12384 4678 12396
rect 4893 12393 4905 12396
rect 4939 12393 4951 12427
rect 4893 12387 4951 12393
rect 5074 12384 5080 12436
rect 5132 12384 5138 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 6457 12427 6515 12433
rect 6457 12424 6469 12427
rect 5592 12396 6469 12424
rect 5592 12384 5598 12396
rect 6457 12393 6469 12396
rect 6503 12393 6515 12427
rect 8478 12424 8484 12436
rect 8439 12396 8484 12424
rect 6457 12387 6515 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 10134 12424 10140 12436
rect 10095 12396 10140 12424
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12492 12396 12537 12424
rect 12492 12384 12498 12396
rect 4982 12316 4988 12368
rect 5040 12356 5046 12368
rect 5092 12356 5120 12384
rect 5040 12328 5120 12356
rect 5040 12316 5046 12328
rect 6546 12316 6552 12368
rect 6604 12356 6610 12368
rect 6914 12356 6920 12368
rect 6604 12328 6920 12356
rect 6604 12316 6610 12328
rect 6914 12316 6920 12328
rect 6972 12316 6978 12368
rect 5074 12288 5080 12300
rect 5035 12260 5080 12288
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 6822 12288 6828 12300
rect 6783 12260 6828 12288
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 8260 12260 8401 12288
rect 8260 12248 8266 12260
rect 8389 12257 8401 12260
rect 8435 12288 8447 12291
rect 9858 12288 9864 12300
rect 8435 12260 9864 12288
rect 8435 12257 8447 12260
rect 8389 12251 8447 12257
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 10870 12288 10876 12300
rect 10831 12260 10876 12288
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11313 12291 11371 12297
rect 11313 12288 11325 12291
rect 11020 12260 11325 12288
rect 11020 12248 11026 12260
rect 11313 12257 11325 12260
rect 11359 12257 11371 12291
rect 11313 12251 11371 12257
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 6914 12220 6920 12232
rect 6696 12192 6920 12220
rect 6696 12180 6702 12192
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12220 7987 12223
rect 8573 12223 8631 12229
rect 8573 12220 8585 12223
rect 7975 12192 8585 12220
rect 7975 12189 7987 12192
rect 7929 12183 7987 12189
rect 8573 12189 8585 12192
rect 8619 12220 8631 12223
rect 8846 12220 8852 12232
rect 8619 12192 8852 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 6730 12112 6736 12164
rect 6788 12152 6794 12164
rect 7024 12152 7052 12183
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 10502 12180 10508 12232
rect 10560 12220 10566 12232
rect 11057 12223 11115 12229
rect 11057 12220 11069 12223
rect 10560 12192 11069 12220
rect 10560 12180 10566 12192
rect 6788 12124 7052 12152
rect 6788 12112 6794 12124
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 9125 12155 9183 12161
rect 9125 12152 9137 12155
rect 9088 12124 9137 12152
rect 9088 12112 9094 12124
rect 9125 12121 9137 12124
rect 9171 12152 9183 12155
rect 10704 12152 10732 12192
rect 11057 12189 11069 12192
rect 11103 12189 11115 12223
rect 11057 12183 11115 12189
rect 9171 12124 10732 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 10704 12096 10732 12124
rect 1762 12044 1768 12096
rect 1820 12084 1826 12096
rect 2498 12084 2504 12096
rect 1820 12056 2504 12084
rect 1820 12044 1826 12056
rect 2498 12044 2504 12056
rect 2556 12044 2562 12096
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5445 12087 5503 12093
rect 5445 12084 5457 12087
rect 5224 12056 5457 12084
rect 5224 12044 5230 12056
rect 5445 12053 5457 12056
rect 5491 12084 5503 12087
rect 5718 12084 5724 12096
rect 5491 12056 5724 12084
rect 5491 12053 5503 12056
rect 5445 12047 5503 12053
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 5994 12084 6000 12096
rect 5955 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6365 12087 6423 12093
rect 6365 12053 6377 12087
rect 6411 12084 6423 12087
rect 7374 12084 7380 12096
rect 6411 12056 7380 12084
rect 6411 12053 6423 12056
rect 6365 12047 6423 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 7558 12084 7564 12096
rect 7519 12056 7564 12084
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 10502 12084 10508 12096
rect 10463 12056 10508 12084
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 4341 11883 4399 11889
rect 4341 11849 4353 11883
rect 4387 11880 4399 11883
rect 5074 11880 5080 11892
rect 4387 11852 5080 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 6549 11883 6607 11889
rect 6549 11849 6561 11883
rect 6595 11880 6607 11883
rect 6730 11880 6736 11892
rect 6595 11852 6736 11880
rect 6595 11849 6607 11852
rect 6549 11843 6607 11849
rect 6730 11840 6736 11852
rect 6788 11840 6794 11892
rect 6822 11840 6828 11892
rect 6880 11880 6886 11892
rect 6917 11883 6975 11889
rect 6917 11880 6929 11883
rect 6880 11852 6929 11880
rect 6880 11840 6886 11852
rect 6917 11849 6929 11852
rect 6963 11849 6975 11883
rect 6917 11843 6975 11849
rect 8021 11883 8079 11889
rect 8021 11849 8033 11883
rect 8067 11880 8079 11883
rect 8202 11880 8208 11892
rect 8067 11852 8208 11880
rect 8067 11849 8079 11852
rect 8021 11843 8079 11849
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 10042 11880 10048 11892
rect 10003 11852 10048 11880
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 11425 11883 11483 11889
rect 11425 11880 11437 11883
rect 10928 11852 11437 11880
rect 10928 11840 10934 11852
rect 11425 11849 11437 11852
rect 11471 11849 11483 11883
rect 11425 11843 11483 11849
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11572 11852 11805 11880
rect 11572 11840 11578 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 4709 11815 4767 11821
rect 4709 11781 4721 11815
rect 4755 11812 4767 11815
rect 5810 11812 5816 11824
rect 4755 11784 5816 11812
rect 4755 11781 4767 11784
rect 4709 11775 4767 11781
rect 5810 11772 5816 11784
rect 5868 11772 5874 11824
rect 8294 11812 8300 11824
rect 7392 11784 8300 11812
rect 7392 11756 7420 11784
rect 8294 11772 8300 11784
rect 8352 11772 8358 11824
rect 8481 11815 8539 11821
rect 8481 11781 8493 11815
rect 8527 11812 8539 11815
rect 8527 11784 10456 11812
rect 8527 11781 8539 11784
rect 8481 11775 8539 11781
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 5718 11744 5724 11756
rect 5679 11716 5724 11744
rect 5718 11704 5724 11716
rect 5776 11704 5782 11756
rect 7374 11744 7380 11756
rect 7335 11716 7380 11744
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 7558 11744 7564 11756
rect 7519 11716 7564 11744
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 8662 11704 8668 11756
rect 8720 11704 8726 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8904 11716 9045 11744
rect 8904 11704 8910 11716
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 5537 11679 5595 11685
rect 5537 11676 5549 11679
rect 1443 11648 2268 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 2240 11552 2268 11648
rect 5000 11648 5549 11676
rect 5000 11552 5028 11648
rect 5537 11645 5549 11648
rect 5583 11645 5595 11679
rect 5537 11639 5595 11645
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 5810 11676 5816 11688
rect 5675 11648 5816 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 5810 11636 5816 11648
rect 5868 11636 5874 11688
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 6052 11648 7297 11676
rect 6052 11636 6058 11648
rect 7285 11645 7297 11648
rect 7331 11676 7343 11679
rect 8018 11676 8024 11688
rect 7331 11648 8024 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 6822 11608 6828 11620
rect 5184 11580 6828 11608
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 4982 11540 4988 11552
rect 4943 11512 4988 11540
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 5184 11549 5212 11580
rect 6822 11568 6828 11580
rect 6880 11568 6886 11620
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11509 5227 11543
rect 5169 11503 5227 11509
rect 8389 11543 8447 11549
rect 8389 11509 8401 11543
rect 8435 11540 8447 11543
rect 8680 11540 8708 11704
rect 10428 11685 10456 11784
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11744 10747 11747
rect 10962 11744 10968 11756
rect 10735 11716 10968 11744
rect 10735 11713 10747 11716
rect 10689 11707 10747 11713
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11676 10471 11679
rect 10502 11676 10508 11688
rect 10459 11648 10508 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 9953 11611 10011 11617
rect 9953 11577 9965 11611
rect 9999 11608 10011 11611
rect 10704 11608 10732 11707
rect 10962 11704 10968 11716
rect 11020 11744 11026 11756
rect 11020 11716 11192 11744
rect 11020 11704 11026 11716
rect 9999 11580 10732 11608
rect 9999 11577 10011 11580
rect 9953 11571 10011 11577
rect 8754 11540 8760 11552
rect 8435 11512 8760 11540
rect 8435 11509 8447 11512
rect 8389 11503 8447 11509
rect 8754 11500 8760 11512
rect 8812 11540 8818 11552
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 8812 11512 8861 11540
rect 8812 11500 8818 11512
rect 8849 11509 8861 11512
rect 8895 11509 8907 11543
rect 8849 11503 8907 11509
rect 8941 11543 8999 11549
rect 8941 11509 8953 11543
rect 8987 11540 8999 11543
rect 9398 11540 9404 11552
rect 8987 11512 9404 11540
rect 8987 11509 8999 11512
rect 8941 11503 8999 11509
rect 9398 11500 9404 11512
rect 9456 11540 9462 11552
rect 9582 11540 9588 11552
rect 9456 11512 9588 11540
rect 9456 11500 9462 11512
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 11164 11549 11192 11716
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10100 11512 10517 11540
rect 10100 11500 10106 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 10505 11503 10563 11509
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11540 11207 11543
rect 11422 11540 11428 11552
rect 11195 11512 11428 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 11422 11500 11428 11512
rect 11480 11500 11486 11552
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 4798 11336 4804 11348
rect 4759 11308 4804 11336
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 5169 11339 5227 11345
rect 5169 11305 5181 11339
rect 5215 11336 5227 11339
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 5215 11308 6377 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 6365 11305 6377 11308
rect 6411 11305 6423 11339
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 6365 11299 6423 11305
rect 4709 11271 4767 11277
rect 4709 11237 4721 11271
rect 4755 11268 4767 11271
rect 5184 11268 5212 11299
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7834 11336 7840 11348
rect 7795 11308 7840 11336
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 8018 11336 8024 11348
rect 7979 11308 8024 11336
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 8478 11336 8484 11348
rect 8439 11308 8484 11336
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 9033 11339 9091 11345
rect 9033 11336 9045 11339
rect 8904 11308 9045 11336
rect 8904 11296 8910 11308
rect 9033 11305 9045 11308
rect 9079 11305 9091 11339
rect 10042 11336 10048 11348
rect 10003 11308 10048 11336
rect 9033 11299 9091 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 10781 11339 10839 11345
rect 10781 11336 10793 11339
rect 10468 11308 10793 11336
rect 10468 11296 10474 11308
rect 10781 11305 10793 11308
rect 10827 11305 10839 11339
rect 10781 11299 10839 11305
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11514 11336 11520 11348
rect 11112 11308 11520 11336
rect 11112 11296 11118 11308
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 4755 11240 5212 11268
rect 5261 11271 5319 11277
rect 4755 11237 4767 11240
rect 4709 11231 4767 11237
rect 5261 11237 5273 11271
rect 5307 11268 5319 11271
rect 5442 11268 5448 11280
rect 5307 11240 5448 11268
rect 5307 11237 5319 11240
rect 5261 11231 5319 11237
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1670 11200 1676 11212
rect 1443 11172 1676 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1670 11160 1676 11172
rect 1728 11200 1734 11212
rect 2406 11200 2412 11212
rect 1728 11172 2412 11200
rect 1728 11160 1734 11172
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 4062 11160 4068 11212
rect 4120 11200 4126 11212
rect 5276 11200 5304 11231
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 5905 11271 5963 11277
rect 5905 11237 5917 11271
rect 5951 11268 5963 11271
rect 7006 11268 7012 11280
rect 5951 11240 7012 11268
rect 5951 11237 5963 11240
rect 5905 11231 5963 11237
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 4120 11172 5304 11200
rect 6196 11172 6745 11200
rect 4120 11160 4126 11172
rect 1578 11132 1584 11144
rect 1539 11104 1584 11132
rect 1578 11092 1584 11104
rect 1636 11092 1642 11144
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 5353 11135 5411 11141
rect 5353 11132 5365 11135
rect 4764 11104 5365 11132
rect 4764 11092 4770 11104
rect 5353 11101 5365 11104
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 6196 11073 6224 11172
rect 6733 11169 6745 11172
rect 6779 11169 6791 11203
rect 7852 11200 7880 11296
rect 8389 11271 8447 11277
rect 8389 11237 8401 11271
rect 8435 11268 8447 11271
rect 9674 11268 9680 11280
rect 8435 11240 9680 11268
rect 8435 11237 8447 11240
rect 8389 11231 8447 11237
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 10689 11271 10747 11277
rect 10689 11237 10701 11271
rect 10735 11268 10747 11271
rect 11422 11268 11428 11280
rect 10735 11240 11428 11268
rect 10735 11237 10747 11240
rect 10689 11231 10747 11237
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 7852 11172 8616 11200
rect 6733 11163 6791 11169
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 8588 11141 8616 11172
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 11149 11203 11207 11209
rect 11149 11200 11161 11203
rect 11112 11172 11161 11200
rect 11112 11160 11118 11172
rect 11149 11169 11161 11172
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 11974 11160 11980 11212
rect 12032 11200 12038 11212
rect 12250 11200 12256 11212
rect 12032 11172 12256 11200
rect 12032 11160 12038 11172
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6696 11104 6929 11132
rect 6696 11092 6702 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11101 8631 11135
rect 11241 11135 11299 11141
rect 11241 11132 11253 11135
rect 8573 11095 8631 11101
rect 11164 11104 11253 11132
rect 6181 11067 6239 11073
rect 6181 11064 6193 11067
rect 5592 11036 6193 11064
rect 5592 11024 5598 11036
rect 6181 11033 6193 11036
rect 6227 11033 6239 11067
rect 6181 11027 6239 11033
rect 2225 10999 2283 11005
rect 2225 10965 2237 10999
rect 2271 10996 2283 10999
rect 2406 10996 2412 11008
rect 2271 10968 2412 10996
rect 2271 10965 2283 10968
rect 2225 10959 2283 10965
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 7469 10999 7527 11005
rect 7469 10965 7481 10999
rect 7515 10996 7527 10999
rect 7558 10996 7564 11008
rect 7515 10968 7564 10996
rect 7515 10965 7527 10968
rect 7469 10959 7527 10965
rect 7558 10956 7564 10968
rect 7616 10956 7622 11008
rect 8588 10996 8616 11095
rect 11164 11076 11192 11104
rect 11241 11101 11253 11104
rect 11287 11101 11299 11135
rect 11422 11132 11428 11144
rect 11383 11104 11428 11132
rect 11241 11095 11299 11101
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 12342 11132 12348 11144
rect 12303 11104 12348 11132
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 11146 11024 11152 11076
rect 11204 11024 11210 11076
rect 8846 10996 8852 11008
rect 8588 10968 8852 10996
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 11330 10996 11336 11008
rect 10836 10968 11336 10996
rect 10836 10956 10842 10968
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4062 10792 4068 10804
rect 4019 10764 4068 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4706 10792 4712 10804
rect 4667 10764 4712 10792
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5534 10792 5540 10804
rect 5215 10764 5540 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 6972 10764 7021 10792
rect 6972 10752 6978 10764
rect 7009 10761 7021 10764
rect 7055 10761 7067 10795
rect 7009 10755 7067 10761
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 8573 10795 8631 10801
rect 8573 10792 8585 10795
rect 8352 10764 8585 10792
rect 8352 10752 8358 10764
rect 8573 10761 8585 10764
rect 8619 10761 8631 10795
rect 9674 10792 9680 10804
rect 9635 10764 9680 10792
rect 8573 10755 8631 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 10594 10792 10600 10804
rect 10555 10764 10600 10792
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 10781 10795 10839 10801
rect 10781 10761 10793 10795
rect 10827 10792 10839 10795
rect 10962 10792 10968 10804
rect 10827 10764 10968 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 12437 10795 12495 10801
rect 12437 10792 12449 10795
rect 11204 10764 12449 10792
rect 11204 10752 11210 10764
rect 12437 10761 12449 10764
rect 12483 10761 12495 10795
rect 12437 10755 12495 10761
rect 8113 10727 8171 10733
rect 8113 10693 8125 10727
rect 8159 10724 8171 10727
rect 8478 10724 8484 10736
rect 8159 10696 8484 10724
rect 8159 10693 8171 10696
rect 8113 10687 8171 10693
rect 8478 10684 8484 10696
rect 8536 10684 8542 10736
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2682 10656 2688 10668
rect 2087 10628 2688 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 5718 10656 5724 10668
rect 4387 10628 5724 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 7064 10628 7481 10656
rect 7064 10616 7070 10628
rect 7469 10625 7481 10628
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7616 10628 7661 10656
rect 7616 10616 7622 10628
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8904 10628 9137 10656
rect 8904 10616 8910 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 10612 10656 10640 10752
rect 11514 10724 11520 10736
rect 11256 10696 11520 10724
rect 11256 10665 11284 10696
rect 11514 10684 11520 10696
rect 11572 10684 11578 10736
rect 12253 10727 12311 10733
rect 12253 10693 12265 10727
rect 12299 10724 12311 10727
rect 12618 10724 12624 10736
rect 12299 10696 12624 10724
rect 12299 10693 12311 10696
rect 12253 10687 12311 10693
rect 12618 10684 12624 10696
rect 12676 10724 12682 10736
rect 12676 10696 12848 10724
rect 12676 10684 12682 10696
rect 11241 10659 11299 10665
rect 11241 10656 11253 10659
rect 10612 10628 11253 10656
rect 9125 10619 9183 10625
rect 11241 10625 11253 10628
rect 11287 10625 11299 10659
rect 11241 10619 11299 10625
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11388 10628 11805 10656
rect 11388 10616 11394 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10588 5135 10591
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5123 10560 5641 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 5629 10557 5641 10560
rect 5675 10588 5687 10591
rect 6178 10588 6184 10600
rect 5675 10560 6184 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 9030 10588 9036 10600
rect 8943 10560 9036 10588
rect 9030 10548 9036 10560
rect 9088 10588 9094 10600
rect 9398 10588 9404 10600
rect 9088 10560 9404 10588
rect 9088 10548 9094 10560
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10588 10379 10591
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 10367 10560 11161 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 11149 10557 11161 10560
rect 11195 10588 11207 10591
rect 12342 10588 12348 10600
rect 11195 10560 12348 10588
rect 11195 10557 11207 10560
rect 11149 10551 11207 10557
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 12820 10597 12848 10696
rect 12986 10656 12992 10668
rect 12947 10628 12992 10656
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10588 12863 10591
rect 15746 10588 15752 10600
rect 12851 10560 15752 10588
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 1673 10523 1731 10529
rect 1673 10489 1685 10523
rect 1719 10520 1731 10523
rect 1719 10492 2360 10520
rect 1719 10489 1731 10492
rect 1673 10483 1731 10489
rect 2130 10452 2136 10464
rect 2091 10424 2136 10452
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 2332 10452 2360 10492
rect 2406 10480 2412 10532
rect 2464 10520 2470 10532
rect 2593 10523 2651 10529
rect 2593 10520 2605 10523
rect 2464 10492 2605 10520
rect 2464 10480 2470 10492
rect 2593 10489 2605 10492
rect 2639 10489 2651 10523
rect 2593 10483 2651 10489
rect 11330 10480 11336 10532
rect 11388 10520 11394 10532
rect 11606 10520 11612 10532
rect 11388 10492 11612 10520
rect 11388 10480 11394 10492
rect 11606 10480 11612 10492
rect 11664 10480 11670 10532
rect 12434 10480 12440 10532
rect 12492 10520 12498 10532
rect 12894 10520 12900 10532
rect 12492 10492 12900 10520
rect 12492 10480 12498 10492
rect 12894 10480 12900 10492
rect 12952 10480 12958 10532
rect 2501 10455 2559 10461
rect 2501 10452 2513 10455
rect 2332 10424 2513 10452
rect 2501 10421 2513 10424
rect 2547 10452 2559 10455
rect 3418 10452 3424 10464
rect 2547 10424 3424 10452
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 5534 10452 5540 10464
rect 5495 10424 5540 10452
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6086 10412 6092 10464
rect 6144 10452 6150 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 6144 10424 6377 10452
rect 6144 10412 6150 10424
rect 6365 10421 6377 10424
rect 6411 10452 6423 10455
rect 6638 10452 6644 10464
rect 6411 10424 6644 10452
rect 6411 10421 6423 10424
rect 6365 10415 6423 10421
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7374 10452 7380 10464
rect 7335 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10452 8539 10455
rect 8938 10452 8944 10464
rect 8527 10424 8944 10452
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 1670 10248 1676 10260
rect 1631 10220 1676 10248
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 3145 10251 3203 10257
rect 3145 10248 3157 10251
rect 2740 10220 3157 10248
rect 2740 10208 2746 10220
rect 3145 10217 3157 10220
rect 3191 10217 3203 10251
rect 3145 10211 3203 10217
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 4065 10251 4123 10257
rect 4065 10248 4077 10251
rect 3476 10220 4077 10248
rect 3476 10208 3482 10220
rect 4065 10217 4077 10220
rect 4111 10217 4123 10251
rect 4065 10211 4123 10217
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10248 5319 10251
rect 5534 10248 5540 10260
rect 5307 10220 5540 10248
rect 5307 10217 5319 10220
rect 5261 10211 5319 10217
rect 5534 10208 5540 10220
rect 5592 10248 5598 10260
rect 5905 10251 5963 10257
rect 5905 10248 5917 10251
rect 5592 10220 5917 10248
rect 5592 10208 5598 10220
rect 5905 10217 5917 10220
rect 5951 10217 5963 10251
rect 5905 10211 5963 10217
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 6822 10248 6828 10260
rect 6503 10220 6828 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7101 10251 7159 10257
rect 7101 10248 7113 10251
rect 7064 10220 7113 10248
rect 7064 10208 7070 10220
rect 7101 10217 7113 10220
rect 7147 10217 7159 10251
rect 7101 10211 7159 10217
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 7248 10220 7481 10248
rect 7248 10208 7254 10220
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 8110 10248 8116 10260
rect 8071 10220 8116 10248
rect 7469 10211 7527 10217
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8846 10208 8852 10260
rect 8904 10248 8910 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8904 10220 8953 10248
rect 8904 10208 8910 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 8941 10211 8999 10217
rect 10229 10251 10287 10257
rect 10229 10217 10241 10251
rect 10275 10248 10287 10251
rect 10962 10248 10968 10260
rect 10275 10220 10968 10248
rect 10275 10217 10287 10220
rect 10229 10211 10287 10217
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 11480 10220 11713 10248
rect 11480 10208 11486 10220
rect 11701 10217 11713 10220
rect 11747 10217 11759 10251
rect 11701 10211 11759 10217
rect 6917 10183 6975 10189
rect 6917 10149 6929 10183
rect 6963 10180 6975 10183
rect 7558 10180 7564 10192
rect 6963 10152 7564 10180
rect 6963 10149 6975 10152
rect 6917 10143 6975 10149
rect 7558 10140 7564 10152
rect 7616 10140 7622 10192
rect 8294 10140 8300 10192
rect 8352 10180 8358 10192
rect 8665 10183 8723 10189
rect 8665 10180 8677 10183
rect 8352 10152 8677 10180
rect 8352 10140 8358 10152
rect 8665 10149 8677 10152
rect 8711 10180 8723 10183
rect 9030 10180 9036 10192
rect 8711 10152 9036 10180
rect 8711 10149 8723 10152
rect 8665 10143 8723 10149
rect 9030 10140 9036 10152
rect 9088 10140 9094 10192
rect 10588 10183 10646 10189
rect 10588 10149 10600 10183
rect 10634 10180 10646 10183
rect 10778 10180 10784 10192
rect 10634 10152 10784 10180
rect 10634 10149 10646 10152
rect 10588 10143 10646 10149
rect 10778 10140 10784 10152
rect 10836 10180 10842 10192
rect 12805 10183 12863 10189
rect 12805 10180 12817 10183
rect 10836 10152 12817 10180
rect 10836 10140 10842 10152
rect 12805 10149 12817 10152
rect 12851 10180 12863 10183
rect 12986 10180 12992 10192
rect 12851 10152 12992 10180
rect 12851 10149 12863 10152
rect 12805 10143 12863 10149
rect 12986 10140 12992 10152
rect 13044 10140 13050 10192
rect 2038 10121 2044 10124
rect 2032 10112 2044 10121
rect 1999 10084 2044 10112
rect 2032 10075 2044 10084
rect 2038 10072 2044 10075
rect 2096 10072 2102 10124
rect 3513 10115 3571 10121
rect 3513 10081 3525 10115
rect 3559 10112 3571 10115
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 3559 10084 4445 10112
rect 3559 10081 3571 10084
rect 3513 10075 3571 10081
rect 4433 10081 4445 10084
rect 4479 10112 4491 10115
rect 5442 10112 5448 10124
rect 4479 10084 5448 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 5810 10112 5816 10124
rect 5771 10084 5816 10112
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 8478 10072 8484 10124
rect 8536 10112 8542 10124
rect 9306 10112 9312 10124
rect 8536 10084 9312 10112
rect 8536 10072 8542 10084
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 10321 10115 10379 10121
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 10410 10112 10416 10124
rect 10367 10084 10416 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10044 3939 10047
rect 4522 10044 4528 10056
rect 3927 10016 4528 10044
rect 3927 10013 3939 10016
rect 3881 10007 3939 10013
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 7558 10044 7564 10056
rect 4672 10016 4717 10044
rect 7519 10016 7564 10044
rect 4672 10004 4678 10016
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 8846 10044 8852 10056
rect 7791 10016 8852 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 5074 9936 5080 9988
rect 5132 9976 5138 9988
rect 5629 9979 5687 9985
rect 5629 9976 5641 9979
rect 5132 9948 5641 9976
rect 5132 9936 5138 9948
rect 5629 9945 5641 9948
rect 5675 9945 5687 9979
rect 5629 9939 5687 9945
rect 9306 9908 9312 9920
rect 9267 9880 9312 9908
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12492 9880 12537 9908
rect 12492 9868 12498 9880
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 3050 9664 3056 9716
rect 3108 9704 3114 9716
rect 3142 9704 3148 9716
rect 3108 9676 3148 9704
rect 3108 9664 3114 9676
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4580 9676 4997 9704
rect 4580 9664 4586 9676
rect 4985 9673 4997 9676
rect 5031 9673 5043 9707
rect 7190 9704 7196 9716
rect 7151 9676 7196 9704
rect 4985 9667 5043 9673
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 7374 9664 7380 9716
rect 7432 9704 7438 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 7432 9676 7757 9704
rect 7432 9664 7438 9676
rect 7745 9673 7757 9676
rect 7791 9704 7803 9707
rect 9306 9704 9312 9716
rect 7791 9676 9312 9704
rect 7791 9673 7803 9676
rect 7745 9667 7803 9673
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10686 9704 10692 9716
rect 10468 9676 10692 9704
rect 10468 9664 10474 9676
rect 10686 9664 10692 9676
rect 10744 9704 10750 9716
rect 10744 9676 11100 9704
rect 10744 9664 10750 9676
rect 1857 9639 1915 9645
rect 1857 9605 1869 9639
rect 1903 9636 1915 9639
rect 2038 9636 2044 9648
rect 1903 9608 2044 9636
rect 1903 9605 1915 9608
rect 1857 9599 1915 9605
rect 2038 9596 2044 9608
rect 2096 9596 2102 9648
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 4157 9639 4215 9645
rect 4157 9636 4169 9639
rect 3936 9608 4169 9636
rect 3936 9596 3942 9608
rect 4157 9605 4169 9608
rect 4203 9636 4215 9639
rect 4614 9636 4620 9648
rect 4203 9608 4620 9636
rect 4203 9605 4215 9608
rect 4157 9599 4215 9605
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 6641 9639 6699 9645
rect 6641 9605 6653 9639
rect 6687 9636 6699 9639
rect 8846 9636 8852 9648
rect 6687 9608 8852 9636
rect 6687 9605 6699 9608
rect 6641 9599 6699 9605
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5500 9540 5549 9568
rect 5500 9528 5506 9540
rect 5537 9537 5549 9540
rect 5583 9568 5595 9571
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5583 9540 6009 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 5997 9537 6009 9540
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 8110 9568 8116 9580
rect 7340 9540 8116 9568
rect 7340 9528 7346 9540
rect 8110 9528 8116 9540
rect 8168 9568 8174 9580
rect 8404 9577 8432 9608
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 10873 9639 10931 9645
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 10962 9636 10968 9648
rect 10919 9608 10968 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 11072 9636 11100 9676
rect 11149 9639 11207 9645
rect 11149 9636 11161 9639
rect 11072 9608 11161 9636
rect 11149 9605 11161 9608
rect 11195 9605 11207 9639
rect 11149 9599 11207 9605
rect 8205 9571 8263 9577
rect 8205 9568 8217 9571
rect 8168 9540 8217 9568
rect 8168 9528 8174 9540
rect 8205 9537 8217 9540
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10778 9568 10784 9580
rect 10459 9540 10784 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2682 9500 2688 9512
rect 2363 9472 2688 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2682 9460 2688 9472
rect 2740 9500 2746 9512
rect 2777 9503 2835 9509
rect 2777 9500 2789 9503
rect 2740 9472 2789 9500
rect 2740 9460 2746 9472
rect 2777 9469 2789 9472
rect 2823 9469 2835 9503
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 2777 9463 2835 9469
rect 9140 9472 9505 9500
rect 9140 9444 9168 9472
rect 9493 9469 9505 9472
rect 9539 9500 9551 9503
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 9539 9472 9781 9500
rect 9539 9469 9551 9472
rect 9493 9463 9551 9469
rect 9769 9469 9781 9472
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 3044 9435 3102 9441
rect 3044 9401 3056 9435
rect 3090 9432 3102 9435
rect 5258 9432 5264 9444
rect 3090 9404 3124 9432
rect 4632 9404 5264 9432
rect 3090 9401 3102 9404
rect 3044 9395 3102 9401
rect 2685 9367 2743 9373
rect 2685 9333 2697 9367
rect 2731 9364 2743 9367
rect 3059 9364 3087 9395
rect 4632 9376 4660 9404
rect 5258 9392 5264 9404
rect 5316 9432 5322 9444
rect 5445 9435 5503 9441
rect 5445 9432 5457 9435
rect 5316 9404 5457 9432
rect 5316 9392 5322 9404
rect 5445 9401 5457 9404
rect 5491 9401 5503 9435
rect 9122 9432 9128 9444
rect 9083 9404 9128 9432
rect 5445 9395 5503 9401
rect 9122 9392 9128 9404
rect 9180 9392 9186 9444
rect 3234 9364 3240 9376
rect 2731 9336 3240 9364
rect 2731 9333 2743 9336
rect 2685 9327 2743 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 4614 9364 4620 9376
rect 4571 9336 4620 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4893 9367 4951 9373
rect 4893 9333 4905 9367
rect 4939 9364 4951 9367
rect 4982 9364 4988 9376
rect 4939 9336 4988 9364
rect 4939 9333 4951 9336
rect 4893 9327 4951 9333
rect 4982 9324 4988 9336
rect 5040 9364 5046 9376
rect 5350 9364 5356 9376
rect 5040 9336 5356 9364
rect 5040 9324 5046 9336
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 7653 9367 7711 9373
rect 7653 9333 7665 9367
rect 7699 9364 7711 9367
rect 8110 9364 8116 9376
rect 7699 9336 8116 9364
rect 7699 9333 7711 9336
rect 7653 9327 7711 9333
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 9306 9364 9312 9376
rect 9267 9336 9312 9364
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 1762 9160 1768 9172
rect 1723 9132 1768 9160
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 2363 9132 2881 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 2869 9129 2881 9132
rect 2915 9160 2927 9163
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 2915 9132 4077 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 5592 9132 5641 9160
rect 5592 9120 5598 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 5629 9123 5687 9129
rect 5994 9120 6000 9172
rect 6052 9120 6058 9172
rect 6089 9163 6147 9169
rect 6089 9129 6101 9163
rect 6135 9160 6147 9163
rect 6178 9160 6184 9172
rect 6135 9132 6184 9160
rect 6135 9129 6147 9132
rect 6089 9123 6147 9129
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6914 9160 6920 9172
rect 6875 9132 6920 9160
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7558 9160 7564 9172
rect 7331 9132 7564 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7558 9120 7564 9132
rect 7616 9160 7622 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 7616 9132 9689 9160
rect 7616 9120 7622 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 10008 9132 10057 9160
rect 10008 9120 10014 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10226 9160 10232 9172
rect 10183 9132 10232 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 2777 9095 2835 9101
rect 2777 9092 2789 9095
rect 2556 9064 2789 9092
rect 2556 9052 2562 9064
rect 2777 9061 2789 9064
rect 2823 9092 2835 9095
rect 6012 9092 6040 9120
rect 2823 9064 6040 9092
rect 2823 9061 2835 9064
rect 2777 9055 2835 9061
rect 3326 8984 3332 9036
rect 3384 9024 3390 9036
rect 3878 9024 3884 9036
rect 3384 8996 3884 9024
rect 3384 8984 3390 8996
rect 3878 8984 3884 8996
rect 3936 8984 3942 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4982 9024 4988 9036
rect 4479 8996 4988 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5994 9024 6000 9036
rect 5955 8996 6000 9024
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 7644 9027 7702 9033
rect 7644 8993 7656 9027
rect 7690 9024 7702 9027
rect 8202 9024 8208 9036
rect 7690 8996 8208 9024
rect 7690 8993 7702 8996
rect 7644 8987 7702 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3234 8956 3240 8968
rect 3099 8928 3240 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3234 8916 3240 8928
rect 3292 8956 3298 8968
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 3292 8928 3433 8956
rect 3292 8916 3298 8928
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 4522 8956 4528 8968
rect 4483 8928 4528 8956
rect 3421 8919 3479 8925
rect 3436 8888 3464 8919
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 4798 8956 4804 8968
rect 4755 8928 4804 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 4798 8916 4804 8928
rect 4856 8956 4862 8968
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 4856 8928 5089 8956
rect 4856 8916 4862 8928
rect 5077 8925 5089 8928
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8925 6239 8959
rect 7374 8956 7380 8968
rect 7335 8928 7380 8956
rect 6181 8919 6239 8925
rect 5442 8888 5448 8900
rect 3436 8860 5448 8888
rect 5442 8848 5448 8860
rect 5500 8888 5506 8900
rect 6196 8888 6224 8919
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 9490 8956 9496 8968
rect 9364 8928 9496 8956
rect 9364 8916 9370 8928
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 10284 8928 10329 8956
rect 10284 8916 10290 8928
rect 5500 8860 6224 8888
rect 8757 8891 8815 8897
rect 5500 8848 5506 8860
rect 8757 8857 8769 8891
rect 8803 8888 8815 8891
rect 8846 8888 8852 8900
rect 8803 8860 8852 8888
rect 8803 8857 8815 8860
rect 8757 8851 8815 8857
rect 8846 8848 8852 8860
rect 8904 8848 8910 8900
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8820 2467 8823
rect 2774 8820 2780 8832
rect 2455 8792 2780 8820
rect 2455 8789 2467 8792
rect 2409 8783 2467 8789
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 5902 8820 5908 8832
rect 4580 8792 5908 8820
rect 4580 8780 4586 8792
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 9217 8823 9275 8829
rect 9217 8789 9229 8823
rect 9263 8820 9275 8823
rect 9490 8820 9496 8832
rect 9263 8792 9496 8820
rect 9263 8789 9275 8792
rect 9217 8783 9275 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 2498 8616 2504 8628
rect 2459 8588 2504 8616
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4522 8616 4528 8628
rect 4203 8588 4528 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4522 8576 4528 8588
rect 4580 8576 4586 8628
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 5629 8619 5687 8625
rect 5629 8616 5641 8619
rect 5500 8588 5641 8616
rect 5500 8576 5506 8588
rect 5629 8585 5641 8588
rect 5675 8585 5687 8619
rect 5629 8579 5687 8585
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 5868 8588 6469 8616
rect 5868 8576 5874 8588
rect 6457 8585 6469 8588
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 5997 8551 6055 8557
rect 5997 8517 6009 8551
rect 6043 8548 6055 8551
rect 6178 8548 6184 8560
rect 6043 8520 6184 8548
rect 6043 8517 6055 8520
rect 5997 8511 6055 8517
rect 6178 8508 6184 8520
rect 6236 8508 6242 8560
rect 6638 8508 6644 8560
rect 6696 8548 6702 8560
rect 6696 8520 6868 8548
rect 6696 8508 6702 8520
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 3234 8480 3240 8492
rect 3195 8452 3240 8480
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1670 8412 1676 8424
rect 1443 8384 1676 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1670 8372 1676 8384
rect 1728 8412 1734 8424
rect 2130 8412 2136 8424
rect 1728 8384 2136 8412
rect 1728 8372 1734 8384
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 2682 8372 2688 8424
rect 2740 8412 2746 8424
rect 4249 8415 4307 8421
rect 4249 8412 4261 8415
rect 2740 8384 4261 8412
rect 2740 8372 2746 8384
rect 4249 8381 4261 8384
rect 4295 8412 4307 8415
rect 5350 8412 5356 8424
rect 4295 8384 5356 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 6840 8421 6868 8520
rect 7098 8421 7104 8424
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 7092 8412 7104 8421
rect 6871 8384 6960 8412
rect 7059 8384 7104 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 3053 8347 3111 8353
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 3786 8344 3792 8356
rect 3099 8316 3792 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 4154 8304 4160 8356
rect 4212 8344 4218 8356
rect 4516 8347 4574 8353
rect 4516 8344 4528 8347
rect 4212 8316 4528 8344
rect 4212 8304 4218 8316
rect 4516 8313 4528 8316
rect 4562 8344 4574 8347
rect 4798 8344 4804 8356
rect 4562 8316 4804 8344
rect 4562 8313 4574 8316
rect 4516 8307 4574 8313
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5534 8304 5540 8356
rect 5592 8344 5598 8356
rect 5994 8344 6000 8356
rect 5592 8316 6000 8344
rect 5592 8304 5598 8316
rect 5994 8304 6000 8316
rect 6052 8344 6058 8356
rect 6273 8347 6331 8353
rect 6273 8344 6285 8347
rect 6052 8316 6285 8344
rect 6052 8304 6058 8316
rect 6273 8313 6285 8316
rect 6319 8313 6331 8347
rect 6656 8344 6684 8375
rect 6932 8344 6960 8384
rect 7092 8375 7104 8384
rect 7098 8372 7104 8375
rect 7156 8372 7162 8424
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 7432 8384 9137 8412
rect 7432 8372 7438 8384
rect 7392 8344 7420 8372
rect 6656 8316 6868 8344
rect 6932 8316 7420 8344
rect 6273 8307 6331 8313
rect 2685 8279 2743 8285
rect 2685 8245 2697 8279
rect 2731 8276 2743 8279
rect 2866 8276 2872 8288
rect 2731 8248 2872 8276
rect 2731 8245 2743 8248
rect 2685 8239 2743 8245
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3145 8279 3203 8285
rect 3145 8245 3157 8279
rect 3191 8276 3203 8279
rect 3418 8276 3424 8288
rect 3191 8248 3424 8276
rect 3191 8245 3203 8248
rect 3145 8239 3203 8245
rect 3418 8236 3424 8248
rect 3476 8236 3482 8288
rect 6840 8276 6868 8316
rect 8772 8288 8800 8384
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 9381 8415 9439 8421
rect 9381 8412 9393 8415
rect 9272 8384 9393 8412
rect 9272 8372 9278 8384
rect 9381 8381 9393 8384
rect 9427 8381 9439 8415
rect 9950 8412 9956 8424
rect 9381 8375 9439 8381
rect 9508 8384 9956 8412
rect 9033 8347 9091 8353
rect 9033 8313 9045 8347
rect 9079 8344 9091 8347
rect 9508 8344 9536 8384
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 9079 8316 9536 8344
rect 9079 8313 9091 8316
rect 9033 8307 9091 8313
rect 7558 8276 7564 8288
rect 6840 8248 7564 8276
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 8202 8276 8208 8288
rect 8163 8248 8208 8276
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8665 8279 8723 8285
rect 8665 8245 8677 8279
rect 8711 8276 8723 8279
rect 8754 8276 8760 8288
rect 8711 8248 8760 8276
rect 8711 8245 8723 8248
rect 8665 8239 8723 8245
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 10505 8279 10563 8285
rect 10505 8276 10517 8279
rect 8996 8248 10517 8276
rect 8996 8236 9002 8248
rect 10505 8245 10517 8248
rect 10551 8245 10563 8279
rect 10505 8239 10563 8245
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 11974 8276 11980 8288
rect 11480 8248 11980 8276
rect 11480 8236 11486 8248
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 1670 8072 1676 8084
rect 1631 8044 1676 8072
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 2406 8072 2412 8084
rect 2367 8044 2412 8072
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 2869 8075 2927 8081
rect 2869 8072 2881 8075
rect 2832 8044 2881 8072
rect 2832 8032 2838 8044
rect 2869 8041 2881 8044
rect 2915 8041 2927 8075
rect 2869 8035 2927 8041
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4062 8072 4068 8084
rect 3927 8044 4068 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 5534 8072 5540 8084
rect 4387 8044 5540 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 6733 8075 6791 8081
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 6822 8072 6828 8084
rect 6779 8044 6828 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 7469 8075 7527 8081
rect 7469 8041 7481 8075
rect 7515 8072 7527 8075
rect 8202 8072 8208 8084
rect 7515 8044 8208 8072
rect 7515 8041 7527 8044
rect 7469 8035 7527 8041
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 10226 8072 10232 8084
rect 10187 8044 10232 8072
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 13262 8072 13268 8084
rect 12124 8044 13268 8072
rect 12124 8032 12130 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 2317 8007 2375 8013
rect 2317 7973 2329 8007
rect 2363 8004 2375 8007
rect 3234 8004 3240 8016
rect 2363 7976 3240 8004
rect 2363 7973 2375 7976
rect 2317 7967 2375 7973
rect 3234 7964 3240 7976
rect 3292 7964 3298 8016
rect 4893 8007 4951 8013
rect 4893 7973 4905 8007
rect 4939 8004 4951 8007
rect 4982 8004 4988 8016
rect 4939 7976 4988 8004
rect 4939 7973 4951 7976
rect 4893 7967 4951 7973
rect 4982 7964 4988 7976
rect 5040 7964 5046 8016
rect 7101 8007 7159 8013
rect 7101 7973 7113 8007
rect 7147 8004 7159 8007
rect 7558 8004 7564 8016
rect 7147 7976 7564 8004
rect 7147 7973 7159 7976
rect 7101 7967 7159 7973
rect 7558 7964 7564 7976
rect 7616 7964 7622 8016
rect 7929 8007 7987 8013
rect 7929 7973 7941 8007
rect 7975 8004 7987 8007
rect 9214 8004 9220 8016
rect 7975 7976 9220 8004
rect 7975 7973 7987 7976
rect 7929 7967 7987 7973
rect 9214 7964 9220 7976
rect 9272 8004 9278 8016
rect 9401 8007 9459 8013
rect 9401 8004 9413 8007
rect 9272 7976 9413 8004
rect 9272 7964 9278 7976
rect 9401 7973 9413 7976
rect 9447 8004 9459 8007
rect 9490 8004 9496 8016
rect 9447 7976 9496 8004
rect 9447 7973 9459 7976
rect 9401 7967 9459 7973
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 2866 7936 2872 7948
rect 2823 7908 2872 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 2866 7896 2872 7908
rect 2924 7936 2930 7948
rect 3142 7936 3148 7948
rect 2924 7908 3148 7936
rect 2924 7896 2930 7908
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 5609 7939 5667 7945
rect 5609 7936 5621 7939
rect 5500 7908 5621 7936
rect 5500 7896 5506 7908
rect 5609 7905 5621 7908
rect 5655 7936 5667 7939
rect 6086 7936 6092 7948
rect 5655 7908 6092 7936
rect 5655 7905 5667 7908
rect 5609 7899 5667 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8846 7936 8852 7948
rect 8435 7908 8852 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3326 7868 3332 7880
rect 3099 7840 3332 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 5350 7868 5356 7880
rect 5311 7840 5356 7868
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 8481 7871 8539 7877
rect 8481 7868 8493 7871
rect 7892 7840 8493 7868
rect 7892 7828 7898 7840
rect 8481 7837 8493 7840
rect 8527 7837 8539 7871
rect 8665 7871 8723 7877
rect 8665 7868 8677 7871
rect 8481 7831 8539 7837
rect 8588 7840 8677 7868
rect 3418 7692 3424 7744
rect 3476 7732 3482 7744
rect 3513 7735 3571 7741
rect 3513 7732 3525 7735
rect 3476 7704 3525 7732
rect 3476 7692 3482 7704
rect 3513 7701 3525 7704
rect 3559 7732 3571 7735
rect 4062 7732 4068 7744
rect 3559 7704 4068 7732
rect 3559 7701 3571 7704
rect 3513 7695 3571 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8202 7732 8208 7744
rect 8067 7704 8208 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8588 7732 8616 7840
rect 8665 7837 8677 7840
rect 8711 7868 8723 7871
rect 8938 7868 8944 7880
rect 8711 7840 8944 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9416 7800 9444 7967
rect 9490 7964 9496 7976
rect 9548 7964 9554 8016
rect 9950 8004 9956 8016
rect 9863 7976 9956 8004
rect 9950 7964 9956 7976
rect 10008 8004 10014 8016
rect 10134 8004 10140 8016
rect 10008 7976 10140 8004
rect 10008 7964 10014 7976
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 10597 7939 10655 7945
rect 10597 7905 10609 7939
rect 10643 7936 10655 7939
rect 10870 7936 10876 7948
rect 10643 7908 10876 7936
rect 10643 7905 10655 7908
rect 10597 7899 10655 7905
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 11054 7896 11060 7948
rect 11112 7936 11118 7948
rect 11221 7939 11279 7945
rect 11221 7936 11233 7939
rect 11112 7908 11233 7936
rect 11112 7896 11118 7908
rect 11221 7905 11233 7908
rect 11267 7905 11279 7939
rect 11221 7899 11279 7905
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 10428 7840 10977 7868
rect 10226 7800 10232 7812
rect 9416 7772 10232 7800
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 8662 7732 8668 7744
rect 8588 7704 8668 7732
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 8812 7704 9137 7732
rect 8812 7692 8818 7704
rect 9125 7701 9137 7704
rect 9171 7732 9183 7735
rect 9582 7732 9588 7744
rect 9171 7704 9588 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 9582 7692 9588 7704
rect 9640 7732 9646 7744
rect 10428 7741 10456 7840
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 10413 7735 10471 7741
rect 10413 7732 10425 7735
rect 9640 7704 10425 7732
rect 9640 7692 9646 7704
rect 10413 7701 10425 7704
rect 10459 7701 10471 7735
rect 12342 7732 12348 7744
rect 12303 7704 12348 7732
rect 10413 7695 10471 7701
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 3142 7528 3148 7540
rect 2832 7500 2877 7528
rect 3103 7500 3148 7528
rect 2832 7488 2838 7500
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 5074 7528 5080 7540
rect 4755 7500 5080 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 2501 7463 2559 7469
rect 2501 7429 2513 7463
rect 2547 7460 2559 7463
rect 3326 7460 3332 7472
rect 2547 7432 3332 7460
rect 2547 7429 2559 7432
rect 2501 7423 2559 7429
rect 3326 7420 3332 7432
rect 3384 7420 3390 7472
rect 5000 7333 5028 7500
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5442 7528 5448 7540
rect 5403 7500 5448 7528
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 6178 7528 6184 7540
rect 6139 7500 6184 7528
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 6638 7528 6644 7540
rect 6599 7500 6644 7528
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7834 7528 7840 7540
rect 7795 7500 7840 7528
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 10505 7531 10563 7537
rect 10505 7497 10517 7531
rect 10551 7528 10563 7531
rect 10870 7528 10876 7540
rect 10551 7500 10876 7528
rect 10551 7497 10563 7500
rect 10505 7491 10563 7497
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 11054 7528 11060 7540
rect 11015 7500 11060 7528
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 8757 7463 8815 7469
rect 8757 7460 8769 7463
rect 5960 7432 8769 7460
rect 5960 7420 5966 7432
rect 8757 7429 8769 7432
rect 8803 7429 8815 7463
rect 8938 7460 8944 7472
rect 8899 7432 8944 7460
rect 8757 7423 8815 7429
rect 8938 7420 8944 7432
rect 8996 7420 9002 7472
rect 8481 7395 8539 7401
rect 8481 7361 8493 7395
rect 8527 7392 8539 7395
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 8527 7364 10057 7392
rect 8527 7361 8539 7364
rect 8481 7355 8539 7361
rect 10045 7361 10057 7364
rect 10091 7392 10103 7395
rect 10226 7392 10232 7404
rect 10091 7364 10232 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 10226 7352 10232 7364
rect 10284 7392 10290 7404
rect 12342 7392 12348 7404
rect 10284 7364 12348 7392
rect 10284 7352 10290 7364
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 4985 7327 5043 7333
rect 4985 7293 4997 7327
rect 5031 7293 5043 7327
rect 4985 7287 5043 7293
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7324 5687 7327
rect 6178 7324 6184 7336
rect 5675 7296 6184 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 8662 7324 8668 7336
rect 7423 7296 8668 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 9766 7284 9772 7336
rect 9824 7324 9830 7336
rect 10410 7324 10416 7336
rect 9824 7296 10416 7324
rect 9824 7284 9830 7296
rect 10410 7284 10416 7296
rect 10468 7284 10474 7336
rect 7466 7216 7472 7268
rect 7524 7256 7530 7268
rect 8205 7259 8263 7265
rect 8205 7256 8217 7259
rect 7524 7228 8217 7256
rect 7524 7216 7530 7228
rect 8205 7225 8217 7228
rect 8251 7225 8263 7259
rect 8205 7219 8263 7225
rect 8757 7259 8815 7265
rect 8757 7225 8769 7259
rect 8803 7256 8815 7259
rect 9861 7259 9919 7265
rect 9861 7256 9873 7259
rect 8803 7228 9873 7256
rect 8803 7225 8815 7228
rect 8757 7219 8815 7225
rect 9232 7200 9260 7228
rect 9861 7225 9873 7228
rect 9907 7225 9919 7259
rect 9861 7219 9919 7225
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 4387 7160 4813 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4801 7157 4813 7160
rect 4847 7188 4859 7191
rect 5442 7188 5448 7200
rect 4847 7160 5448 7188
rect 4847 7157 4859 7160
rect 4801 7151 4859 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5813 7191 5871 7197
rect 5813 7157 5825 7191
rect 5859 7188 5871 7191
rect 6086 7188 6092 7200
rect 5859 7160 6092 7188
rect 5859 7157 5871 7160
rect 5813 7151 5871 7157
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 6730 7148 6736 7200
rect 6788 7188 6794 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 6788 7160 7757 7188
rect 6788 7148 6794 7160
rect 7745 7157 7757 7160
rect 7791 7188 7803 7191
rect 8110 7188 8116 7200
rect 7791 7160 8116 7188
rect 7791 7157 7803 7160
rect 7745 7151 7803 7157
rect 8110 7148 8116 7160
rect 8168 7188 8174 7200
rect 8297 7191 8355 7197
rect 8297 7188 8309 7191
rect 8168 7160 8309 7188
rect 8168 7148 8174 7160
rect 8297 7157 8309 7160
rect 8343 7157 8355 7191
rect 9214 7188 9220 7200
rect 9175 7160 9220 7188
rect 8297 7151 8355 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 9398 7188 9404 7200
rect 9359 7160 9404 7188
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9766 7188 9772 7200
rect 9727 7160 9772 7188
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11020 7160 11345 7188
rect 11020 7148 11026 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 2038 6944 2044 6996
rect 2096 6984 2102 6996
rect 2133 6987 2191 6993
rect 2133 6984 2145 6987
rect 2096 6956 2145 6984
rect 2096 6944 2102 6956
rect 2133 6953 2145 6956
rect 2179 6984 2191 6987
rect 3418 6984 3424 6996
rect 2179 6956 3424 6984
rect 2179 6953 2191 6956
rect 2133 6947 2191 6953
rect 3418 6944 3424 6956
rect 3476 6944 3482 6996
rect 7193 6987 7251 6993
rect 7193 6953 7205 6987
rect 7239 6984 7251 6987
rect 7834 6984 7840 6996
rect 7239 6956 7840 6984
rect 7239 6953 7251 6956
rect 7193 6947 7251 6953
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 8481 6987 8539 6993
rect 8481 6953 8493 6987
rect 8527 6984 8539 6987
rect 8846 6984 8852 6996
rect 8527 6956 8852 6984
rect 8527 6953 8539 6956
rect 8481 6947 8539 6953
rect 8846 6944 8852 6956
rect 8904 6984 8910 6996
rect 9398 6984 9404 6996
rect 8904 6956 9404 6984
rect 8904 6944 8910 6956
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 10226 6984 10232 6996
rect 10187 6956 10232 6984
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 7466 6876 7472 6928
rect 7524 6916 7530 6928
rect 7929 6919 7987 6925
rect 7929 6916 7941 6919
rect 7524 6888 7941 6916
rect 7524 6876 7530 6888
rect 7929 6885 7941 6888
rect 7975 6885 7987 6919
rect 9766 6916 9772 6928
rect 7929 6879 7987 6885
rect 9416 6888 9772 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1578 6848 1584 6860
rect 1443 6820 1584 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 2498 6848 2504 6860
rect 2459 6820 2504 6848
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 5074 6848 5080 6860
rect 5035 6820 5080 6848
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 6178 6848 6184 6860
rect 6139 6820 6184 6848
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 7561 6851 7619 6857
rect 7561 6817 7573 6851
rect 7607 6848 7619 6851
rect 8386 6848 8392 6860
rect 7607 6820 8392 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 8754 6848 8760 6860
rect 8536 6820 8760 6848
rect 8536 6808 8542 6820
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8662 6780 8668 6792
rect 7984 6752 8668 6780
rect 7984 6740 7990 6752
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 566 6672 572 6724
rect 624 6712 630 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 624 6684 2697 6712
rect 624 6672 630 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 4890 6672 4896 6724
rect 4948 6712 4954 6724
rect 6365 6715 6423 6721
rect 6365 6712 6377 6715
rect 4948 6684 6377 6712
rect 4948 6672 4954 6684
rect 6365 6681 6377 6684
rect 6411 6681 6423 6715
rect 6365 6675 6423 6681
rect 8294 6672 8300 6724
rect 8352 6712 8358 6724
rect 9416 6721 9444 6888
rect 9766 6876 9772 6888
rect 9824 6876 9830 6928
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9548 6820 9689 6848
rect 9548 6808 9554 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 11020 6820 11069 6848
rect 11020 6808 11026 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11313 6851 11371 6857
rect 11313 6848 11325 6851
rect 11204 6820 11325 6848
rect 11204 6808 11210 6820
rect 11313 6817 11325 6820
rect 11359 6817 11371 6851
rect 11313 6811 11371 6817
rect 9401 6715 9459 6721
rect 9401 6712 9413 6715
rect 8352 6684 9413 6712
rect 8352 6672 8358 6684
rect 9401 6681 9413 6684
rect 9447 6681 9459 6715
rect 9401 6675 9459 6681
rect 1302 6604 1308 6656
rect 1360 6644 1366 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1360 6616 1593 6644
rect 1360 6604 1366 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 5258 6644 5264 6656
rect 5219 6616 5264 6644
rect 1581 6607 1639 6613
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 5721 6647 5779 6653
rect 5721 6644 5733 6647
rect 5500 6616 5733 6644
rect 5500 6604 5506 6616
rect 5721 6613 5733 6616
rect 5767 6644 5779 6647
rect 5902 6644 5908 6656
rect 5767 6616 5908 6644
rect 5767 6613 5779 6616
rect 5721 6607 5779 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 8021 6647 8079 6653
rect 8021 6613 8033 6647
rect 8067 6644 8079 6647
rect 8478 6644 8484 6656
rect 8067 6616 8484 6644
rect 8067 6613 8079 6616
rect 8021 6607 8079 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9858 6644 9864 6656
rect 9819 6616 9864 6644
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 11974 6644 11980 6656
rect 11112 6616 11980 6644
rect 11112 6604 11118 6616
rect 11974 6604 11980 6616
rect 12032 6644 12038 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 12032 6616 12449 6644
rect 12032 6604 12038 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 12437 6607 12495 6613
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6440 1642 6452
rect 1636 6412 2452 6440
rect 1636 6400 1642 6412
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 2225 6375 2283 6381
rect 2225 6372 2237 6375
rect 1452 6344 2237 6372
rect 1452 6332 1458 6344
rect 2225 6341 2237 6344
rect 2271 6341 2283 6375
rect 2225 6335 2283 6341
rect 2424 6304 2452 6412
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 2593 6443 2651 6449
rect 2593 6440 2605 6443
rect 2556 6412 2605 6440
rect 2556 6400 2562 6412
rect 2593 6409 2605 6412
rect 2639 6409 2651 6443
rect 2593 6403 2651 6409
rect 4982 6400 4988 6452
rect 5040 6440 5046 6452
rect 5077 6443 5135 6449
rect 5077 6440 5089 6443
rect 5040 6412 5089 6440
rect 5040 6400 5046 6412
rect 5077 6409 5089 6412
rect 5123 6409 5135 6443
rect 5534 6440 5540 6452
rect 5495 6412 5540 6440
rect 5077 6403 5135 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 6178 6440 6184 6452
rect 6139 6412 6184 6440
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 6638 6440 6644 6452
rect 6599 6412 6644 6440
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 7561 6443 7619 6449
rect 7561 6409 7573 6443
rect 7607 6440 7619 6443
rect 8018 6440 8024 6452
rect 7607 6412 8024 6440
rect 7607 6409 7619 6412
rect 7561 6403 7619 6409
rect 4709 6375 4767 6381
rect 4709 6341 4721 6375
rect 4755 6372 4767 6375
rect 5718 6372 5724 6384
rect 4755 6344 5724 6372
rect 4755 6341 4767 6344
rect 4709 6335 4767 6341
rect 5718 6332 5724 6344
rect 5776 6332 5782 6384
rect 6178 6304 6184 6316
rect 2424 6276 6184 6304
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 2038 6236 2044 6248
rect 1999 6208 2044 6236
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 4430 6236 4436 6248
rect 4391 6208 4436 6236
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4525 6239 4583 6245
rect 4525 6205 4537 6239
rect 4571 6236 4583 6239
rect 4706 6236 4712 6248
rect 4571 6208 4712 6236
rect 4571 6205 4583 6208
rect 4525 6199 4583 6205
rect 4706 6196 4712 6208
rect 4764 6236 4770 6248
rect 4982 6236 4988 6248
rect 4764 6208 4988 6236
rect 4764 6196 4770 6208
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 5629 6239 5687 6245
rect 5629 6236 5641 6239
rect 5592 6208 5641 6236
rect 5592 6196 5598 6208
rect 5629 6205 5641 6208
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6236 6975 6239
rect 7576 6236 7604 6403
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 8444 6412 9597 6440
rect 8444 6400 8450 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 9585 6403 9643 6409
rect 11057 6443 11115 6449
rect 11057 6409 11069 6443
rect 11103 6440 11115 6443
rect 11146 6440 11152 6452
rect 11103 6412 11152 6440
rect 11103 6409 11115 6412
rect 11057 6403 11115 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 7926 6372 7932 6384
rect 7887 6344 7932 6372
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 9125 6375 9183 6381
rect 9125 6341 9137 6375
rect 9171 6372 9183 6375
rect 9490 6372 9496 6384
rect 9171 6344 9496 6372
rect 9171 6341 9183 6344
rect 9125 6335 9183 6341
rect 9490 6332 9496 6344
rect 9548 6332 9554 6384
rect 7944 6304 7972 6332
rect 8662 6304 8668 6316
rect 7944 6276 8524 6304
rect 8623 6276 8668 6304
rect 6963 6208 7604 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 8294 6196 8300 6248
rect 8352 6236 8358 6248
rect 8389 6239 8447 6245
rect 8389 6236 8401 6239
rect 8352 6208 8401 6236
rect 8352 6196 8358 6208
rect 8389 6205 8401 6208
rect 8435 6205 8447 6239
rect 8496 6236 8524 6276
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 10226 6304 10232 6316
rect 10187 6276 10232 6304
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 8570 6236 8576 6248
rect 8496 6208 8576 6236
rect 8389 6199 8447 6205
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9732 6208 9965 6236
rect 9732 6196 9738 6208
rect 9953 6205 9965 6208
rect 9999 6236 10011 6239
rect 10597 6239 10655 6245
rect 10597 6236 10609 6239
rect 9999 6208 10609 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10597 6205 10609 6208
rect 10643 6205 10655 6239
rect 10597 6199 10655 6205
rect 11149 6239 11207 6245
rect 11149 6205 11161 6239
rect 11195 6236 11207 6239
rect 11514 6236 11520 6248
rect 11195 6208 11520 6236
rect 11195 6205 11207 6208
rect 11149 6199 11207 6205
rect 11514 6196 11520 6208
rect 11572 6236 11578 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11572 6208 11713 6236
rect 11572 6196 11578 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 5813 6103 5871 6109
rect 5813 6100 5825 6103
rect 5592 6072 5825 6100
rect 5592 6060 5598 6072
rect 5813 6069 5825 6072
rect 5859 6069 5871 6103
rect 5813 6063 5871 6069
rect 7006 6060 7012 6112
rect 7064 6100 7070 6112
rect 7101 6103 7159 6109
rect 7101 6100 7113 6103
rect 7064 6072 7113 6100
rect 7064 6060 7070 6072
rect 7101 6069 7113 6072
rect 7147 6069 7159 6103
rect 7101 6063 7159 6069
rect 7926 6060 7932 6112
rect 7984 6100 7990 6112
rect 8021 6103 8079 6109
rect 8021 6100 8033 6103
rect 7984 6072 8033 6100
rect 7984 6060 7990 6072
rect 8021 6069 8033 6072
rect 8067 6069 8079 6103
rect 8021 6063 8079 6069
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 9490 6100 9496 6112
rect 8536 6072 8581 6100
rect 9403 6072 9496 6100
rect 8536 6060 8542 6072
rect 9490 6060 9496 6072
rect 9548 6100 9554 6112
rect 9766 6100 9772 6112
rect 9548 6072 9772 6100
rect 9548 6060 9554 6072
rect 9766 6060 9772 6072
rect 9824 6100 9830 6112
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 9824 6072 10057 6100
rect 9824 6060 9830 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 11112 6072 11345 6100
rect 11112 6060 11118 6072
rect 11333 6069 11345 6072
rect 11379 6069 11391 6103
rect 11333 6063 11391 6069
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 6273 5899 6331 5905
rect 6273 5865 6285 5899
rect 6319 5896 6331 5899
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 6319 5868 7849 5896
rect 6319 5865 6331 5868
rect 6273 5859 6331 5865
rect 7837 5865 7849 5868
rect 7883 5896 7895 5899
rect 9677 5899 9735 5905
rect 9677 5896 9689 5899
rect 7883 5868 9689 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 9677 5865 9689 5868
rect 9723 5865 9735 5899
rect 9677 5859 9735 5865
rect 9766 5856 9772 5908
rect 9824 5896 9830 5908
rect 10781 5899 10839 5905
rect 10781 5896 10793 5899
rect 9824 5868 10793 5896
rect 9824 5856 9830 5868
rect 10781 5865 10793 5868
rect 10827 5896 10839 5899
rect 10962 5896 10968 5908
rect 10827 5868 10968 5896
rect 10827 5865 10839 5868
rect 10781 5859 10839 5865
rect 10962 5856 10968 5868
rect 11020 5896 11026 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 11020 5868 11069 5896
rect 11020 5856 11026 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 11333 5899 11391 5905
rect 11333 5896 11345 5899
rect 11296 5868 11345 5896
rect 11296 5856 11302 5868
rect 11333 5865 11345 5868
rect 11379 5865 11391 5899
rect 11333 5859 11391 5865
rect 7377 5831 7435 5837
rect 7377 5797 7389 5831
rect 7423 5828 7435 5831
rect 8478 5828 8484 5840
rect 7423 5800 8484 5828
rect 7423 5797 7435 5800
rect 7377 5791 7435 5797
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 8846 5828 8852 5840
rect 8807 5800 8852 5828
rect 8846 5788 8852 5800
rect 8904 5788 8910 5840
rect 10137 5831 10195 5837
rect 10137 5828 10149 5831
rect 9692 5800 10149 5828
rect 9692 5772 9720 5800
rect 10137 5797 10149 5800
rect 10183 5797 10195 5831
rect 10137 5791 10195 5797
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5760 2191 5763
rect 3050 5760 3056 5772
rect 2179 5732 3056 5760
rect 2179 5729 2191 5732
rect 2133 5723 2191 5729
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 5074 5760 5080 5772
rect 5035 5732 5080 5760
rect 5074 5720 5080 5732
rect 5132 5720 5138 5772
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5760 6423 5763
rect 6638 5760 6644 5772
rect 6411 5732 6644 5760
rect 6411 5729 6423 5732
rect 6365 5723 6423 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 9674 5720 9680 5772
rect 9732 5720 9738 5772
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5692 4675 5695
rect 5166 5692 5172 5704
rect 4663 5664 5172 5692
rect 4663 5661 4675 5664
rect 4617 5655 4675 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 5276 5568 5304 5655
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7926 5692 7932 5704
rect 6972 5664 7932 5692
rect 6972 5652 6978 5664
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 6549 5627 6607 5633
rect 6549 5624 6561 5627
rect 5552 5596 6561 5624
rect 1762 5516 1768 5568
rect 1820 5556 1826 5568
rect 2317 5559 2375 5565
rect 2317 5556 2329 5559
rect 1820 5528 2329 5556
rect 1820 5516 1826 5528
rect 2317 5525 2329 5528
rect 2363 5525 2375 5559
rect 3418 5556 3424 5568
rect 3379 5528 3424 5556
rect 2317 5519 2375 5525
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4709 5559 4767 5565
rect 4709 5556 4721 5559
rect 4120 5528 4721 5556
rect 4120 5516 4126 5528
rect 4709 5525 4721 5528
rect 4755 5525 4767 5559
rect 4709 5519 4767 5525
rect 5258 5516 5264 5568
rect 5316 5516 5322 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 5552 5556 5580 5596
rect 6549 5593 6561 5596
rect 6595 5593 6607 5627
rect 7466 5624 7472 5636
rect 7427 5596 7472 5624
rect 6549 5587 6607 5593
rect 7466 5584 7472 5596
rect 7524 5584 7530 5636
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 8444 5596 9413 5624
rect 8444 5584 8450 5596
rect 9401 5593 9413 5596
rect 9447 5624 9459 5627
rect 10060 5624 10088 5723
rect 11514 5720 11520 5772
rect 11572 5760 11578 5772
rect 11701 5763 11759 5769
rect 11701 5760 11713 5763
rect 11572 5732 11713 5760
rect 11572 5720 11578 5732
rect 11701 5729 11713 5732
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 10229 5655 10287 5661
rect 10244 5624 10272 5655
rect 11146 5652 11152 5704
rect 11204 5692 11210 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11204 5664 11805 5692
rect 11204 5652 11210 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11974 5692 11980 5704
rect 11935 5664 11980 5692
rect 11793 5655 11851 5661
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 9447 5596 10088 5624
rect 10152 5596 10272 5624
rect 9447 5593 9459 5596
rect 9401 5587 9459 5593
rect 5902 5556 5908 5568
rect 5500 5528 5580 5556
rect 5863 5528 5908 5556
rect 5500 5516 5506 5528
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 7009 5559 7067 5565
rect 7009 5525 7021 5559
rect 7055 5556 7067 5559
rect 7098 5556 7104 5568
rect 7055 5528 7104 5556
rect 7055 5525 7067 5528
rect 7009 5519 7067 5525
rect 7098 5516 7104 5528
rect 7156 5556 7162 5568
rect 8110 5556 8116 5568
rect 7156 5528 8116 5556
rect 7156 5516 7162 5528
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8573 5559 8631 5565
rect 8573 5525 8585 5559
rect 8619 5556 8631 5559
rect 8662 5556 8668 5568
rect 8619 5528 8668 5556
rect 8619 5525 8631 5528
rect 8573 5519 8631 5525
rect 8662 5516 8668 5528
rect 8720 5556 8726 5568
rect 8846 5556 8852 5568
rect 8720 5528 8852 5556
rect 8720 5516 8726 5528
rect 8846 5516 8852 5528
rect 8904 5556 8910 5568
rect 10152 5556 10180 5596
rect 8904 5528 10180 5556
rect 8904 5516 8910 5528
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 4798 5352 4804 5364
rect 4759 5324 4804 5352
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5258 5352 5264 5364
rect 5215 5324 5264 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5537 5355 5595 5361
rect 5537 5321 5549 5355
rect 5583 5352 5595 5355
rect 5626 5352 5632 5364
rect 5583 5324 5632 5352
rect 5583 5321 5595 5324
rect 5537 5315 5595 5321
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 6638 5352 6644 5364
rect 6503 5324 6644 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 8168 5324 8585 5352
rect 8168 5312 8174 5324
rect 8573 5321 8585 5324
rect 8619 5352 8631 5355
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 8619 5324 10425 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 12032 5324 12173 5352
rect 12032 5312 12038 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 12161 5315 12219 5321
rect 2961 5287 3019 5293
rect 2961 5253 2973 5287
rect 3007 5284 3019 5287
rect 3050 5284 3056 5296
rect 3007 5256 3056 5284
rect 3007 5253 3019 5256
rect 2961 5247 3019 5253
rect 3050 5244 3056 5256
rect 3108 5244 3114 5296
rect 11054 5244 11060 5296
rect 11112 5284 11118 5296
rect 11425 5287 11483 5293
rect 11425 5284 11437 5287
rect 11112 5256 11437 5284
rect 11112 5244 11118 5256
rect 11425 5253 11437 5256
rect 11471 5253 11483 5287
rect 11425 5247 11483 5253
rect 2314 5216 2320 5228
rect 2275 5188 2320 5216
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5148 2099 5151
rect 2133 5151 2191 5157
rect 2133 5148 2145 5151
rect 2087 5120 2145 5148
rect 2087 5117 2099 5120
rect 2041 5111 2099 5117
rect 2133 5117 2145 5120
rect 2179 5148 2191 5151
rect 2406 5148 2412 5160
rect 2179 5120 2412 5148
rect 2179 5117 2191 5120
rect 2133 5111 2191 5117
rect 2406 5108 2412 5120
rect 2464 5108 2470 5160
rect 3418 5148 3424 5160
rect 3379 5120 3424 5148
rect 3418 5108 3424 5120
rect 3476 5108 3482 5160
rect 5626 5148 5632 5160
rect 5587 5120 5632 5148
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 5960 5120 6837 5148
rect 5960 5108 5966 5120
rect 6825 5117 6837 5120
rect 6871 5148 6883 5151
rect 6914 5148 6920 5160
rect 6871 5120 6920 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7098 5157 7104 5160
rect 7092 5148 7104 5157
rect 7059 5120 7104 5148
rect 7092 5111 7104 5120
rect 7098 5108 7104 5111
rect 7156 5108 7162 5160
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5148 9091 5151
rect 11241 5151 11299 5157
rect 9079 5120 9536 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 9508 5092 9536 5120
rect 11241 5117 11253 5151
rect 11287 5148 11299 5151
rect 11606 5148 11612 5160
rect 11287 5120 11612 5148
rect 11287 5117 11299 5120
rect 11241 5111 11299 5117
rect 11606 5108 11612 5120
rect 11664 5148 11670 5160
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 11664 5120 11805 5148
rect 11664 5108 11670 5120
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 3329 5083 3387 5089
rect 3329 5049 3341 5083
rect 3375 5080 3387 5083
rect 3688 5083 3746 5089
rect 3688 5080 3700 5083
rect 3375 5052 3700 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 3688 5049 3700 5052
rect 3734 5080 3746 5083
rect 3970 5080 3976 5092
rect 3734 5052 3976 5080
rect 3734 5049 3746 5052
rect 3688 5043 3746 5049
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 9278 5083 9336 5089
rect 9278 5080 9290 5083
rect 8864 5052 9290 5080
rect 8864 5024 8892 5052
rect 9278 5049 9290 5052
rect 9324 5049 9336 5083
rect 9278 5043 9336 5049
rect 9490 5040 9496 5092
rect 9548 5040 9554 5092
rect 10781 5083 10839 5089
rect 10781 5049 10793 5083
rect 10827 5080 10839 5083
rect 11514 5080 11520 5092
rect 10827 5052 11520 5080
rect 10827 5049 10839 5052
rect 10781 5043 10839 5049
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 5813 5015 5871 5021
rect 5813 5012 5825 5015
rect 5684 4984 5825 5012
rect 5684 4972 5690 4984
rect 5813 4981 5825 4984
rect 5859 4981 5871 5015
rect 5813 4975 5871 4981
rect 6638 4972 6644 5024
rect 6696 5012 6702 5024
rect 7098 5012 7104 5024
rect 6696 4984 7104 5012
rect 6696 4972 6702 4984
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 8202 5012 8208 5024
rect 8163 4984 8208 5012
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 8846 5012 8852 5024
rect 8807 4984 8852 5012
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 11146 5012 11152 5024
rect 11107 4984 11152 5012
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 12710 5012 12716 5024
rect 12483 4984 12716 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 2777 4811 2835 4817
rect 2777 4808 2789 4811
rect 2608 4780 2789 4808
rect 1949 4743 2007 4749
rect 1949 4709 1961 4743
rect 1995 4740 2007 4743
rect 2314 4740 2320 4752
rect 1995 4712 2320 4740
rect 1995 4709 2007 4712
rect 1949 4703 2007 4709
rect 2314 4700 2320 4712
rect 2372 4740 2378 4752
rect 2608 4740 2636 4780
rect 2777 4777 2789 4780
rect 2823 4777 2835 4811
rect 2777 4771 2835 4777
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 5997 4811 6055 4817
rect 5997 4808 6009 4811
rect 5316 4780 6009 4808
rect 5316 4768 5322 4780
rect 5997 4777 6009 4780
rect 6043 4777 6055 4811
rect 5997 4771 6055 4777
rect 6365 4811 6423 4817
rect 6365 4777 6377 4811
rect 6411 4808 6423 4811
rect 6822 4808 6828 4820
rect 6411 4780 6828 4808
rect 6411 4777 6423 4780
rect 6365 4771 6423 4777
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 8570 4808 8576 4820
rect 8531 4780 8576 4808
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 9953 4811 10011 4817
rect 9953 4808 9965 4811
rect 9824 4780 9965 4808
rect 9824 4768 9830 4780
rect 9953 4777 9965 4780
rect 9999 4808 10011 4811
rect 10226 4808 10232 4820
rect 9999 4780 10232 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 11793 4811 11851 4817
rect 11793 4808 11805 4811
rect 11572 4780 11805 4808
rect 11572 4768 11578 4780
rect 11793 4777 11805 4780
rect 11839 4777 11851 4811
rect 11793 4771 11851 4777
rect 2869 4743 2927 4749
rect 2869 4740 2881 4743
rect 2372 4712 2636 4740
rect 2792 4712 2881 4740
rect 2372 4700 2378 4712
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2792 4604 2820 4712
rect 2869 4709 2881 4712
rect 2915 4740 2927 4743
rect 4062 4740 4068 4752
rect 2915 4712 4068 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 6638 4700 6644 4752
rect 6696 4740 6702 4752
rect 6733 4743 6791 4749
rect 6733 4740 6745 4743
rect 6696 4712 6745 4740
rect 6696 4700 6702 4712
rect 6733 4709 6745 4712
rect 6779 4740 6791 4743
rect 7092 4743 7150 4749
rect 7092 4740 7104 4743
rect 6779 4712 7104 4740
rect 6779 4709 6791 4712
rect 6733 4703 6791 4709
rect 7092 4709 7104 4712
rect 7138 4740 7150 4743
rect 7374 4740 7380 4752
rect 7138 4712 7380 4740
rect 7138 4709 7150 4712
rect 7092 4703 7150 4709
rect 7374 4700 7380 4712
rect 7432 4740 7438 4752
rect 8202 4740 8208 4752
rect 7432 4712 8208 4740
rect 7432 4700 7438 4712
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 11701 4743 11759 4749
rect 11701 4709 11713 4743
rect 11747 4740 11759 4743
rect 12253 4743 12311 4749
rect 12253 4740 12265 4743
rect 11747 4712 12265 4740
rect 11747 4709 11759 4712
rect 11701 4703 11759 4709
rect 12253 4709 12265 4712
rect 12299 4740 12311 4743
rect 12434 4740 12440 4752
rect 12299 4712 12440 4740
rect 12299 4709 12311 4712
rect 12253 4703 12311 4709
rect 12434 4700 12440 4712
rect 12492 4700 12498 4752
rect 4522 4672 4528 4684
rect 4483 4644 4528 4672
rect 4522 4632 4528 4644
rect 4580 4672 4586 4684
rect 4873 4675 4931 4681
rect 4873 4672 4885 4675
rect 4580 4644 4885 4672
rect 4580 4632 4586 4644
rect 4873 4641 4885 4644
rect 4919 4641 4931 4675
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 4873 4635 4931 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 12158 4672 12164 4684
rect 11379 4644 12164 4672
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 12805 4675 12863 4681
rect 12805 4672 12817 4675
rect 12268 4644 12817 4672
rect 2363 4576 2820 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 2924 4576 3065 4604
rect 2924 4564 2930 4576
rect 3053 4573 3065 4576
rect 3099 4604 3111 4607
rect 3970 4604 3976 4616
rect 3099 4576 3976 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 6822 4604 6828 4616
rect 6783 4576 6828 4604
rect 4617 4567 4675 4573
rect 3878 4536 3884 4548
rect 3839 4508 3884 4536
rect 3878 4496 3884 4508
rect 3936 4496 3942 4548
rect 3418 4428 3424 4480
rect 3476 4468 3482 4480
rect 3513 4471 3571 4477
rect 3513 4468 3525 4471
rect 3476 4440 3525 4468
rect 3476 4428 3482 4440
rect 3513 4437 3525 4440
rect 3559 4468 3571 4471
rect 4632 4468 4660 4567
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 10686 4604 10692 4616
rect 10647 4576 10692 4604
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 8294 4496 8300 4548
rect 8352 4536 8358 4548
rect 9401 4539 9459 4545
rect 9401 4536 9413 4539
rect 8352 4508 9413 4536
rect 8352 4496 8358 4508
rect 9401 4505 9413 4508
rect 9447 4536 9459 4539
rect 9582 4536 9588 4548
rect 9447 4508 9588 4536
rect 9447 4505 9459 4508
rect 9401 4499 9459 4505
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 10229 4539 10287 4545
rect 10229 4505 10241 4539
rect 10275 4536 10287 4539
rect 12268 4536 12296 4644
rect 12805 4641 12817 4644
rect 12851 4672 12863 4675
rect 12894 4672 12900 4684
rect 12851 4644 12900 4672
rect 12851 4641 12863 4644
rect 12805 4635 12863 4641
rect 12894 4632 12900 4644
rect 12952 4632 12958 4684
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4604 12495 4607
rect 12618 4604 12624 4616
rect 12483 4576 12624 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 10275 4508 12296 4536
rect 10275 4505 10287 4508
rect 10229 4499 10287 4505
rect 5902 4468 5908 4480
rect 3559 4440 5908 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 6880 4440 8217 4468
rect 6880 4428 6886 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 8904 4440 9045 4468
rect 8904 4428 8910 4440
rect 9033 4437 9045 4440
rect 9079 4437 9091 4471
rect 9033 4431 9091 4437
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 12250 4468 12256 4480
rect 11388 4440 12256 4468
rect 11388 4428 11394 4440
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 2501 4267 2559 4273
rect 2501 4233 2513 4267
rect 2547 4264 2559 4267
rect 2866 4264 2872 4276
rect 2547 4236 2872 4264
rect 2547 4233 2559 4236
rect 2501 4227 2559 4233
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 3326 4264 3332 4276
rect 2976 4236 3332 4264
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 2976 4137 3004 4236
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 3970 4224 3976 4276
rect 4028 4264 4034 4276
rect 4341 4267 4399 4273
rect 4341 4264 4353 4267
rect 4028 4236 4353 4264
rect 4028 4224 4034 4236
rect 4341 4233 4353 4236
rect 4387 4233 4399 4267
rect 5166 4264 5172 4276
rect 5127 4236 5172 4264
rect 4341 4227 4399 4233
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 6178 4264 6184 4276
rect 6139 4236 6184 4264
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 6457 4267 6515 4273
rect 6457 4233 6469 4267
rect 6503 4264 6515 4267
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 6503 4236 6837 4264
rect 6503 4233 6515 4236
rect 6457 4227 6515 4233
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 8386 4264 8392 4276
rect 8347 4236 8392 4264
rect 6825 4227 6883 4233
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 10965 4267 11023 4273
rect 10965 4264 10977 4267
rect 10928 4236 10977 4264
rect 10928 4224 10934 4236
rect 10965 4233 10977 4236
rect 11011 4233 11023 4267
rect 10965 4227 11023 4233
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 12437 4267 12495 4273
rect 12437 4264 12449 4267
rect 11204 4236 12449 4264
rect 11204 4224 11210 4236
rect 12437 4233 12449 4236
rect 12483 4233 12495 4267
rect 12437 4227 12495 4233
rect 5258 4196 5264 4208
rect 4080 4168 5264 4196
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1486 4060 1492 4072
rect 1443 4032 1492 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1486 4020 1492 4032
rect 1544 4020 1550 4072
rect 3228 4063 3286 4069
rect 3228 4060 3240 4063
rect 3160 4032 3240 4060
rect 2869 3995 2927 4001
rect 2869 3961 2881 3995
rect 2915 3992 2927 3995
rect 3050 3992 3056 4004
rect 2915 3964 3056 3992
rect 2915 3961 2927 3964
rect 2869 3955 2927 3961
rect 3050 3952 3056 3964
rect 3108 3992 3114 4004
rect 3160 3992 3188 4032
rect 3228 4029 3240 4032
rect 3274 4060 3286 4063
rect 4080 4060 4108 4168
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 7190 4196 7196 4208
rect 6564 4168 7196 4196
rect 4522 4088 4528 4140
rect 4580 4128 4586 4140
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4580 4100 4721 4128
rect 4580 4088 4586 4100
rect 4709 4097 4721 4100
rect 4755 4128 4767 4131
rect 5810 4128 5816 4140
rect 4755 4100 5816 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 3274 4032 4108 4060
rect 5077 4063 5135 4069
rect 3274 4029 3286 4032
rect 3228 4023 3286 4029
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5123 4032 5549 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5537 4029 5549 4032
rect 5583 4060 5595 4063
rect 6564 4060 6592 4168
rect 7190 4156 7196 4168
rect 7248 4156 7254 4208
rect 7374 4156 7380 4208
rect 7432 4196 7438 4208
rect 7432 4168 7512 4196
rect 7432 4156 7438 4168
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7282 4128 7288 4140
rect 6972 4100 7288 4128
rect 6972 4088 6978 4100
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7484 4137 7512 4168
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 11793 4199 11851 4205
rect 11793 4196 11805 4199
rect 11296 4168 11805 4196
rect 11296 4156 11302 4168
rect 11793 4165 11805 4168
rect 11839 4196 11851 4199
rect 12161 4199 12219 4205
rect 12161 4196 12173 4199
rect 11839 4168 12173 4196
rect 11839 4165 11851 4168
rect 11793 4159 11851 4165
rect 12161 4165 12173 4168
rect 12207 4196 12219 4199
rect 12342 4196 12348 4208
rect 12207 4168 12348 4196
rect 12207 4165 12219 4168
rect 12161 4159 12219 4165
rect 12342 4156 12348 4168
rect 12400 4196 12406 4208
rect 12618 4196 12624 4208
rect 12400 4168 12624 4196
rect 12400 4156 12406 4168
rect 12618 4156 12624 4168
rect 12676 4196 12682 4208
rect 12676 4168 13032 4196
rect 12676 4156 12682 4168
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 8570 4128 8576 4140
rect 7708 4100 8576 4128
rect 7708 4088 7714 4100
rect 8570 4088 8576 4100
rect 8628 4128 8634 4140
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8628 4100 8953 4128
rect 8628 4088 8634 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9824 4100 9873 4128
rect 9824 4088 9830 4100
rect 9861 4097 9873 4100
rect 9907 4128 9919 4131
rect 10318 4128 10324 4140
rect 9907 4100 10324 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 10318 4088 10324 4100
rect 10376 4128 10382 4140
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 10376 4100 10425 4128
rect 10376 4088 10382 4100
rect 10413 4097 10425 4100
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 12894 4128 12900 4140
rect 10560 4100 10605 4128
rect 12855 4100 12900 4128
rect 10560 4088 10566 4100
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13004 4137 13032 4168
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 5583 4032 6592 4060
rect 6641 4063 6699 4069
rect 5583 4029 5595 4032
rect 5537 4023 5595 4029
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 8297 4063 8355 4069
rect 6687 4032 7420 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 3108 3964 3188 3992
rect 3108 3952 3114 3964
rect 4522 3952 4528 4004
rect 4580 3992 4586 4004
rect 5442 3992 5448 4004
rect 4580 3964 5448 3992
rect 4580 3952 4586 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 6457 3995 6515 4001
rect 6457 3992 6469 3995
rect 5644 3964 6469 3992
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 5644 3933 5672 3964
rect 6457 3961 6469 3964
rect 6503 3961 6515 3995
rect 6457 3955 6515 3961
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 5040 3896 5641 3924
rect 5040 3884 5046 3896
rect 5629 3893 5641 3896
rect 5675 3893 5687 3927
rect 5629 3887 5687 3893
rect 6178 3884 6184 3936
rect 6236 3924 6242 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 6236 3896 7205 3924
rect 6236 3884 6242 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 7193 3887 7251 3893
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7392 3924 7420 4032
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 8343 4032 8861 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8849 4029 8861 4032
rect 8895 4060 8907 4063
rect 9306 4060 9312 4072
rect 8895 4032 9312 4060
rect 8895 4029 8907 4032
rect 8849 4023 8907 4029
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 10042 4060 10048 4072
rect 9407 4032 10048 4060
rect 7929 3995 7987 4001
rect 7929 3961 7941 3995
rect 7975 3992 7987 3995
rect 8754 3992 8760 4004
rect 7975 3964 8760 3992
rect 7975 3961 7987 3964
rect 7929 3955 7987 3961
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 9407 3992 9435 4032
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 11054 3992 11060 4004
rect 9232 3964 9435 3992
rect 9968 3964 11060 3992
rect 7340 3896 7420 3924
rect 7340 3884 7346 3896
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 9232 3924 9260 3964
rect 8444 3896 9260 3924
rect 8444 3884 8450 3896
rect 9306 3884 9312 3936
rect 9364 3924 9370 3936
rect 9968 3933 9996 3964
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 12676 3964 12817 3992
rect 12676 3952 12682 3964
rect 12805 3961 12817 3964
rect 12851 3992 12863 3995
rect 13449 3995 13507 4001
rect 13449 3992 13461 3995
rect 12851 3964 13461 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 13449 3961 13461 3964
rect 13495 3961 13507 3995
rect 13449 3955 13507 3961
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 9364 3896 9413 3924
rect 9364 3884 9370 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 9401 3887 9459 3893
rect 9953 3927 10011 3933
rect 9953 3893 9965 3927
rect 9999 3893 10011 3927
rect 9953 3887 10011 3893
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10284 3896 10333 3924
rect 10284 3884 10290 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 11330 3924 11336 3936
rect 11291 3896 11336 3924
rect 10321 3887 10379 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 13354 3924 13360 3936
rect 13044 3896 13360 3924
rect 13044 3884 13050 3896
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 1486 3680 1492 3732
rect 1544 3720 1550 3732
rect 1581 3723 1639 3729
rect 1581 3720 1593 3723
rect 1544 3692 1593 3720
rect 1544 3680 1550 3692
rect 1581 3689 1593 3692
rect 1627 3689 1639 3723
rect 1581 3683 1639 3689
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 2409 3723 2467 3729
rect 2409 3720 2421 3723
rect 2372 3692 2421 3720
rect 2372 3680 2378 3692
rect 2409 3689 2421 3692
rect 2455 3689 2467 3723
rect 3418 3720 3424 3732
rect 3379 3692 3424 3720
rect 2409 3683 2467 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4982 3720 4988 3732
rect 3927 3692 4988 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5169 3723 5227 3729
rect 5169 3720 5181 3723
rect 5132 3692 5181 3720
rect 5132 3680 5138 3692
rect 5169 3689 5181 3692
rect 5215 3689 5227 3723
rect 6638 3720 6644 3732
rect 6599 3692 6644 3720
rect 5169 3683 5227 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7561 3723 7619 3729
rect 7561 3689 7573 3723
rect 7607 3720 7619 3723
rect 7650 3720 7656 3732
rect 7607 3692 7656 3720
rect 7607 3689 7619 3692
rect 7561 3683 7619 3689
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 8018 3720 8024 3732
rect 7979 3692 8024 3720
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8386 3720 8392 3732
rect 8347 3692 8392 3720
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8536 3692 9045 3720
rect 8536 3680 8542 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9033 3683 9091 3689
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3720 9919 3723
rect 10594 3720 10600 3732
rect 9907 3692 10600 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 10594 3680 10600 3692
rect 10652 3720 10658 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10652 3692 10885 3720
rect 10652 3680 10658 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 10873 3683 10931 3689
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11146 3720 11152 3732
rect 11020 3692 11152 3720
rect 11020 3680 11026 3692
rect 11146 3680 11152 3692
rect 11204 3720 11210 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 11204 3692 11253 3720
rect 11204 3680 11210 3692
rect 11241 3689 11253 3692
rect 11287 3689 11299 3723
rect 11241 3683 11299 3689
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 6273 3655 6331 3661
rect 2832 3624 2877 3652
rect 2832 3612 2838 3624
rect 6273 3621 6285 3655
rect 6319 3652 6331 3655
rect 6822 3652 6828 3664
rect 6319 3624 6828 3652
rect 6319 3621 6331 3624
rect 6273 3615 6331 3621
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3200 3556 4077 3584
rect 3200 3544 3206 3556
rect 4065 3553 4077 3556
rect 4111 3584 4123 3587
rect 4338 3584 4344 3596
rect 4111 3556 4344 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 4338 3544 4344 3556
rect 4396 3584 4402 3596
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4396 3556 4629 3584
rect 4396 3544 4402 3556
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3584 5595 3587
rect 5994 3584 6000 3596
rect 5583 3556 6000 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 6288 3528 6316 3615
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 9674 3612 9680 3664
rect 9732 3652 9738 3664
rect 10321 3655 10379 3661
rect 10321 3652 10333 3655
rect 9732 3624 10333 3652
rect 9732 3612 9738 3624
rect 10321 3621 10333 3624
rect 10367 3621 10379 3655
rect 11256 3652 11284 3683
rect 12342 3680 12348 3732
rect 12400 3720 12406 3732
rect 12805 3723 12863 3729
rect 12805 3720 12817 3723
rect 12400 3692 12817 3720
rect 12400 3680 12406 3692
rect 12805 3689 12817 3692
rect 12851 3689 12863 3723
rect 12805 3683 12863 3689
rect 11670 3655 11728 3661
rect 11670 3652 11682 3655
rect 11256 3624 11682 3652
rect 10321 3615 10379 3621
rect 11670 3621 11682 3624
rect 11716 3621 11728 3655
rect 11670 3615 11728 3621
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 6914 3584 6920 3596
rect 6779 3556 6920 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3516 2375 3519
rect 2682 3516 2688 3528
rect 2363 3488 2688 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3516 2872 3528
rect 2827 3488 2872 3516
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3050 3516 3056 3528
rect 3011 3488 3056 3516
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3485 5687 3519
rect 5810 3516 5816 3528
rect 5723 3488 5816 3516
rect 5629 3479 5687 3485
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 3068 3448 3096 3476
rect 2004 3420 3096 3448
rect 2004 3408 2010 3420
rect 4430 3408 4436 3460
rect 4488 3448 4494 3460
rect 5644 3448 5672 3479
rect 5810 3476 5816 3488
rect 5868 3516 5874 3528
rect 6270 3516 6276 3528
rect 5868 3488 6276 3516
rect 5868 3476 5874 3488
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 6748 3448 6776 3547
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 9950 3584 9956 3596
rect 8496 3556 9956 3584
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8496 3525 8524 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10226 3584 10232 3596
rect 10187 3556 10232 3584
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 8168 3488 8493 3516
rect 8168 3476 8174 3488
rect 8481 3485 8493 3488
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 10502 3516 10508 3528
rect 10459 3488 10508 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 8588 3448 8616 3479
rect 9306 3448 9312 3460
rect 4488 3420 6776 3448
rect 7852 3420 9312 3448
rect 4488 3408 4494 3420
rect 198 3340 204 3392
rect 256 3380 262 3392
rect 1302 3380 1308 3392
rect 256 3352 1308 3380
rect 256 3340 262 3352
rect 1302 3340 1308 3352
rect 1360 3340 1366 3392
rect 2406 3340 2412 3392
rect 2464 3380 2470 3392
rect 3418 3380 3424 3392
rect 2464 3352 3424 3380
rect 2464 3340 2470 3352
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 4246 3380 4252 3392
rect 4207 3352 4252 3380
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4982 3380 4988 3392
rect 4943 3352 4988 3380
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 6914 3380 6920 3392
rect 6875 3352 6920 3380
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 7852 3389 7880 3420
rect 9306 3408 9312 3420
rect 9364 3448 9370 3460
rect 10428 3448 10456 3479
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 9364 3420 10456 3448
rect 9364 3408 9370 3420
rect 7837 3383 7895 3389
rect 7837 3380 7849 3383
rect 7248 3352 7849 3380
rect 7248 3340 7254 3352
rect 7837 3349 7849 3352
rect 7883 3349 7895 3383
rect 9490 3380 9496 3392
rect 9451 3352 9496 3380
rect 7837 3343 7895 3349
rect 9490 3340 9496 3352
rect 9548 3380 9554 3392
rect 11440 3380 11468 3479
rect 13081 3383 13139 3389
rect 13081 3380 13093 3383
rect 9548 3352 13093 3380
rect 9548 3340 9554 3352
rect 13081 3349 13093 3352
rect 13127 3349 13139 3383
rect 13081 3343 13139 3349
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 1946 3176 1952 3188
rect 1907 3148 1952 3176
rect 1946 3136 1952 3148
rect 2004 3136 2010 3188
rect 2774 3136 2780 3188
rect 2832 3176 2838 3188
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 2832 3148 4905 3176
rect 2832 3136 2838 3148
rect 4893 3145 4905 3148
rect 4939 3145 4951 3179
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 4893 3139 4951 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 7009 3179 7067 3185
rect 7009 3176 7021 3179
rect 6880 3148 7021 3176
rect 6880 3136 6886 3148
rect 7009 3145 7021 3148
rect 7055 3145 7067 3179
rect 7834 3176 7840 3188
rect 7009 3139 7067 3145
rect 7208 3148 7840 3176
rect 4430 3108 4436 3120
rect 4391 3080 4436 3108
rect 4430 3068 4436 3080
rect 4488 3068 4494 3120
rect 4706 3108 4712 3120
rect 4667 3080 4712 3108
rect 4706 3068 4712 3080
rect 4764 3108 4770 3120
rect 5994 3108 6000 3120
rect 4764 3080 5396 3108
rect 5907 3080 6000 3108
rect 4764 3068 4770 3080
rect 5368 3049 5396 3080
rect 5994 3068 6000 3080
rect 6052 3108 6058 3120
rect 7208 3108 7236 3148
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 8941 3179 8999 3185
rect 8941 3176 8953 3179
rect 8904 3148 8953 3176
rect 8904 3136 8910 3148
rect 8941 3145 8953 3148
rect 8987 3145 8999 3179
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 8941 3139 8999 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 11146 3176 11152 3188
rect 11107 3148 11152 3176
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 12434 3176 12440 3188
rect 12395 3148 12440 3176
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 6052 3080 7236 3108
rect 6052 3068 6058 3080
rect 8570 3068 8576 3120
rect 8628 3108 8634 3120
rect 9398 3108 9404 3120
rect 8628 3080 9404 3108
rect 8628 3068 8634 3080
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3040 1455 3043
rect 5353 3043 5411 3049
rect 1443 3012 2544 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 2406 2972 2412 2984
rect 1728 2944 2412 2972
rect 1728 2932 1734 2944
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 2516 2972 2544 3012
rect 5353 3009 5365 3043
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 5810 3040 5816 3052
rect 5583 3012 5816 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 9217 3043 9275 3049
rect 9217 3040 9229 3043
rect 8588 3012 9229 3040
rect 4982 2972 4988 2984
rect 2516 2944 4988 2972
rect 4982 2932 4988 2944
rect 5040 2972 5046 2984
rect 5261 2975 5319 2981
rect 5261 2972 5273 2975
rect 5040 2944 5273 2972
rect 5040 2932 5046 2944
rect 5261 2941 5273 2944
rect 5307 2941 5319 2975
rect 5261 2935 5319 2941
rect 7466 2932 7472 2984
rect 7524 2972 7530 2984
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7524 2944 7573 2972
rect 7524 2932 7530 2944
rect 7561 2941 7573 2944
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 7817 2975 7875 2981
rect 7817 2972 7829 2975
rect 7708 2944 7829 2972
rect 7708 2932 7714 2944
rect 7817 2941 7829 2944
rect 7863 2941 7875 2975
rect 7817 2935 7875 2941
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 8588 2972 8616 3012
rect 9217 3009 9229 3012
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 11204 3012 13093 3040
rect 11204 3000 11210 3012
rect 13081 3009 13093 3012
rect 13127 3040 13139 3043
rect 13170 3040 13176 3052
rect 13127 3012 13176 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13170 3000 13176 3012
rect 13228 3040 13234 3052
rect 13449 3043 13507 3049
rect 13449 3040 13461 3043
rect 13228 3012 13461 3040
rect 13228 3000 13234 3012
rect 13449 3009 13461 3012
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 9490 2972 9496 2984
rect 8444 2944 8616 2972
rect 9232 2944 9496 2972
rect 8444 2932 8450 2944
rect 2222 2904 2228 2916
rect 2183 2876 2228 2904
rect 2222 2864 2228 2876
rect 2280 2904 2286 2916
rect 2654 2907 2712 2913
rect 2654 2904 2666 2907
rect 2280 2876 2666 2904
rect 2280 2864 2286 2876
rect 2654 2873 2666 2876
rect 2700 2873 2712 2907
rect 2654 2867 2712 2873
rect 7282 2864 7288 2916
rect 7340 2904 7346 2916
rect 7377 2907 7435 2913
rect 7377 2904 7389 2907
rect 7340 2876 7389 2904
rect 7340 2864 7346 2876
rect 7377 2873 7389 2876
rect 7423 2904 7435 2907
rect 8110 2904 8116 2916
rect 7423 2876 8116 2904
rect 7423 2873 7435 2876
rect 7377 2867 7435 2873
rect 8110 2864 8116 2876
rect 8168 2864 8174 2916
rect 3789 2839 3847 2845
rect 3789 2805 3801 2839
rect 3835 2836 3847 2839
rect 7190 2836 7196 2848
rect 3835 2808 7196 2836
rect 3835 2805 3847 2808
rect 3789 2799 3847 2805
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 9232 2836 9260 2944
rect 9490 2932 9496 2944
rect 9548 2972 9554 2984
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 9548 2944 9781 2972
rect 9548 2932 9554 2944
rect 9769 2941 9781 2944
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 11885 2975 11943 2981
rect 11885 2941 11897 2975
rect 11931 2972 11943 2975
rect 12526 2972 12532 2984
rect 11931 2944 12532 2972
rect 11931 2941 11943 2944
rect 11885 2935 11943 2941
rect 12526 2932 12532 2944
rect 12584 2972 12590 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12584 2944 12909 2972
rect 12584 2932 12590 2944
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 9306 2864 9312 2916
rect 9364 2904 9370 2916
rect 9582 2904 9588 2916
rect 9364 2876 9588 2904
rect 9364 2864 9370 2876
rect 9582 2864 9588 2876
rect 9640 2904 9646 2916
rect 10014 2907 10072 2913
rect 10014 2904 10026 2907
rect 9640 2876 10026 2904
rect 9640 2864 9646 2876
rect 10014 2873 10026 2876
rect 10060 2904 10072 2907
rect 11425 2907 11483 2913
rect 11425 2904 11437 2907
rect 10060 2876 11437 2904
rect 10060 2873 10072 2876
rect 10014 2867 10072 2873
rect 11425 2873 11437 2876
rect 11471 2873 11483 2907
rect 11425 2867 11483 2873
rect 12805 2907 12863 2913
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 13078 2904 13084 2916
rect 12851 2876 13084 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 7524 2808 9260 2836
rect 12253 2839 12311 2845
rect 7524 2796 7530 2808
rect 12253 2805 12265 2839
rect 12299 2836 12311 2839
rect 12820 2836 12848 2867
rect 13078 2864 13084 2876
rect 13136 2864 13142 2916
rect 12299 2808 12848 2836
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 1670 2632 1676 2644
rect 1631 2604 1676 2632
rect 1670 2592 1676 2604
rect 1728 2592 1734 2644
rect 2406 2632 2412 2644
rect 2367 2604 2412 2632
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 2866 2632 2872 2644
rect 2792 2604 2872 2632
rect 1765 2499 1823 2505
rect 1765 2465 1777 2499
rect 1811 2496 1823 2499
rect 2424 2496 2452 2592
rect 1811 2468 2452 2496
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 2792 2437 2820 2604
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 4338 2632 4344 2644
rect 4299 2604 4344 2632
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 4614 2632 4620 2644
rect 4575 2604 4620 2632
rect 4614 2592 4620 2604
rect 4672 2632 4678 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 4672 2604 5181 2632
rect 4672 2592 4678 2604
rect 5169 2601 5181 2604
rect 5215 2601 5227 2635
rect 5810 2632 5816 2644
rect 5771 2604 5816 2632
rect 5169 2595 5227 2601
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 7156 2604 7573 2632
rect 7156 2592 7162 2604
rect 7561 2601 7573 2604
rect 7607 2632 7619 2635
rect 8113 2635 8171 2641
rect 7607 2604 7972 2632
rect 7607 2601 7619 2604
rect 7561 2595 7619 2601
rect 3878 2564 3884 2576
rect 3839 2536 3884 2564
rect 3878 2524 3884 2536
rect 3936 2524 3942 2576
rect 4356 2564 4384 2592
rect 5261 2567 5319 2573
rect 5261 2564 5273 2567
rect 4356 2536 5273 2564
rect 5261 2533 5273 2536
rect 5307 2533 5319 2567
rect 5261 2527 5319 2533
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 2958 2496 2964 2508
rect 2915 2468 2964 2496
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 2958 2456 2964 2468
rect 3016 2496 3022 2508
rect 3421 2499 3479 2505
rect 3421 2496 3433 2499
rect 3016 2468 3433 2496
rect 3016 2456 3022 2468
rect 3421 2465 3433 2468
rect 3467 2465 3479 2499
rect 3421 2459 3479 2465
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6779 2468 6929 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 6917 2465 6929 2468
rect 6963 2496 6975 2499
rect 7558 2496 7564 2508
rect 6963 2468 7564 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7558 2456 7564 2468
rect 7616 2456 7622 2508
rect 7944 2496 7972 2604
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 8202 2632 8208 2644
rect 8159 2604 8208 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10045 2635 10103 2641
rect 10045 2601 10057 2635
rect 10091 2632 10103 2635
rect 10226 2632 10232 2644
rect 10091 2604 10232 2632
rect 10091 2601 10103 2604
rect 10045 2595 10103 2601
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10686 2632 10692 2644
rect 10647 2604 10692 2632
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 11112 2604 11161 2632
rect 11112 2592 11118 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 11149 2595 11207 2601
rect 12069 2635 12127 2641
rect 12069 2601 12081 2635
rect 12115 2632 12127 2635
rect 12710 2632 12716 2644
rect 12115 2604 12716 2632
rect 12115 2601 12127 2604
rect 12069 2595 12127 2601
rect 8021 2567 8079 2573
rect 8021 2533 8033 2567
rect 8067 2564 8079 2567
rect 8496 2564 8524 2592
rect 8067 2536 8524 2564
rect 11164 2564 11192 2595
rect 12710 2592 12716 2604
rect 12768 2632 12774 2644
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 12768 2604 13001 2632
rect 12768 2592 12774 2604
rect 12989 2601 13001 2604
rect 13035 2601 13047 2635
rect 12989 2595 13047 2601
rect 13078 2592 13084 2644
rect 13136 2632 13142 2644
rect 13446 2632 13452 2644
rect 13136 2604 13452 2632
rect 13136 2592 13142 2604
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 14001 2567 14059 2573
rect 14001 2564 14013 2567
rect 11164 2536 14013 2564
rect 8067 2533 8079 2536
rect 8021 2527 8079 2533
rect 14001 2533 14013 2536
rect 14047 2533 14059 2567
rect 14001 2527 14059 2533
rect 8573 2499 8631 2505
rect 8573 2496 8585 2499
rect 7944 2468 8585 2496
rect 8573 2465 8585 2468
rect 8619 2465 8631 2499
rect 8573 2459 8631 2465
rect 10410 2456 10416 2508
rect 10468 2496 10474 2508
rect 10597 2499 10655 2505
rect 10597 2496 10609 2499
rect 10468 2468 10609 2496
rect 10468 2456 10474 2468
rect 10597 2465 10609 2468
rect 10643 2496 10655 2499
rect 11057 2499 11115 2505
rect 11057 2496 11069 2499
rect 10643 2468 11069 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 11057 2465 11069 2468
rect 11103 2496 11115 2499
rect 12066 2496 12072 2508
rect 11103 2468 12072 2496
rect 11103 2465 11115 2468
rect 11057 2459 11115 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12437 2499 12495 2505
rect 12437 2465 12449 2499
rect 12483 2496 12495 2499
rect 13078 2496 13084 2508
rect 12483 2468 13084 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 13078 2456 13084 2468
rect 13136 2456 13142 2508
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 5445 2431 5503 2437
rect 2823 2400 4844 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 1949 2363 2007 2369
rect 1949 2329 1961 2363
rect 1995 2360 2007 2363
rect 2958 2360 2964 2372
rect 1995 2332 2964 2360
rect 1995 2329 2007 2332
rect 1949 2323 2007 2329
rect 2958 2320 2964 2332
rect 3016 2320 3022 2372
rect 4816 2369 4844 2400
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5810 2428 5816 2440
rect 5491 2400 5816 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 7650 2428 7656 2440
rect 6411 2400 7656 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 7650 2388 7656 2400
rect 7708 2428 7714 2440
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 7708 2400 8677 2428
rect 7708 2388 7714 2400
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 11146 2428 11152 2440
rect 9263 2400 11152 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 11146 2388 11152 2400
rect 11204 2428 11210 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 11204 2400 11253 2428
rect 11204 2388 11210 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13228 2400 13645 2428
rect 13228 2388 13234 2400
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 4801 2363 4859 2369
rect 4801 2329 4813 2363
rect 4847 2329 4859 2363
rect 4801 2323 4859 2329
rect 12158 2320 12164 2372
rect 12216 2360 12222 2372
rect 12621 2363 12679 2369
rect 12621 2360 12633 2363
rect 12216 2332 12633 2360
rect 12216 2320 12222 2332
rect 12621 2329 12633 2332
rect 12667 2329 12679 2363
rect 12621 2323 12679 2329
rect 3053 2295 3111 2301
rect 3053 2261 3065 2295
rect 3099 2292 3111 2295
rect 3326 2292 3332 2304
rect 3099 2264 3332 2292
rect 3099 2261 3111 2264
rect 3053 2255 3111 2261
rect 3326 2252 3332 2264
rect 3384 2252 3390 2304
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 3786 1980 3792 2032
rect 3844 2020 3850 2032
rect 5626 2020 5632 2032
rect 3844 1992 5632 2020
rect 3844 1980 3850 1992
rect 5626 1980 5632 1992
rect 5684 1980 5690 2032
rect 11790 1368 11796 1420
rect 11848 1408 11854 1420
rect 12250 1408 12256 1420
rect 11848 1380 12256 1408
rect 11848 1368 11854 1380
rect 12250 1368 12256 1380
rect 12308 1368 12314 1420
rect 9398 552 9404 604
rect 9456 592 9462 604
rect 9490 592 9496 604
rect 9456 564 9496 592
rect 9456 552 9462 564
rect 9490 552 9496 564
rect 9548 552 9554 604
<< via1 >>
rect 11336 37816 11388 37868
rect 12256 37816 12308 37868
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 13912 37136 13964 37188
rect 14556 37136 14608 37188
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 7288 36363 7340 36372
rect 7288 36329 7297 36363
rect 7297 36329 7331 36363
rect 7331 36329 7340 36363
rect 7288 36320 7340 36329
rect 7196 36184 7248 36236
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 4988 35776 5040 35828
rect 6920 35776 6972 35828
rect 7288 35572 7340 35624
rect 6000 35436 6052 35488
rect 7196 35436 7248 35488
rect 8208 35436 8260 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 3332 35232 3384 35284
rect 4252 35275 4304 35284
rect 4252 35241 4261 35275
rect 4261 35241 4295 35275
rect 4295 35241 4304 35275
rect 4252 35232 4304 35241
rect 5448 35232 5500 35284
rect 6644 35232 6696 35284
rect 7380 35232 7432 35284
rect 3056 35096 3108 35148
rect 4252 35096 4304 35148
rect 5172 35139 5224 35148
rect 5172 35105 5181 35139
rect 5181 35105 5215 35139
rect 5215 35105 5224 35139
rect 5172 35096 5224 35105
rect 6828 35096 6880 35148
rect 7472 35139 7524 35148
rect 7472 35105 7481 35139
rect 7481 35105 7515 35139
rect 7515 35105 7524 35139
rect 7472 35096 7524 35105
rect 11152 35096 11204 35148
rect 7288 34892 7340 34944
rect 8116 34935 8168 34944
rect 8116 34901 8125 34935
rect 8125 34901 8159 34935
rect 8159 34901 8168 34935
rect 8116 34892 8168 34901
rect 10048 34935 10100 34944
rect 10048 34901 10057 34935
rect 10057 34901 10091 34935
rect 10091 34901 10100 34935
rect 10048 34892 10100 34901
rect 12532 34892 12584 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 572 34688 624 34740
rect 2964 34688 3016 34740
rect 4252 34731 4304 34740
rect 4252 34697 4261 34731
rect 4261 34697 4295 34731
rect 4295 34697 4304 34731
rect 4252 34688 4304 34697
rect 6184 34688 6236 34740
rect 7472 34731 7524 34740
rect 7472 34697 7481 34731
rect 7481 34697 7515 34731
rect 7515 34697 7524 34731
rect 7472 34688 7524 34697
rect 8208 34688 8260 34740
rect 13636 34731 13688 34740
rect 13636 34697 13645 34731
rect 13645 34697 13679 34731
rect 13679 34697 13688 34731
rect 13636 34688 13688 34697
rect 204 34620 256 34672
rect 1308 34620 1360 34672
rect 1400 34620 1452 34672
rect 3056 34552 3108 34604
rect 2044 34527 2096 34536
rect 2044 34493 2053 34527
rect 2053 34493 2087 34527
rect 2087 34493 2096 34527
rect 2044 34484 2096 34493
rect 3332 34552 3384 34604
rect 3240 34484 3292 34536
rect 4804 34484 4856 34536
rect 5172 34527 5224 34536
rect 5172 34493 5181 34527
rect 5181 34493 5215 34527
rect 5215 34493 5224 34527
rect 5172 34484 5224 34493
rect 5724 34484 5776 34536
rect 6828 34484 6880 34536
rect 7840 34527 7892 34536
rect 7840 34493 7849 34527
rect 7849 34493 7883 34527
rect 7883 34493 7892 34527
rect 7840 34484 7892 34493
rect 8116 34527 8168 34536
rect 8116 34493 8150 34527
rect 8150 34493 8168 34527
rect 8116 34484 8168 34493
rect 11060 34620 11112 34672
rect 10048 34527 10100 34536
rect 8024 34416 8076 34468
rect 10048 34493 10057 34527
rect 10057 34493 10091 34527
rect 10091 34493 10100 34527
rect 10048 34484 10100 34493
rect 13452 34527 13504 34536
rect 13452 34493 13461 34527
rect 13461 34493 13495 34527
rect 13495 34493 13504 34527
rect 13452 34484 13504 34493
rect 12072 34348 12124 34400
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 940 34144 992 34196
rect 1768 34144 1820 34196
rect 4160 34144 4212 34196
rect 5540 34144 5592 34196
rect 7748 34187 7800 34196
rect 7748 34153 7757 34187
rect 7757 34153 7791 34187
rect 7791 34153 7800 34187
rect 7748 34144 7800 34153
rect 2412 34008 2464 34060
rect 3148 34008 3200 34060
rect 4252 34008 4304 34060
rect 6092 34008 6144 34060
rect 7840 34008 7892 34060
rect 9680 34008 9732 34060
rect 10048 34144 10100 34196
rect 11152 34187 11204 34196
rect 11152 34153 11161 34187
rect 11161 34153 11195 34187
rect 11195 34153 11204 34187
rect 11152 34144 11204 34153
rect 11244 34144 11296 34196
rect 10048 34051 10100 34060
rect 10048 34017 10082 34051
rect 10082 34017 10100 34051
rect 10048 34008 10100 34017
rect 12072 34076 12124 34128
rect 11152 34008 11204 34060
rect 13452 34008 13504 34060
rect 12532 33983 12584 33992
rect 12532 33949 12541 33983
rect 12541 33949 12575 33983
rect 12575 33949 12584 33983
rect 12532 33940 12584 33949
rect 10784 33872 10836 33924
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 1400 33600 1452 33652
rect 2136 33600 2188 33652
rect 7380 33643 7432 33652
rect 7380 33609 7389 33643
rect 7389 33609 7423 33643
rect 7423 33609 7432 33643
rect 7380 33600 7432 33609
rect 7840 33600 7892 33652
rect 8576 33600 8628 33652
rect 9312 33643 9364 33652
rect 9312 33609 9321 33643
rect 9321 33609 9355 33643
rect 9355 33609 9364 33643
rect 9312 33600 9364 33609
rect 10048 33464 10100 33516
rect 10968 33600 11020 33652
rect 11244 33600 11296 33652
rect 13452 33643 13504 33652
rect 13452 33609 13461 33643
rect 13461 33609 13495 33643
rect 13495 33609 13504 33643
rect 13452 33600 13504 33609
rect 12072 33464 12124 33516
rect 2688 33396 2740 33448
rect 7748 33439 7800 33448
rect 7748 33405 7757 33439
rect 7757 33405 7791 33439
rect 7791 33405 7800 33439
rect 7748 33396 7800 33405
rect 3148 33371 3200 33380
rect 3148 33337 3157 33371
rect 3157 33337 3191 33371
rect 3191 33337 3200 33371
rect 3148 33328 3200 33337
rect 4712 33328 4764 33380
rect 9312 33328 9364 33380
rect 12348 33396 12400 33448
rect 12164 33371 12216 33380
rect 12164 33337 12173 33371
rect 12173 33337 12207 33371
rect 12207 33337 12216 33371
rect 12900 33371 12952 33380
rect 12164 33328 12216 33337
rect 12900 33337 12909 33371
rect 12909 33337 12943 33371
rect 12943 33337 12952 33371
rect 12900 33328 12952 33337
rect 2044 33303 2096 33312
rect 2044 33269 2053 33303
rect 2053 33269 2087 33303
rect 2087 33269 2096 33303
rect 2044 33260 2096 33269
rect 2412 33303 2464 33312
rect 2412 33269 2421 33303
rect 2421 33269 2455 33303
rect 2455 33269 2464 33303
rect 2412 33260 2464 33269
rect 4252 33303 4304 33312
rect 4252 33269 4261 33303
rect 4261 33269 4295 33303
rect 4295 33269 4304 33303
rect 4252 33260 4304 33269
rect 5172 33303 5224 33312
rect 5172 33269 5181 33303
rect 5181 33269 5215 33303
rect 5215 33269 5224 33303
rect 5172 33260 5224 33269
rect 6092 33260 6144 33312
rect 9496 33303 9548 33312
rect 9496 33269 9505 33303
rect 9505 33269 9539 33303
rect 9539 33269 9548 33303
rect 9496 33260 9548 33269
rect 11428 33303 11480 33312
rect 11428 33269 11437 33303
rect 11437 33269 11471 33303
rect 11471 33269 11480 33303
rect 11428 33260 11480 33269
rect 12072 33260 12124 33312
rect 12440 33303 12492 33312
rect 12440 33269 12449 33303
rect 12449 33269 12483 33303
rect 12483 33269 12492 33303
rect 12808 33303 12860 33312
rect 12440 33260 12492 33269
rect 12808 33269 12817 33303
rect 12817 33269 12851 33303
rect 12851 33269 12860 33303
rect 12808 33260 12860 33269
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 5172 33056 5224 33108
rect 9496 33056 9548 33108
rect 10876 33056 10928 33108
rect 12808 33056 12860 33108
rect 1492 32988 1544 33040
rect 11612 32988 11664 33040
rect 1768 32920 1820 32972
rect 6920 32963 6972 32972
rect 6920 32929 6954 32963
rect 6954 32929 6972 32963
rect 6920 32920 6972 32929
rect 9680 32920 9732 32972
rect 10048 32920 10100 32972
rect 5540 32895 5592 32904
rect 5540 32861 5549 32895
rect 5549 32861 5583 32895
rect 5583 32861 5592 32895
rect 5540 32852 5592 32861
rect 6644 32895 6696 32904
rect 2688 32716 2740 32768
rect 5448 32716 5500 32768
rect 6644 32861 6653 32895
rect 6653 32861 6687 32895
rect 6687 32861 6696 32895
rect 6644 32852 6696 32861
rect 11060 32852 11112 32904
rect 11980 32895 12032 32904
rect 11244 32784 11296 32836
rect 11980 32861 11989 32895
rect 11989 32861 12023 32895
rect 12023 32861 12032 32895
rect 11980 32852 12032 32861
rect 12072 32895 12124 32904
rect 12072 32861 12081 32895
rect 12081 32861 12115 32895
rect 12115 32861 12124 32895
rect 12072 32852 12124 32861
rect 7012 32716 7064 32768
rect 9312 32716 9364 32768
rect 11520 32759 11572 32768
rect 11520 32725 11529 32759
rect 11529 32725 11563 32759
rect 11563 32725 11572 32759
rect 11520 32716 11572 32725
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 4988 32555 5040 32564
rect 4988 32521 4997 32555
rect 4997 32521 5031 32555
rect 5031 32521 5040 32555
rect 4988 32512 5040 32521
rect 5172 32555 5224 32564
rect 5172 32521 5181 32555
rect 5181 32521 5215 32555
rect 5215 32521 5224 32555
rect 5172 32512 5224 32521
rect 6184 32512 6236 32564
rect 6552 32555 6604 32564
rect 6552 32521 6561 32555
rect 6561 32521 6595 32555
rect 6595 32521 6604 32555
rect 6552 32512 6604 32521
rect 8300 32512 8352 32564
rect 10048 32555 10100 32564
rect 10048 32521 10057 32555
rect 10057 32521 10091 32555
rect 10091 32521 10100 32555
rect 10048 32512 10100 32521
rect 10324 32555 10376 32564
rect 10324 32521 10333 32555
rect 10333 32521 10367 32555
rect 10367 32521 10376 32555
rect 10324 32512 10376 32521
rect 10968 32512 11020 32564
rect 11612 32555 11664 32564
rect 11612 32521 11621 32555
rect 11621 32521 11655 32555
rect 11655 32521 11664 32555
rect 11612 32512 11664 32521
rect 11980 32555 12032 32564
rect 11980 32521 11989 32555
rect 11989 32521 12023 32555
rect 12023 32521 12032 32555
rect 11980 32512 12032 32521
rect 5540 32444 5592 32496
rect 6920 32444 6972 32496
rect 5908 32308 5960 32360
rect 8576 32376 8628 32428
rect 11060 32419 11112 32428
rect 11060 32385 11069 32419
rect 11069 32385 11103 32419
rect 11103 32385 11112 32419
rect 11060 32376 11112 32385
rect 12808 32376 12860 32428
rect 6920 32308 6972 32360
rect 7932 32308 7984 32360
rect 9312 32351 9364 32360
rect 9312 32317 9321 32351
rect 9321 32317 9355 32351
rect 9355 32317 9364 32351
rect 9312 32308 9364 32317
rect 10324 32308 10376 32360
rect 6552 32240 6604 32292
rect 6736 32240 6788 32292
rect 8668 32240 8720 32292
rect 1768 32172 1820 32224
rect 5632 32172 5684 32224
rect 7380 32172 7432 32224
rect 8852 32215 8904 32224
rect 8852 32181 8861 32215
rect 8861 32181 8895 32215
rect 8895 32181 8904 32215
rect 8852 32172 8904 32181
rect 10968 32215 11020 32224
rect 10968 32181 10977 32215
rect 10977 32181 11011 32215
rect 11011 32181 11020 32215
rect 10968 32172 11020 32181
rect 11980 32172 12032 32224
rect 12624 32172 12676 32224
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 5540 31968 5592 32020
rect 5908 31968 5960 32020
rect 6920 32011 6972 32020
rect 1676 31943 1728 31952
rect 1676 31909 1685 31943
rect 1685 31909 1719 31943
rect 1719 31909 1728 31943
rect 1676 31900 1728 31909
rect 5632 31900 5684 31952
rect 6920 31977 6929 32011
rect 6929 31977 6963 32011
rect 6963 31977 6972 32011
rect 6920 31968 6972 31977
rect 8300 31968 8352 32020
rect 9496 32011 9548 32020
rect 9496 31977 9505 32011
rect 9505 31977 9539 32011
rect 9539 31977 9548 32011
rect 9496 31968 9548 31977
rect 11060 31968 11112 32020
rect 11520 32011 11572 32020
rect 11520 31977 11529 32011
rect 11529 31977 11563 32011
rect 11563 31977 11572 32011
rect 11520 31968 11572 31977
rect 7196 31943 7248 31952
rect 7196 31909 7205 31943
rect 7205 31909 7239 31943
rect 7239 31909 7248 31943
rect 7196 31900 7248 31909
rect 7472 31900 7524 31952
rect 8576 31900 8628 31952
rect 9588 31900 9640 31952
rect 10968 31900 11020 31952
rect 1676 31764 1728 31816
rect 3424 31628 3476 31680
rect 5172 31875 5224 31884
rect 5172 31841 5206 31875
rect 5206 31841 5224 31875
rect 5172 31832 5224 31841
rect 6552 31832 6604 31884
rect 7380 31875 7432 31884
rect 7380 31841 7389 31875
rect 7389 31841 7423 31875
rect 7423 31841 7432 31875
rect 7380 31832 7432 31841
rect 12348 31832 12400 31884
rect 9956 31764 10008 31816
rect 11428 31696 11480 31748
rect 14924 31764 14976 31816
rect 14740 31696 14792 31748
rect 10508 31628 10560 31680
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 5632 31424 5684 31476
rect 6552 31467 6604 31476
rect 6552 31433 6561 31467
rect 6561 31433 6595 31467
rect 6595 31433 6604 31467
rect 6552 31424 6604 31433
rect 7472 31424 7524 31476
rect 11520 31467 11572 31476
rect 11520 31433 11529 31467
rect 11529 31433 11563 31467
rect 11563 31433 11572 31467
rect 11520 31424 11572 31433
rect 12348 31424 12400 31476
rect 8024 31288 8076 31340
rect 11520 31288 11572 31340
rect 1676 31263 1728 31272
rect 1676 31229 1685 31263
rect 1685 31229 1719 31263
rect 1719 31229 1728 31263
rect 1676 31220 1728 31229
rect 3424 31220 3476 31272
rect 10508 31263 10560 31272
rect 10508 31229 10517 31263
rect 10517 31229 10551 31263
rect 10551 31229 10560 31263
rect 10508 31220 10560 31229
rect 10784 31220 10836 31272
rect 4344 31152 4396 31204
rect 8024 31195 8076 31204
rect 8024 31161 8033 31195
rect 8033 31161 8067 31195
rect 8067 31161 8076 31195
rect 8024 31152 8076 31161
rect 4160 31084 4212 31136
rect 5172 31084 5224 31136
rect 6920 31084 6972 31136
rect 8116 31127 8168 31136
rect 8116 31093 8125 31127
rect 8125 31093 8159 31127
rect 8159 31093 8168 31127
rect 8116 31084 8168 31093
rect 10140 31127 10192 31136
rect 10140 31093 10149 31127
rect 10149 31093 10183 31127
rect 10183 31093 10192 31127
rect 10140 31084 10192 31093
rect 11244 31127 11296 31136
rect 11244 31093 11253 31127
rect 11253 31093 11287 31127
rect 11287 31093 11296 31127
rect 11244 31084 11296 31093
rect 11428 31084 11480 31136
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 7288 30880 7340 30932
rect 8116 30923 8168 30932
rect 8116 30889 8125 30923
rect 8125 30889 8159 30923
rect 8159 30889 8168 30923
rect 8116 30880 8168 30889
rect 10784 30880 10836 30932
rect 11520 30880 11572 30932
rect 11244 30812 11296 30864
rect 4436 30787 4488 30796
rect 4436 30753 4445 30787
rect 4445 30753 4479 30787
rect 4479 30753 4488 30787
rect 4436 30744 4488 30753
rect 4988 30744 5040 30796
rect 7104 30787 7156 30796
rect 7104 30753 7113 30787
rect 7113 30753 7147 30787
rect 7147 30753 7156 30787
rect 7104 30744 7156 30753
rect 7380 30744 7432 30796
rect 9680 30744 9732 30796
rect 10232 30744 10284 30796
rect 4344 30676 4396 30728
rect 5632 30719 5684 30728
rect 5632 30685 5641 30719
rect 5641 30685 5675 30719
rect 5675 30685 5684 30719
rect 5632 30676 5684 30685
rect 7196 30719 7248 30728
rect 7196 30685 7205 30719
rect 7205 30685 7239 30719
rect 7239 30685 7248 30719
rect 7196 30676 7248 30685
rect 2964 30583 3016 30592
rect 2964 30549 2973 30583
rect 2973 30549 3007 30583
rect 3007 30549 3016 30583
rect 2964 30540 3016 30549
rect 4068 30583 4120 30592
rect 4068 30549 4077 30583
rect 4077 30549 4111 30583
rect 4111 30549 4120 30583
rect 4068 30540 4120 30549
rect 5264 30540 5316 30592
rect 5540 30583 5592 30592
rect 5540 30549 5549 30583
rect 5549 30549 5583 30583
rect 5583 30549 5592 30583
rect 5540 30540 5592 30549
rect 6644 30583 6696 30592
rect 6644 30549 6653 30583
rect 6653 30549 6687 30583
rect 6687 30549 6696 30583
rect 6644 30540 6696 30549
rect 7840 30540 7892 30592
rect 8760 30540 8812 30592
rect 9312 30540 9364 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 2228 30311 2280 30320
rect 2228 30277 2237 30311
rect 2237 30277 2271 30311
rect 2271 30277 2280 30311
rect 2228 30268 2280 30277
rect 7196 30336 7248 30388
rect 8116 30336 8168 30388
rect 8576 30268 8628 30320
rect 9956 30311 10008 30320
rect 1584 30243 1636 30252
rect 1584 30209 1593 30243
rect 1593 30209 1627 30243
rect 1627 30209 1636 30243
rect 1584 30200 1636 30209
rect 5356 30200 5408 30252
rect 7104 30200 7156 30252
rect 7288 30200 7340 30252
rect 8208 30200 8260 30252
rect 8392 30200 8444 30252
rect 9956 30277 9965 30311
rect 9965 30277 9999 30311
rect 9999 30277 10008 30311
rect 9956 30268 10008 30277
rect 2964 30132 3016 30184
rect 3424 30132 3476 30184
rect 3516 30064 3568 30116
rect 5724 30064 5776 30116
rect 7748 30107 7800 30116
rect 7748 30073 7757 30107
rect 7757 30073 7791 30107
rect 7791 30073 7800 30107
rect 7748 30064 7800 30073
rect 4344 29996 4396 30048
rect 4896 30039 4948 30048
rect 4896 30005 4905 30039
rect 4905 30005 4939 30039
rect 4939 30005 4948 30039
rect 4896 29996 4948 30005
rect 4988 29996 5040 30048
rect 5264 29996 5316 30048
rect 7380 29996 7432 30048
rect 7840 30039 7892 30048
rect 7840 30005 7849 30039
rect 7849 30005 7883 30039
rect 7883 30005 7892 30039
rect 7840 29996 7892 30005
rect 9312 30132 9364 30184
rect 11244 30336 11296 30388
rect 10600 30200 10652 30252
rect 10140 29996 10192 30048
rect 10508 30039 10560 30048
rect 10508 30005 10517 30039
rect 10517 30005 10551 30039
rect 10551 30005 10560 30039
rect 10508 29996 10560 30005
rect 10968 30039 11020 30048
rect 10968 30005 10977 30039
rect 10977 30005 11011 30039
rect 11011 30005 11020 30039
rect 10968 29996 11020 30005
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 2780 29835 2832 29844
rect 2780 29801 2789 29835
rect 2789 29801 2823 29835
rect 2823 29801 2832 29835
rect 2780 29792 2832 29801
rect 4068 29792 4120 29844
rect 4436 29792 4488 29844
rect 5540 29792 5592 29844
rect 6644 29792 6696 29844
rect 7748 29835 7800 29844
rect 7748 29801 7757 29835
rect 7757 29801 7791 29835
rect 7791 29801 7800 29835
rect 7748 29792 7800 29801
rect 8024 29835 8076 29844
rect 8024 29801 8033 29835
rect 8033 29801 8067 29835
rect 8067 29801 8076 29835
rect 8024 29792 8076 29801
rect 8300 29792 8352 29844
rect 8852 29792 8904 29844
rect 10232 29835 10284 29844
rect 10232 29801 10241 29835
rect 10241 29801 10275 29835
rect 10275 29801 10284 29835
rect 10232 29792 10284 29801
rect 4988 29724 5040 29776
rect 5172 29724 5224 29776
rect 5632 29724 5684 29776
rect 8576 29724 8628 29776
rect 10508 29724 10560 29776
rect 2872 29699 2924 29708
rect 2872 29665 2881 29699
rect 2881 29665 2915 29699
rect 2915 29665 2924 29699
rect 2872 29656 2924 29665
rect 5448 29656 5500 29708
rect 6276 29656 6328 29708
rect 11244 29792 11296 29844
rect 10968 29724 11020 29776
rect 11520 29724 11572 29776
rect 2964 29631 3016 29640
rect 2964 29597 2973 29631
rect 2973 29597 3007 29631
rect 3007 29597 3016 29631
rect 2964 29588 3016 29597
rect 4160 29588 4212 29640
rect 5080 29588 5132 29640
rect 5632 29588 5684 29640
rect 7012 29588 7064 29640
rect 8208 29588 8260 29640
rect 10508 29588 10560 29640
rect 5448 29520 5500 29572
rect 8760 29520 8812 29572
rect 9588 29520 9640 29572
rect 1400 29452 1452 29504
rect 3516 29495 3568 29504
rect 3516 29461 3525 29495
rect 3525 29461 3559 29495
rect 3559 29461 3568 29495
rect 3516 29452 3568 29461
rect 4344 29495 4396 29504
rect 4344 29461 4353 29495
rect 4353 29461 4387 29495
rect 4387 29461 4396 29495
rect 4344 29452 4396 29461
rect 4620 29452 4672 29504
rect 5816 29495 5868 29504
rect 5816 29461 5825 29495
rect 5825 29461 5859 29495
rect 5859 29461 5868 29495
rect 5816 29452 5868 29461
rect 9496 29452 9548 29504
rect 11520 29452 11572 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 1584 29291 1636 29300
rect 1584 29257 1593 29291
rect 1593 29257 1627 29291
rect 1627 29257 1636 29291
rect 1584 29248 1636 29257
rect 2964 29248 3016 29300
rect 5080 29248 5132 29300
rect 7012 29291 7064 29300
rect 7012 29257 7021 29291
rect 7021 29257 7055 29291
rect 7055 29257 7064 29291
rect 7012 29248 7064 29257
rect 8208 29248 8260 29300
rect 10968 29291 11020 29300
rect 10968 29257 10977 29291
rect 10977 29257 11011 29291
rect 11011 29257 11020 29291
rect 10968 29248 11020 29257
rect 11244 29291 11296 29300
rect 11244 29257 11253 29291
rect 11253 29257 11287 29291
rect 11287 29257 11296 29291
rect 11244 29248 11296 29257
rect 4160 29180 4212 29232
rect 5356 29180 5408 29232
rect 9588 29180 9640 29232
rect 2044 29155 2096 29164
rect 2044 29121 2053 29155
rect 2053 29121 2087 29155
rect 2087 29121 2096 29155
rect 2044 29112 2096 29121
rect 3516 29112 3568 29164
rect 4344 29112 4396 29164
rect 5448 29112 5500 29164
rect 5632 29155 5684 29164
rect 5632 29121 5641 29155
rect 5641 29121 5675 29155
rect 5675 29121 5684 29155
rect 5632 29112 5684 29121
rect 5816 29155 5868 29164
rect 5816 29121 5825 29155
rect 5825 29121 5859 29155
rect 5859 29121 5868 29155
rect 5816 29112 5868 29121
rect 9496 29112 9548 29164
rect 5540 29087 5592 29096
rect 5540 29053 5549 29087
rect 5549 29053 5583 29087
rect 5583 29053 5592 29087
rect 5540 29044 5592 29053
rect 8852 29044 8904 29096
rect 3240 28976 3292 29028
rect 3976 28976 4028 29028
rect 6000 28976 6052 29028
rect 6276 29019 6328 29028
rect 6276 28985 6285 29019
rect 6285 28985 6319 29019
rect 6319 28985 6328 29019
rect 6276 28976 6328 28985
rect 8944 29019 8996 29028
rect 8944 28985 8953 29019
rect 8953 28985 8987 29019
rect 8987 28985 8996 29019
rect 8944 28976 8996 28985
rect 9680 28976 9732 29028
rect 10048 28976 10100 29028
rect 10324 28976 10376 29028
rect 10508 29019 10560 29028
rect 10508 28985 10517 29019
rect 10517 28985 10551 29019
rect 10551 28985 10560 29019
rect 10508 28976 10560 28985
rect 11980 28976 12032 29028
rect 12072 28976 12124 29028
rect 2872 28951 2924 28960
rect 2872 28917 2881 28951
rect 2881 28917 2915 28951
rect 2915 28917 2924 28951
rect 2872 28908 2924 28917
rect 3516 28908 3568 28960
rect 6920 28908 6972 28960
rect 7472 28908 7524 28960
rect 8392 28908 8444 28960
rect 9220 28908 9272 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 2780 28704 2832 28756
rect 2872 28704 2924 28756
rect 4160 28704 4212 28756
rect 5172 28747 5224 28756
rect 5172 28713 5181 28747
rect 5181 28713 5215 28747
rect 5215 28713 5224 28747
rect 5172 28704 5224 28713
rect 6644 28704 6696 28756
rect 7012 28747 7064 28756
rect 7012 28713 7021 28747
rect 7021 28713 7055 28747
rect 7055 28713 7064 28747
rect 7012 28704 7064 28713
rect 8208 28747 8260 28756
rect 8208 28713 8217 28747
rect 8217 28713 8251 28747
rect 8251 28713 8260 28747
rect 8208 28704 8260 28713
rect 8576 28747 8628 28756
rect 8576 28713 8585 28747
rect 8585 28713 8619 28747
rect 8619 28713 8628 28747
rect 8576 28704 8628 28713
rect 10232 28704 10284 28756
rect 3516 28679 3568 28688
rect 3516 28645 3525 28679
rect 3525 28645 3559 28679
rect 3559 28645 3568 28679
rect 3516 28636 3568 28645
rect 4988 28636 5040 28688
rect 7104 28636 7156 28688
rect 7472 28679 7524 28688
rect 7472 28645 7481 28679
rect 7481 28645 7515 28679
rect 7515 28645 7524 28679
rect 7472 28636 7524 28645
rect 5448 28568 5500 28620
rect 5724 28568 5776 28620
rect 5908 28611 5960 28620
rect 5908 28577 5917 28611
rect 5917 28577 5951 28611
rect 5951 28577 5960 28611
rect 5908 28568 5960 28577
rect 7564 28611 7616 28620
rect 7564 28577 7573 28611
rect 7573 28577 7607 28611
rect 7607 28577 7616 28611
rect 7564 28568 7616 28577
rect 4620 28543 4672 28552
rect 4620 28509 4629 28543
rect 4629 28509 4663 28543
rect 4663 28509 4672 28543
rect 4620 28500 4672 28509
rect 7012 28500 7064 28552
rect 7748 28500 7800 28552
rect 7932 28500 7984 28552
rect 9220 28500 9272 28552
rect 11060 28568 11112 28620
rect 9680 28500 9732 28552
rect 10784 28543 10836 28552
rect 10784 28509 10793 28543
rect 10793 28509 10827 28543
rect 10827 28509 10836 28543
rect 10784 28500 10836 28509
rect 11520 28500 11572 28552
rect 4528 28432 4580 28484
rect 5540 28432 5592 28484
rect 4068 28364 4120 28416
rect 5264 28364 5316 28416
rect 6920 28364 6972 28416
rect 8116 28364 8168 28416
rect 10324 28407 10376 28416
rect 10324 28373 10333 28407
rect 10333 28373 10367 28407
rect 10367 28373 10376 28407
rect 10324 28364 10376 28373
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 2044 28203 2096 28212
rect 2044 28169 2053 28203
rect 2053 28169 2087 28203
rect 2087 28169 2096 28203
rect 2044 28160 2096 28169
rect 3332 28160 3384 28212
rect 4620 28203 4672 28212
rect 2596 28092 2648 28144
rect 2044 27956 2096 28008
rect 4620 28169 4629 28203
rect 4629 28169 4663 28203
rect 4663 28169 4672 28203
rect 4620 28160 4672 28169
rect 6828 28160 6880 28212
rect 3700 28024 3752 28076
rect 4344 28024 4396 28076
rect 5632 28067 5684 28076
rect 5632 28033 5641 28067
rect 5641 28033 5675 28067
rect 5675 28033 5684 28067
rect 5632 28024 5684 28033
rect 5816 28067 5868 28076
rect 5816 28033 5825 28067
rect 5825 28033 5859 28067
rect 5859 28033 5868 28067
rect 5816 28024 5868 28033
rect 6736 28024 6788 28076
rect 5540 27999 5592 28008
rect 5540 27965 5549 27999
rect 5549 27965 5583 27999
rect 5583 27965 5592 27999
rect 5540 27956 5592 27965
rect 4068 27931 4120 27940
rect 4068 27897 4077 27931
rect 4077 27897 4111 27931
rect 4111 27897 4120 27931
rect 4068 27888 4120 27897
rect 7472 28160 7524 28212
rect 10600 28160 10652 28212
rect 10784 28203 10836 28212
rect 10784 28169 10793 28203
rect 10793 28169 10827 28203
rect 10827 28169 10836 28203
rect 10784 28160 10836 28169
rect 11060 28203 11112 28212
rect 11060 28169 11069 28203
rect 11069 28169 11103 28203
rect 11103 28169 11112 28203
rect 11060 28160 11112 28169
rect 11520 28203 11572 28212
rect 11520 28169 11529 28203
rect 11529 28169 11563 28203
rect 11563 28169 11572 28203
rect 11520 28160 11572 28169
rect 8116 28092 8168 28144
rect 8760 28092 8812 28144
rect 7472 28067 7524 28076
rect 7472 28033 7481 28067
rect 7481 28033 7515 28067
rect 7515 28033 7524 28067
rect 7472 28024 7524 28033
rect 7748 28024 7800 28076
rect 8208 27956 8260 28008
rect 8392 27956 8444 28008
rect 7564 27888 7616 27940
rect 10232 27956 10284 28008
rect 9496 27888 9548 27940
rect 4528 27820 4580 27872
rect 5448 27820 5500 27872
rect 8760 27863 8812 27872
rect 8760 27829 8769 27863
rect 8769 27829 8803 27863
rect 8803 27829 8812 27863
rect 8760 27820 8812 27829
rect 9220 27820 9272 27872
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 3700 27659 3752 27668
rect 3700 27625 3709 27659
rect 3709 27625 3743 27659
rect 3743 27625 3752 27659
rect 3700 27616 3752 27625
rect 4528 27616 4580 27668
rect 4160 27548 4212 27600
rect 5632 27616 5684 27668
rect 7104 27659 7156 27668
rect 7104 27625 7113 27659
rect 7113 27625 7147 27659
rect 7147 27625 7156 27659
rect 7104 27616 7156 27625
rect 7472 27616 7524 27668
rect 9496 27616 9548 27668
rect 10324 27616 10376 27668
rect 10784 27616 10836 27668
rect 11520 27548 11572 27600
rect 5264 27480 5316 27532
rect 6828 27480 6880 27532
rect 7196 27480 7248 27532
rect 9128 27480 9180 27532
rect 9772 27480 9824 27532
rect 4620 27276 4672 27328
rect 4896 27276 4948 27328
rect 6736 27276 6788 27328
rect 10232 27412 10284 27464
rect 11428 27412 11480 27464
rect 7564 27276 7616 27328
rect 9312 27276 9364 27328
rect 10692 27276 10744 27328
rect 12900 27319 12952 27328
rect 12900 27285 12909 27319
rect 12909 27285 12943 27319
rect 12943 27285 12952 27319
rect 12900 27276 12952 27285
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 3424 27115 3476 27124
rect 3424 27081 3433 27115
rect 3433 27081 3467 27115
rect 3467 27081 3476 27115
rect 3424 27072 3476 27081
rect 5264 27072 5316 27124
rect 5724 27072 5776 27124
rect 5908 27072 5960 27124
rect 6644 27072 6696 27124
rect 6828 27072 6880 27124
rect 11520 27115 11572 27124
rect 11520 27081 11529 27115
rect 11529 27081 11563 27115
rect 11563 27081 11572 27115
rect 11520 27072 11572 27081
rect 4160 26936 4212 26988
rect 6184 26936 6236 26988
rect 10784 26936 10836 26988
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 6000 26868 6052 26920
rect 6828 26868 6880 26920
rect 7472 26911 7524 26920
rect 7472 26877 7481 26911
rect 7481 26877 7515 26911
rect 7515 26877 7524 26911
rect 7472 26868 7524 26877
rect 12808 26868 12860 26920
rect 13360 26868 13412 26920
rect 4896 26800 4948 26852
rect 5816 26800 5868 26852
rect 6552 26800 6604 26852
rect 10692 26800 10744 26852
rect 7288 26775 7340 26784
rect 7288 26741 7297 26775
rect 7297 26741 7331 26775
rect 7331 26741 7340 26775
rect 7288 26732 7340 26741
rect 8760 26732 8812 26784
rect 9772 26732 9824 26784
rect 10048 26775 10100 26784
rect 10048 26741 10057 26775
rect 10057 26741 10091 26775
rect 10091 26741 10100 26775
rect 10048 26732 10100 26741
rect 10232 26732 10284 26784
rect 10416 26775 10468 26784
rect 10416 26741 10425 26775
rect 10425 26741 10459 26775
rect 10459 26741 10468 26775
rect 10416 26732 10468 26741
rect 11428 26732 11480 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 4068 26571 4120 26580
rect 4068 26537 4077 26571
rect 4077 26537 4111 26571
rect 4111 26537 4120 26571
rect 4068 26528 4120 26537
rect 5356 26528 5408 26580
rect 5632 26528 5684 26580
rect 9680 26528 9732 26580
rect 10692 26528 10744 26580
rect 1676 26503 1728 26512
rect 1676 26469 1685 26503
rect 1685 26469 1719 26503
rect 1719 26469 1728 26503
rect 1676 26460 1728 26469
rect 4528 26460 4580 26512
rect 6276 26460 6328 26512
rect 6736 26460 6788 26512
rect 10968 26460 11020 26512
rect 1492 26392 1544 26444
rect 7472 26392 7524 26444
rect 10048 26435 10100 26444
rect 10048 26401 10057 26435
rect 10057 26401 10091 26435
rect 10091 26401 10100 26435
rect 10048 26392 10100 26401
rect 4436 26324 4488 26376
rect 4896 26324 4948 26376
rect 5540 26324 5592 26376
rect 5908 26367 5960 26376
rect 5908 26333 5917 26367
rect 5917 26333 5951 26367
rect 5951 26333 5960 26367
rect 5908 26324 5960 26333
rect 9496 26324 9548 26376
rect 10600 26324 10652 26376
rect 7288 26299 7340 26308
rect 7288 26265 7297 26299
rect 7297 26265 7331 26299
rect 7331 26265 7340 26299
rect 7288 26256 7340 26265
rect 9680 26299 9732 26308
rect 9680 26265 9689 26299
rect 9689 26265 9723 26299
rect 9723 26265 9732 26299
rect 9680 26256 9732 26265
rect 7196 26188 7248 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 4436 25984 4488 26036
rect 6276 26027 6328 26036
rect 6276 25993 6285 26027
rect 6285 25993 6319 26027
rect 6319 25993 6328 26027
rect 6276 25984 6328 25993
rect 6644 26027 6696 26036
rect 6644 25993 6653 26027
rect 6653 25993 6687 26027
rect 6687 25993 6696 26027
rect 6644 25984 6696 25993
rect 7104 25984 7156 26036
rect 7288 25984 7340 26036
rect 7564 25984 7616 26036
rect 1492 25916 1544 25968
rect 9496 25916 9548 25968
rect 9680 25916 9732 25968
rect 10048 25916 10100 25968
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 5540 25848 5592 25900
rect 10232 25984 10284 26036
rect 5632 25823 5684 25832
rect 5632 25789 5641 25823
rect 5641 25789 5675 25823
rect 5675 25789 5684 25823
rect 5632 25780 5684 25789
rect 4528 25755 4580 25764
rect 4528 25721 4537 25755
rect 4537 25721 4571 25755
rect 4571 25721 4580 25755
rect 4528 25712 4580 25721
rect 5540 25755 5592 25764
rect 5540 25721 5549 25755
rect 5549 25721 5583 25755
rect 5583 25721 5592 25755
rect 5540 25712 5592 25721
rect 11520 25984 11572 26036
rect 10508 25780 10560 25832
rect 2504 25687 2556 25696
rect 2504 25653 2513 25687
rect 2513 25653 2547 25687
rect 2547 25653 2556 25687
rect 2504 25644 2556 25653
rect 4896 25687 4948 25696
rect 4896 25653 4905 25687
rect 4905 25653 4939 25687
rect 4939 25653 4948 25687
rect 4896 25644 4948 25653
rect 5080 25644 5132 25696
rect 5632 25644 5684 25696
rect 7656 25644 7708 25696
rect 9680 25687 9732 25696
rect 9680 25653 9689 25687
rect 9689 25653 9723 25687
rect 9723 25653 9732 25687
rect 9680 25644 9732 25653
rect 9864 25687 9916 25696
rect 9864 25653 9873 25687
rect 9873 25653 9907 25687
rect 9907 25653 9916 25687
rect 9864 25644 9916 25653
rect 10140 25687 10192 25696
rect 10140 25653 10149 25687
rect 10149 25653 10183 25687
rect 10183 25653 10192 25687
rect 10140 25644 10192 25653
rect 10600 25687 10652 25696
rect 10600 25653 10609 25687
rect 10609 25653 10643 25687
rect 10643 25653 10652 25687
rect 10600 25644 10652 25653
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 4896 25440 4948 25492
rect 5540 25440 5592 25492
rect 9588 25440 9640 25492
rect 10048 25372 10100 25424
rect 10600 25440 10652 25492
rect 12624 25483 12676 25492
rect 12624 25449 12633 25483
rect 12633 25449 12667 25483
rect 12667 25449 12676 25483
rect 12624 25440 12676 25449
rect 12900 25440 12952 25492
rect 1400 25347 1452 25356
rect 1400 25313 1409 25347
rect 1409 25313 1443 25347
rect 1443 25313 1452 25347
rect 1400 25304 1452 25313
rect 4160 25304 4212 25356
rect 6644 25304 6696 25356
rect 10600 25304 10652 25356
rect 12532 25347 12584 25356
rect 12532 25313 12541 25347
rect 12541 25313 12575 25347
rect 12575 25313 12584 25347
rect 12532 25304 12584 25313
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 4068 25279 4120 25288
rect 4068 25245 4077 25279
rect 4077 25245 4111 25279
rect 4111 25245 4120 25279
rect 4068 25236 4120 25245
rect 10048 25236 10100 25288
rect 10416 25236 10468 25288
rect 9496 25168 9548 25220
rect 10784 25168 10836 25220
rect 12900 25236 12952 25288
rect 5908 25100 5960 25152
rect 6736 25100 6788 25152
rect 7196 25143 7248 25152
rect 7196 25109 7205 25143
rect 7205 25109 7239 25143
rect 7239 25109 7248 25143
rect 7196 25100 7248 25109
rect 7472 25143 7524 25152
rect 7472 25109 7481 25143
rect 7481 25109 7515 25143
rect 7515 25109 7524 25143
rect 7472 25100 7524 25109
rect 9588 25100 9640 25152
rect 12348 25100 12400 25152
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 1400 24896 1452 24948
rect 6644 24896 6696 24948
rect 10600 24939 10652 24948
rect 10600 24905 10609 24939
rect 10609 24905 10643 24939
rect 10643 24905 10652 24939
rect 10600 24896 10652 24905
rect 12532 24896 12584 24948
rect 13176 24896 13228 24948
rect 7196 24828 7248 24880
rect 5908 24760 5960 24812
rect 12900 24828 12952 24880
rect 8300 24760 8352 24812
rect 9496 24803 9548 24812
rect 9496 24769 9505 24803
rect 9505 24769 9539 24803
rect 9539 24769 9548 24803
rect 9496 24760 9548 24769
rect 5264 24692 5316 24744
rect 5448 24692 5500 24744
rect 6920 24692 6972 24744
rect 7472 24735 7524 24744
rect 7472 24701 7481 24735
rect 7481 24701 7515 24735
rect 7515 24701 7524 24735
rect 7472 24692 7524 24701
rect 9312 24692 9364 24744
rect 10140 24760 10192 24812
rect 10232 24692 10284 24744
rect 10416 24735 10468 24744
rect 10416 24701 10425 24735
rect 10425 24701 10459 24735
rect 10459 24701 10468 24735
rect 10416 24692 10468 24701
rect 3148 24556 3200 24608
rect 4068 24624 4120 24676
rect 7012 24624 7064 24676
rect 4160 24599 4212 24608
rect 4160 24565 4169 24599
rect 4169 24565 4203 24599
rect 4203 24565 4212 24599
rect 4160 24556 4212 24565
rect 5080 24599 5132 24608
rect 5080 24565 5089 24599
rect 5089 24565 5123 24599
rect 5123 24565 5132 24599
rect 5080 24556 5132 24565
rect 5172 24556 5224 24608
rect 7104 24599 7156 24608
rect 7104 24565 7113 24599
rect 7113 24565 7147 24599
rect 7147 24565 7156 24599
rect 7104 24556 7156 24565
rect 9036 24599 9088 24608
rect 9036 24565 9045 24599
rect 9045 24565 9079 24599
rect 9079 24565 9088 24599
rect 9036 24556 9088 24565
rect 9588 24556 9640 24608
rect 9864 24556 9916 24608
rect 10784 24624 10836 24676
rect 10968 24692 11020 24744
rect 12164 24667 12216 24676
rect 12164 24633 12173 24667
rect 12173 24633 12207 24667
rect 12207 24633 12216 24667
rect 12164 24624 12216 24633
rect 11980 24556 12032 24608
rect 12624 24556 12676 24608
rect 12992 24556 13044 24608
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 5172 24395 5224 24404
rect 5172 24361 5181 24395
rect 5181 24361 5215 24395
rect 5215 24361 5224 24395
rect 5172 24352 5224 24361
rect 6000 24352 6052 24404
rect 8300 24395 8352 24404
rect 8300 24361 8309 24395
rect 8309 24361 8343 24395
rect 8343 24361 8352 24395
rect 8300 24352 8352 24361
rect 9496 24352 9548 24404
rect 10048 24352 10100 24404
rect 10140 24352 10192 24404
rect 10968 24352 11020 24404
rect 12716 24395 12768 24404
rect 12716 24361 12725 24395
rect 12725 24361 12759 24395
rect 12759 24361 12768 24395
rect 12716 24352 12768 24361
rect 6092 24216 6144 24268
rect 7196 24259 7248 24268
rect 7196 24225 7230 24259
rect 7230 24225 7248 24259
rect 7196 24216 7248 24225
rect 10692 24216 10744 24268
rect 12900 24352 12952 24404
rect 13176 24395 13228 24404
rect 13176 24361 13185 24395
rect 13185 24361 13219 24395
rect 13219 24361 13228 24395
rect 13176 24352 13228 24361
rect 13176 24216 13228 24268
rect 5908 24191 5960 24200
rect 5908 24157 5917 24191
rect 5917 24157 5951 24191
rect 5951 24157 5960 24191
rect 5908 24148 5960 24157
rect 3148 24055 3200 24064
rect 3148 24021 3157 24055
rect 3157 24021 3191 24055
rect 3191 24021 3200 24055
rect 3148 24012 3200 24021
rect 5356 24055 5408 24064
rect 5356 24021 5365 24055
rect 5365 24021 5399 24055
rect 5399 24021 5408 24055
rect 5356 24012 5408 24021
rect 6736 24012 6788 24064
rect 6920 24012 6972 24064
rect 8668 24055 8720 24064
rect 8668 24021 8677 24055
rect 8677 24021 8711 24055
rect 8711 24021 8720 24055
rect 8668 24012 8720 24021
rect 12348 24055 12400 24064
rect 12348 24021 12357 24055
rect 12357 24021 12391 24055
rect 12391 24021 12400 24055
rect 12348 24012 12400 24021
rect 12440 24012 12492 24064
rect 12716 24012 12768 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 4436 23808 4488 23860
rect 5908 23808 5960 23860
rect 7012 23851 7064 23860
rect 7012 23817 7021 23851
rect 7021 23817 7055 23851
rect 7055 23817 7064 23851
rect 7012 23808 7064 23817
rect 9864 23808 9916 23860
rect 11520 23851 11572 23860
rect 6000 23740 6052 23792
rect 5172 23672 5224 23724
rect 7932 23740 7984 23792
rect 3148 23604 3200 23656
rect 3884 23604 3936 23656
rect 5632 23604 5684 23656
rect 6000 23604 6052 23656
rect 6644 23647 6696 23656
rect 6644 23613 6653 23647
rect 6653 23613 6687 23647
rect 6687 23613 6696 23647
rect 6644 23604 6696 23613
rect 7196 23604 7248 23656
rect 8208 23672 8260 23724
rect 8668 23672 8720 23724
rect 9220 23715 9272 23724
rect 9220 23681 9229 23715
rect 9229 23681 9263 23715
rect 9263 23681 9272 23715
rect 9220 23672 9272 23681
rect 11520 23817 11529 23851
rect 11529 23817 11563 23851
rect 11563 23817 11572 23851
rect 11520 23808 11572 23817
rect 12532 23808 12584 23860
rect 12900 23740 12952 23792
rect 3516 23536 3568 23588
rect 6092 23536 6144 23588
rect 6920 23536 6972 23588
rect 8392 23604 8444 23656
rect 12440 23672 12492 23724
rect 13268 23672 13320 23724
rect 8024 23536 8076 23588
rect 9680 23579 9732 23588
rect 9680 23545 9689 23579
rect 9689 23545 9723 23579
rect 9723 23545 9732 23579
rect 9680 23536 9732 23545
rect 10692 23536 10744 23588
rect 12348 23536 12400 23588
rect 12624 23604 12676 23656
rect 12716 23536 12768 23588
rect 4160 23468 4212 23520
rect 4620 23468 4672 23520
rect 5172 23468 5224 23520
rect 12440 23511 12492 23520
rect 12440 23477 12449 23511
rect 12449 23477 12483 23511
rect 12483 23477 12492 23511
rect 12440 23468 12492 23477
rect 12624 23468 12676 23520
rect 13176 23468 13228 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 3056 23264 3108 23316
rect 4804 23264 4856 23316
rect 6828 23264 6880 23316
rect 7564 23307 7616 23316
rect 7564 23273 7573 23307
rect 7573 23273 7607 23307
rect 7607 23273 7616 23307
rect 7564 23264 7616 23273
rect 8024 23307 8076 23316
rect 8024 23273 8033 23307
rect 8033 23273 8067 23307
rect 8067 23273 8076 23307
rect 8024 23264 8076 23273
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 12256 23264 12308 23316
rect 12900 23264 12952 23316
rect 2780 23239 2832 23248
rect 2780 23205 2789 23239
rect 2789 23205 2823 23239
rect 2823 23205 2832 23239
rect 2780 23196 2832 23205
rect 4436 23239 4488 23248
rect 4436 23205 4470 23239
rect 4470 23205 4488 23239
rect 4436 23196 4488 23205
rect 7932 23239 7984 23248
rect 7932 23205 7941 23239
rect 7941 23205 7975 23239
rect 7975 23205 7984 23239
rect 7932 23196 7984 23205
rect 10692 23196 10744 23248
rect 11428 23196 11480 23248
rect 12532 23196 12584 23248
rect 2872 23171 2924 23180
rect 2872 23137 2881 23171
rect 2881 23137 2915 23171
rect 2915 23137 2924 23171
rect 3884 23171 3936 23180
rect 2872 23128 2924 23137
rect 3884 23137 3893 23171
rect 3893 23137 3927 23171
rect 3927 23137 3936 23171
rect 6828 23171 6880 23180
rect 3884 23128 3936 23137
rect 6828 23137 6837 23171
rect 6837 23137 6871 23171
rect 6871 23137 6880 23171
rect 6828 23128 6880 23137
rect 8208 23128 8260 23180
rect 10232 23128 10284 23180
rect 12440 23128 12492 23180
rect 2964 23103 3016 23112
rect 2964 23069 2973 23103
rect 2973 23069 3007 23103
rect 3007 23069 3016 23103
rect 2964 23060 3016 23069
rect 4068 23060 4120 23112
rect 4160 23103 4212 23112
rect 4160 23069 4169 23103
rect 4169 23069 4203 23103
rect 4203 23069 4212 23103
rect 4160 23060 4212 23069
rect 6184 23060 6236 23112
rect 6920 23103 6972 23112
rect 6920 23069 6929 23103
rect 6929 23069 6963 23103
rect 6963 23069 6972 23103
rect 6920 23060 6972 23069
rect 6644 22992 6696 23044
rect 7196 23060 7248 23112
rect 8760 23060 8812 23112
rect 9680 23103 9732 23112
rect 9680 23069 9689 23103
rect 9689 23069 9723 23103
rect 9723 23069 9732 23103
rect 9680 23060 9732 23069
rect 2412 22967 2464 22976
rect 2412 22933 2421 22967
rect 2421 22933 2455 22967
rect 2455 22933 2464 22967
rect 2412 22924 2464 22933
rect 4896 22924 4948 22976
rect 9680 22924 9732 22976
rect 9864 22924 9916 22976
rect 13452 22924 13504 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2872 22720 2924 22772
rect 5356 22763 5408 22772
rect 4436 22652 4488 22704
rect 1584 22627 1636 22636
rect 1584 22593 1593 22627
rect 1593 22593 1627 22627
rect 1627 22593 1636 22627
rect 1584 22584 1636 22593
rect 2964 22584 3016 22636
rect 1676 22516 1728 22568
rect 2412 22516 2464 22568
rect 3056 22516 3108 22568
rect 3240 22516 3292 22568
rect 3516 22584 3568 22636
rect 4344 22584 4396 22636
rect 5356 22729 5365 22763
rect 5365 22729 5399 22763
rect 5399 22729 5408 22763
rect 5356 22720 5408 22729
rect 6184 22763 6236 22772
rect 6184 22729 6193 22763
rect 6193 22729 6227 22763
rect 6227 22729 6236 22763
rect 6184 22720 6236 22729
rect 6644 22720 6696 22772
rect 8300 22720 8352 22772
rect 8668 22720 8720 22772
rect 10968 22720 11020 22772
rect 11428 22763 11480 22772
rect 11428 22729 11437 22763
rect 11437 22729 11471 22763
rect 11471 22729 11480 22763
rect 11428 22720 11480 22729
rect 12440 22720 12492 22772
rect 7196 22695 7248 22704
rect 7196 22661 7205 22695
rect 7205 22661 7239 22695
rect 7239 22661 7248 22695
rect 7196 22652 7248 22661
rect 12532 22652 12584 22704
rect 4896 22584 4948 22636
rect 10232 22627 10284 22636
rect 10232 22593 10241 22627
rect 10241 22593 10275 22627
rect 10275 22593 10284 22627
rect 10232 22584 10284 22593
rect 6828 22516 6880 22568
rect 7380 22559 7432 22568
rect 7380 22525 7389 22559
rect 7389 22525 7423 22559
rect 7423 22525 7432 22559
rect 7380 22516 7432 22525
rect 8024 22516 8076 22568
rect 4344 22448 4396 22500
rect 2964 22380 3016 22432
rect 3424 22380 3476 22432
rect 4988 22448 5040 22500
rect 7564 22448 7616 22500
rect 8300 22448 8352 22500
rect 8484 22448 8536 22500
rect 4620 22380 4672 22432
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 1676 22219 1728 22228
rect 1676 22185 1685 22219
rect 1685 22185 1719 22219
rect 1719 22185 1728 22219
rect 1676 22176 1728 22185
rect 2964 22176 3016 22228
rect 3240 22219 3292 22228
rect 3240 22185 3249 22219
rect 3249 22185 3283 22219
rect 3283 22185 3292 22219
rect 3240 22176 3292 22185
rect 4068 22176 4120 22228
rect 5080 22176 5132 22228
rect 2872 22108 2924 22160
rect 3516 22108 3568 22160
rect 4896 22108 4948 22160
rect 4436 21972 4488 22024
rect 6736 22108 6788 22160
rect 7380 22108 7432 22160
rect 5816 22040 5868 22092
rect 8760 22176 8812 22228
rect 11152 22176 11204 22228
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 11152 22040 11204 22092
rect 13452 22083 13504 22092
rect 13452 22049 13461 22083
rect 13461 22049 13495 22083
rect 13495 22049 13504 22083
rect 13452 22040 13504 22049
rect 5724 21972 5776 22024
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 9864 21972 9916 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 2780 21904 2832 21956
rect 13636 21947 13688 21956
rect 13636 21913 13645 21947
rect 13645 21913 13679 21947
rect 13679 21913 13688 21947
rect 13636 21904 13688 21913
rect 4620 21836 4672 21888
rect 4804 21836 4856 21888
rect 7104 21836 7156 21888
rect 8208 21836 8260 21888
rect 8484 21836 8536 21888
rect 9312 21836 9364 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 3516 21632 3568 21684
rect 4804 21675 4856 21684
rect 4804 21641 4813 21675
rect 4813 21641 4847 21675
rect 4847 21641 4856 21675
rect 4804 21632 4856 21641
rect 6920 21632 6972 21684
rect 8392 21632 8444 21684
rect 10048 21632 10100 21684
rect 4068 21564 4120 21616
rect 4344 21539 4396 21548
rect 4344 21505 4353 21539
rect 4353 21505 4387 21539
rect 4387 21505 4396 21539
rect 5448 21539 5500 21548
rect 4344 21496 4396 21505
rect 5448 21505 5457 21539
rect 5457 21505 5491 21539
rect 5491 21505 5500 21539
rect 5448 21496 5500 21505
rect 7564 21496 7616 21548
rect 9312 21539 9364 21548
rect 9312 21505 9321 21539
rect 9321 21505 9355 21539
rect 9355 21505 9364 21539
rect 9312 21496 9364 21505
rect 9496 21539 9548 21548
rect 9496 21505 9505 21539
rect 9505 21505 9539 21539
rect 9539 21505 9548 21539
rect 9496 21496 9548 21505
rect 5540 21428 5592 21480
rect 5908 21428 5960 21480
rect 7380 21428 7432 21480
rect 8116 21428 8168 21480
rect 5172 21403 5224 21412
rect 5172 21369 5181 21403
rect 5181 21369 5215 21403
rect 5215 21369 5224 21403
rect 5172 21360 5224 21369
rect 4620 21292 4672 21344
rect 5908 21335 5960 21344
rect 5908 21301 5917 21335
rect 5917 21301 5951 21335
rect 5951 21301 5960 21335
rect 5908 21292 5960 21301
rect 7748 21335 7800 21344
rect 7748 21301 7757 21335
rect 7757 21301 7791 21335
rect 7791 21301 7800 21335
rect 7748 21292 7800 21301
rect 8576 21292 8628 21344
rect 9864 21335 9916 21344
rect 9864 21301 9873 21335
rect 9873 21301 9907 21335
rect 9907 21301 9916 21335
rect 9864 21292 9916 21301
rect 12440 21292 12492 21344
rect 13452 21335 13504 21344
rect 13452 21301 13461 21335
rect 13461 21301 13495 21335
rect 13495 21301 13504 21335
rect 13452 21292 13504 21301
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 4436 21131 4488 21140
rect 4436 21097 4445 21131
rect 4445 21097 4479 21131
rect 4479 21097 4488 21131
rect 4436 21088 4488 21097
rect 6092 21131 6144 21140
rect 6092 21097 6101 21131
rect 6101 21097 6135 21131
rect 6135 21097 6144 21131
rect 6092 21088 6144 21097
rect 7380 21131 7432 21140
rect 7380 21097 7389 21131
rect 7389 21097 7423 21131
rect 7423 21097 7432 21131
rect 7380 21088 7432 21097
rect 7840 21088 7892 21140
rect 8208 21131 8260 21140
rect 8208 21097 8217 21131
rect 8217 21097 8251 21131
rect 8251 21097 8260 21131
rect 8208 21088 8260 21097
rect 8484 21088 8536 21140
rect 8944 21088 8996 21140
rect 10232 21088 10284 21140
rect 7564 21020 7616 21072
rect 6460 20995 6512 21004
rect 6460 20961 6469 20995
rect 6469 20961 6503 20995
rect 6503 20961 6512 20995
rect 6460 20952 6512 20961
rect 9496 21020 9548 21072
rect 10508 20995 10560 21004
rect 10508 20961 10542 20995
rect 10542 20961 10560 20995
rect 10508 20952 10560 20961
rect 5540 20884 5592 20936
rect 6092 20884 6144 20936
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 8116 20884 8168 20936
rect 8392 20927 8444 20936
rect 8392 20893 8401 20927
rect 8401 20893 8435 20927
rect 8435 20893 8444 20927
rect 8392 20884 8444 20893
rect 10140 20884 10192 20936
rect 2780 20816 2832 20868
rect 4160 20816 4212 20868
rect 5724 20816 5776 20868
rect 6828 20816 6880 20868
rect 7012 20816 7064 20868
rect 4620 20748 4672 20800
rect 10048 20748 10100 20800
rect 12532 20791 12584 20800
rect 12532 20757 12541 20791
rect 12541 20757 12575 20791
rect 12575 20757 12584 20791
rect 12532 20748 12584 20757
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 5908 20544 5960 20596
rect 6736 20544 6788 20596
rect 8300 20544 8352 20596
rect 9496 20544 9548 20596
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 10140 20544 10192 20596
rect 10968 20544 11020 20596
rect 11152 20544 11204 20596
rect 12532 20408 12584 20460
rect 10048 20383 10100 20392
rect 10048 20349 10082 20383
rect 10082 20349 10100 20383
rect 10048 20340 10100 20349
rect 11152 20340 11204 20392
rect 12348 20340 12400 20392
rect 5816 20272 5868 20324
rect 6460 20315 6512 20324
rect 6460 20281 6469 20315
rect 6469 20281 6503 20315
rect 6503 20281 6512 20315
rect 6460 20272 6512 20281
rect 6920 20272 6972 20324
rect 12072 20272 12124 20324
rect 5908 20204 5960 20256
rect 6092 20247 6144 20256
rect 6092 20213 6101 20247
rect 6101 20213 6135 20247
rect 6135 20213 6144 20247
rect 6092 20204 6144 20213
rect 10968 20204 11020 20256
rect 12348 20204 12400 20256
rect 12440 20247 12492 20256
rect 12440 20213 12449 20247
rect 12449 20213 12483 20247
rect 12483 20213 12492 20247
rect 12440 20204 12492 20213
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 6828 20000 6880 20052
rect 8392 20000 8444 20052
rect 10508 20000 10560 20052
rect 12348 20000 12400 20052
rect 9956 19907 10008 19916
rect 9956 19873 9965 19907
rect 9965 19873 9999 19907
rect 9999 19873 10008 19907
rect 9956 19864 10008 19873
rect 11244 19864 11296 19916
rect 11152 19839 11204 19848
rect 11152 19805 11161 19839
rect 11161 19805 11195 19839
rect 11195 19805 11204 19839
rect 11152 19796 11204 19805
rect 2780 19703 2832 19712
rect 2780 19669 2789 19703
rect 2789 19669 2823 19703
rect 2823 19669 2832 19703
rect 2780 19660 2832 19669
rect 5264 19660 5316 19712
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 8208 19660 8260 19712
rect 10508 19660 10560 19712
rect 12992 19660 13044 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 10048 19456 10100 19508
rect 12532 19456 12584 19508
rect 4252 19388 4304 19440
rect 4804 19388 4856 19440
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 10508 19363 10560 19372
rect 10508 19329 10517 19363
rect 10517 19329 10551 19363
rect 10551 19329 10560 19363
rect 10508 19320 10560 19329
rect 11244 19320 11296 19372
rect 12532 19320 12584 19372
rect 12992 19363 13044 19372
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 9956 19252 10008 19304
rect 11060 19252 11112 19304
rect 5172 19184 5224 19236
rect 7564 19227 7616 19236
rect 7564 19193 7573 19227
rect 7573 19193 7607 19227
rect 7607 19193 7616 19227
rect 7564 19184 7616 19193
rect 11796 19227 11848 19236
rect 11796 19193 11805 19227
rect 11805 19193 11839 19227
rect 11839 19193 11848 19227
rect 11796 19184 11848 19193
rect 12624 19184 12676 19236
rect 4068 19116 4120 19168
rect 4528 19159 4580 19168
rect 4528 19125 4537 19159
rect 4537 19125 4571 19159
rect 4571 19125 4580 19159
rect 4528 19116 4580 19125
rect 4988 19159 5040 19168
rect 4988 19125 4997 19159
rect 4997 19125 5031 19159
rect 5031 19125 5040 19159
rect 4988 19116 5040 19125
rect 5264 19116 5316 19168
rect 6828 19116 6880 19168
rect 8760 19116 8812 19168
rect 10048 19159 10100 19168
rect 10048 19125 10057 19159
rect 10057 19125 10091 19159
rect 10091 19125 10100 19159
rect 10048 19116 10100 19125
rect 11244 19159 11296 19168
rect 11244 19125 11253 19159
rect 11253 19125 11287 19159
rect 11287 19125 11296 19159
rect 11244 19116 11296 19125
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 4988 18912 5040 18964
rect 5448 18912 5500 18964
rect 6736 18955 6788 18964
rect 6736 18921 6745 18955
rect 6745 18921 6779 18955
rect 6779 18921 6788 18955
rect 6736 18912 6788 18921
rect 10324 18912 10376 18964
rect 10600 18912 10652 18964
rect 11152 18912 11204 18964
rect 12072 18912 12124 18964
rect 1676 18887 1728 18896
rect 1676 18853 1685 18887
rect 1685 18853 1719 18887
rect 1719 18853 1728 18887
rect 1676 18844 1728 18853
rect 4252 18844 4304 18896
rect 4804 18844 4856 18896
rect 10140 18887 10192 18896
rect 10140 18853 10149 18887
rect 10149 18853 10183 18887
rect 10183 18853 10192 18887
rect 10140 18844 10192 18853
rect 11336 18844 11388 18896
rect 11888 18844 11940 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 7104 18819 7156 18828
rect 7104 18785 7113 18819
rect 7113 18785 7147 18819
rect 7147 18785 7156 18819
rect 7104 18776 7156 18785
rect 10600 18776 10652 18828
rect 11520 18776 11572 18828
rect 12348 18819 12400 18828
rect 12348 18785 12357 18819
rect 12357 18785 12391 18819
rect 12391 18785 12400 18819
rect 12348 18776 12400 18785
rect 3976 18708 4028 18760
rect 7196 18751 7248 18760
rect 7196 18717 7205 18751
rect 7205 18717 7239 18751
rect 7239 18717 7248 18751
rect 7196 18708 7248 18717
rect 6644 18640 6696 18692
rect 6920 18640 6972 18692
rect 8208 18708 8260 18760
rect 9680 18708 9732 18760
rect 9864 18708 9916 18760
rect 9588 18640 9640 18692
rect 9956 18640 10008 18692
rect 10968 18708 11020 18760
rect 12532 18751 12584 18760
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 5540 18572 5592 18624
rect 9680 18615 9732 18624
rect 9680 18581 9689 18615
rect 9689 18581 9723 18615
rect 9723 18581 9732 18615
rect 9680 18572 9732 18581
rect 11060 18615 11112 18624
rect 11060 18581 11069 18615
rect 11069 18581 11103 18615
rect 11103 18581 11112 18615
rect 11060 18572 11112 18581
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 6644 18411 6696 18420
rect 6644 18377 6653 18411
rect 6653 18377 6687 18411
rect 6687 18377 6696 18411
rect 6644 18368 6696 18377
rect 7196 18368 7248 18420
rect 7840 18368 7892 18420
rect 10140 18411 10192 18420
rect 10140 18377 10149 18411
rect 10149 18377 10183 18411
rect 10183 18377 10192 18411
rect 10140 18368 10192 18377
rect 10508 18368 10560 18420
rect 4160 18300 4212 18352
rect 8208 18343 8260 18352
rect 8208 18309 8217 18343
rect 8217 18309 8251 18343
rect 8251 18309 8260 18343
rect 8208 18300 8260 18309
rect 10692 18300 10744 18352
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 2964 18164 3016 18216
rect 3976 18164 4028 18216
rect 2228 18139 2280 18148
rect 2228 18105 2237 18139
rect 2237 18105 2271 18139
rect 2271 18105 2280 18139
rect 2228 18096 2280 18105
rect 3056 18096 3108 18148
rect 4068 18096 4120 18148
rect 9588 18275 9640 18284
rect 9588 18241 9597 18275
rect 9597 18241 9631 18275
rect 9631 18241 9640 18275
rect 9588 18232 9640 18241
rect 10324 18232 10376 18284
rect 12348 18232 12400 18284
rect 5448 18207 5500 18216
rect 5448 18173 5457 18207
rect 5457 18173 5491 18207
rect 5491 18173 5500 18207
rect 5448 18164 5500 18173
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 8300 18164 8352 18216
rect 8576 18164 8628 18216
rect 12256 18164 12308 18216
rect 13912 18164 13964 18216
rect 8116 18096 8168 18148
rect 10232 18096 10284 18148
rect 11060 18139 11112 18148
rect 11060 18105 11069 18139
rect 11069 18105 11103 18139
rect 11103 18105 11112 18139
rect 11060 18096 11112 18105
rect 11888 18096 11940 18148
rect 4252 18071 4304 18080
rect 4252 18037 4261 18071
rect 4261 18037 4295 18071
rect 4295 18037 4304 18071
rect 4252 18028 4304 18037
rect 5448 18028 5500 18080
rect 8944 18028 8996 18080
rect 9312 18028 9364 18080
rect 9864 18028 9916 18080
rect 10048 18028 10100 18080
rect 10508 18071 10560 18080
rect 10508 18037 10517 18071
rect 10517 18037 10551 18071
rect 10551 18037 10560 18071
rect 10508 18028 10560 18037
rect 10968 18071 11020 18080
rect 10968 18037 10977 18071
rect 10977 18037 11011 18071
rect 11011 18037 11020 18071
rect 10968 18028 11020 18037
rect 11428 18028 11480 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 1400 17824 1452 17876
rect 1768 17824 1820 17876
rect 4068 17824 4120 17876
rect 5264 17824 5316 17876
rect 7104 17824 7156 17876
rect 11060 17867 11112 17876
rect 11060 17833 11069 17867
rect 11069 17833 11103 17867
rect 11103 17833 11112 17867
rect 11060 17824 11112 17833
rect 5540 17756 5592 17808
rect 9956 17799 10008 17808
rect 9956 17765 9990 17799
rect 9990 17765 10008 17799
rect 9956 17756 10008 17765
rect 2780 17688 2832 17740
rect 4620 17688 4672 17740
rect 5448 17688 5500 17740
rect 7932 17731 7984 17740
rect 7932 17697 7941 17731
rect 7941 17697 7975 17731
rect 7975 17697 7984 17731
rect 7932 17688 7984 17697
rect 8944 17688 8996 17740
rect 9772 17688 9824 17740
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 4252 17620 4304 17672
rect 4896 17620 4948 17672
rect 5172 17620 5224 17672
rect 8116 17663 8168 17672
rect 8116 17629 8125 17663
rect 8125 17629 8159 17663
rect 8159 17629 8168 17663
rect 8116 17620 8168 17629
rect 8852 17620 8904 17672
rect 7104 17552 7156 17604
rect 2412 17527 2464 17536
rect 2412 17493 2421 17527
rect 2421 17493 2455 17527
rect 2455 17493 2464 17527
rect 2412 17484 2464 17493
rect 4068 17484 4120 17536
rect 4528 17484 4580 17536
rect 4988 17484 5040 17536
rect 6736 17527 6788 17536
rect 6736 17493 6745 17527
rect 6745 17493 6779 17527
rect 6779 17493 6788 17527
rect 6736 17484 6788 17493
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 8576 17484 8628 17536
rect 11336 17527 11388 17536
rect 11336 17493 11345 17527
rect 11345 17493 11379 17527
rect 11379 17493 11388 17527
rect 11336 17484 11388 17493
rect 11888 17484 11940 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 1768 17323 1820 17332
rect 1768 17289 1777 17323
rect 1777 17289 1811 17323
rect 1811 17289 1820 17323
rect 1768 17280 1820 17289
rect 2872 17323 2924 17332
rect 2872 17289 2881 17323
rect 2881 17289 2915 17323
rect 2915 17289 2924 17323
rect 2872 17280 2924 17289
rect 5448 17280 5500 17332
rect 8116 17280 8168 17332
rect 8852 17323 8904 17332
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 9956 17280 10008 17332
rect 10600 17323 10652 17332
rect 10600 17289 10609 17323
rect 10609 17289 10643 17323
rect 10643 17289 10652 17323
rect 10600 17280 10652 17289
rect 10968 17280 11020 17332
rect 11336 17280 11388 17332
rect 2964 17212 3016 17264
rect 9772 17212 9824 17264
rect 11520 17212 11572 17264
rect 3056 17144 3108 17196
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 10324 17144 10376 17196
rect 11244 17144 11296 17196
rect 11888 17144 11940 17196
rect 12072 17144 12124 17196
rect 2964 17076 3016 17128
rect 4344 17119 4396 17128
rect 2504 17008 2556 17060
rect 4344 17085 4353 17119
rect 4353 17085 4387 17119
rect 4387 17085 4396 17119
rect 4344 17076 4396 17085
rect 4712 17076 4764 17128
rect 5172 17076 5224 17128
rect 7012 17076 7064 17128
rect 8300 17076 8352 17128
rect 9772 17076 9824 17128
rect 10416 17076 10468 17128
rect 10600 17076 10652 17128
rect 12164 17076 12216 17128
rect 3608 16940 3660 16992
rect 4068 16940 4120 16992
rect 6828 17008 6880 17060
rect 7196 17008 7248 17060
rect 7748 17008 7800 17060
rect 7932 17008 7984 17060
rect 10784 17008 10836 17060
rect 12624 17008 12676 17060
rect 5540 16983 5592 16992
rect 5540 16949 5549 16983
rect 5549 16949 5583 16983
rect 5583 16949 5592 16983
rect 5540 16940 5592 16949
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 11244 16983 11296 16992
rect 11244 16949 11253 16983
rect 11253 16949 11287 16983
rect 11287 16949 11296 16983
rect 11244 16940 11296 16949
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 2872 16736 2924 16788
rect 3056 16736 3108 16788
rect 3608 16736 3660 16788
rect 4160 16736 4212 16788
rect 4620 16736 4672 16788
rect 5724 16736 5776 16788
rect 6736 16736 6788 16788
rect 7840 16779 7892 16788
rect 7840 16745 7849 16779
rect 7849 16745 7883 16779
rect 7883 16745 7892 16779
rect 7840 16736 7892 16745
rect 8668 16736 8720 16788
rect 8852 16736 8904 16788
rect 9588 16736 9640 16788
rect 10232 16779 10284 16788
rect 10232 16745 10241 16779
rect 10241 16745 10275 16779
rect 10275 16745 10284 16779
rect 10232 16736 10284 16745
rect 11244 16779 11296 16788
rect 11244 16745 11253 16779
rect 11253 16745 11287 16779
rect 11287 16745 11296 16779
rect 11244 16736 11296 16745
rect 12072 16736 12124 16788
rect 3976 16668 4028 16720
rect 6184 16668 6236 16720
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 4160 16532 4212 16584
rect 4988 16532 5040 16584
rect 5908 16532 5960 16584
rect 6644 16532 6696 16584
rect 8116 16668 8168 16720
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 8668 16600 8720 16652
rect 10600 16643 10652 16652
rect 10600 16609 10609 16643
rect 10609 16609 10643 16643
rect 10643 16609 10652 16643
rect 10600 16600 10652 16609
rect 10692 16643 10744 16652
rect 10692 16609 10701 16643
rect 10701 16609 10735 16643
rect 10735 16609 10744 16643
rect 10692 16600 10744 16609
rect 11520 16600 11572 16652
rect 11888 16600 11940 16652
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 8392 16532 8444 16541
rect 10324 16532 10376 16584
rect 4528 16464 4580 16516
rect 7472 16464 7524 16516
rect 8484 16464 8536 16516
rect 5632 16439 5684 16448
rect 5632 16405 5641 16439
rect 5641 16405 5675 16439
rect 5675 16405 5684 16439
rect 5632 16396 5684 16405
rect 5908 16439 5960 16448
rect 5908 16405 5917 16439
rect 5917 16405 5951 16439
rect 5951 16405 5960 16439
rect 5908 16396 5960 16405
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 3976 16192 4028 16244
rect 4620 16192 4672 16244
rect 6184 16235 6236 16244
rect 6184 16201 6193 16235
rect 6193 16201 6227 16235
rect 6227 16201 6236 16235
rect 6184 16192 6236 16201
rect 6736 16192 6788 16244
rect 11244 16192 11296 16244
rect 11520 16192 11572 16244
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 7748 16056 7800 16108
rect 8484 16056 8536 16108
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 11152 16056 11204 16108
rect 11888 16056 11940 16108
rect 5172 15988 5224 16040
rect 5908 15988 5960 16040
rect 7472 16031 7524 16040
rect 7472 15997 7481 16031
rect 7481 15997 7515 16031
rect 7515 15997 7524 16031
rect 7472 15988 7524 15997
rect 7564 16031 7616 16040
rect 7564 15997 7573 16031
rect 7573 15997 7607 16031
rect 7607 15997 7616 16031
rect 7564 15988 7616 15997
rect 8024 15988 8076 16040
rect 9588 15988 9640 16040
rect 5356 15920 5408 15972
rect 6276 15920 6328 15972
rect 7196 15920 7248 15972
rect 8852 15920 8904 15972
rect 11336 15920 11388 15972
rect 4160 15852 4212 15904
rect 5448 15852 5500 15904
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 6000 15852 6052 15904
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 8024 15852 8076 15904
rect 8208 15852 8260 15904
rect 10416 15852 10468 15904
rect 12256 15852 12308 15904
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 3976 15648 4028 15700
rect 5172 15691 5224 15700
rect 5172 15657 5181 15691
rect 5181 15657 5215 15691
rect 5215 15657 5224 15691
rect 5172 15648 5224 15657
rect 5816 15648 5868 15700
rect 6184 15648 6236 15700
rect 6828 15691 6880 15700
rect 6828 15657 6837 15691
rect 6837 15657 6871 15691
rect 6871 15657 6880 15691
rect 6828 15648 6880 15657
rect 7656 15648 7708 15700
rect 7932 15648 7984 15700
rect 8208 15691 8260 15700
rect 8208 15657 8217 15691
rect 8217 15657 8251 15691
rect 8251 15657 8260 15691
rect 8208 15648 8260 15657
rect 8392 15648 8444 15700
rect 10600 15648 10652 15700
rect 4436 15623 4488 15632
rect 4436 15589 4445 15623
rect 4445 15589 4479 15623
rect 4479 15589 4488 15623
rect 4436 15580 4488 15589
rect 4712 15580 4764 15632
rect 5908 15580 5960 15632
rect 7104 15580 7156 15632
rect 8852 15580 8904 15632
rect 10324 15623 10376 15632
rect 10324 15589 10333 15623
rect 10333 15589 10367 15623
rect 10367 15589 10376 15623
rect 10324 15580 10376 15589
rect 10968 15580 11020 15632
rect 4252 15512 4304 15564
rect 7564 15512 7616 15564
rect 8208 15512 8260 15564
rect 8392 15512 8444 15564
rect 8576 15512 8628 15564
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 5356 15376 5408 15428
rect 6644 15444 6696 15496
rect 6828 15444 6880 15496
rect 7288 15444 7340 15496
rect 7932 15444 7984 15496
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 10048 15444 10100 15496
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 3516 15308 3568 15360
rect 5632 15351 5684 15360
rect 5632 15317 5641 15351
rect 5641 15317 5675 15351
rect 5675 15317 5684 15351
rect 5632 15308 5684 15317
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 2504 15104 2556 15156
rect 6000 15104 6052 15156
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 8668 15147 8720 15156
rect 8668 15113 8677 15147
rect 8677 15113 8711 15147
rect 8711 15113 8720 15147
rect 8668 15104 8720 15113
rect 9680 15104 9732 15156
rect 10048 15147 10100 15156
rect 10048 15113 10057 15147
rect 10057 15113 10091 15147
rect 10091 15113 10100 15147
rect 10048 15104 10100 15113
rect 10692 15104 10744 15156
rect 11152 15104 11204 15156
rect 5908 15036 5960 15088
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 4068 14968 4120 15020
rect 4804 14968 4856 15020
rect 5724 15011 5776 15020
rect 5724 14977 5733 15011
rect 5733 14977 5767 15011
rect 5767 14977 5776 15011
rect 5724 14968 5776 14977
rect 8208 15036 8260 15088
rect 6828 14968 6880 15020
rect 6920 14968 6972 15020
rect 7288 14968 7340 15020
rect 8852 14968 8904 15020
rect 9312 15011 9364 15020
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 9312 14968 9364 14977
rect 10968 14968 11020 15020
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 7472 14900 7524 14952
rect 8668 14900 8720 14952
rect 9404 14900 9456 14952
rect 10324 14900 10376 14952
rect 2228 14875 2280 14884
rect 2228 14841 2237 14875
rect 2237 14841 2271 14875
rect 2271 14841 2280 14875
rect 2228 14832 2280 14841
rect 5908 14832 5960 14884
rect 7564 14832 7616 14884
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 4252 14807 4304 14816
rect 3608 14764 3660 14773
rect 4252 14773 4261 14807
rect 4261 14773 4295 14807
rect 4295 14773 4304 14807
rect 4252 14764 4304 14773
rect 4712 14764 4764 14816
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 5632 14807 5684 14816
rect 5632 14773 5641 14807
rect 5641 14773 5675 14807
rect 5675 14773 5684 14807
rect 5632 14764 5684 14773
rect 6000 14764 6052 14816
rect 8852 14764 8904 14816
rect 10232 14764 10284 14816
rect 11244 14832 11296 14884
rect 10784 14764 10836 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 3608 14560 3660 14612
rect 5172 14560 5224 14612
rect 7012 14560 7064 14612
rect 7288 14603 7340 14612
rect 7288 14569 7297 14603
rect 7297 14569 7331 14603
rect 7331 14569 7340 14603
rect 7288 14560 7340 14569
rect 7472 14560 7524 14612
rect 8760 14560 8812 14612
rect 8852 14560 8904 14612
rect 9864 14560 9916 14612
rect 10968 14560 11020 14612
rect 11152 14603 11204 14612
rect 11152 14569 11161 14603
rect 11161 14569 11195 14603
rect 11195 14569 11204 14603
rect 11152 14560 11204 14569
rect 5540 14492 5592 14544
rect 6368 14492 6420 14544
rect 9588 14492 9640 14544
rect 9956 14492 10008 14544
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 4528 14467 4580 14476
rect 4528 14433 4537 14467
rect 4537 14433 4571 14467
rect 4571 14433 4580 14467
rect 5172 14467 5224 14476
rect 4528 14424 4580 14433
rect 5172 14433 5181 14467
rect 5181 14433 5215 14467
rect 5215 14433 5224 14467
rect 5172 14424 5224 14433
rect 5724 14424 5776 14476
rect 8484 14424 8536 14476
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 5816 14356 5868 14408
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 6736 14356 6788 14408
rect 9680 14356 9732 14408
rect 11520 14467 11572 14476
rect 11520 14433 11529 14467
rect 11529 14433 11563 14467
rect 11563 14433 11572 14467
rect 11520 14424 11572 14433
rect 11796 14467 11848 14476
rect 11796 14433 11830 14467
rect 11830 14433 11848 14467
rect 11796 14424 11848 14433
rect 4160 14288 4212 14340
rect 5632 14263 5684 14272
rect 5632 14229 5641 14263
rect 5641 14229 5675 14263
rect 5675 14229 5684 14263
rect 5632 14220 5684 14229
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 10140 14220 10192 14272
rect 10784 14220 10836 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 3516 14016 3568 14068
rect 4068 14016 4120 14068
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 7564 14016 7616 14068
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 9864 14016 9916 14068
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 10968 14016 11020 14068
rect 11520 14016 11572 14068
rect 8944 13948 8996 14000
rect 2780 13812 2832 13864
rect 3884 13855 3936 13864
rect 3884 13821 3893 13855
rect 3893 13821 3927 13855
rect 3927 13821 3936 13855
rect 3884 13812 3936 13821
rect 4160 13855 4212 13864
rect 4160 13821 4194 13855
rect 4194 13821 4212 13855
rect 4160 13812 4212 13821
rect 8392 13812 8444 13864
rect 8760 13812 8812 13864
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 9496 13880 9548 13932
rect 10048 13880 10100 13932
rect 8944 13812 8996 13821
rect 9680 13812 9732 13864
rect 11796 13812 11848 13864
rect 12348 13812 12400 13864
rect 4528 13744 4580 13796
rect 7196 13744 7248 13796
rect 5816 13676 5868 13728
rect 6184 13676 6236 13728
rect 8484 13719 8536 13728
rect 8484 13685 8493 13719
rect 8493 13685 8527 13719
rect 8527 13685 8536 13719
rect 8484 13676 8536 13685
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 2780 13472 2832 13524
rect 4160 13472 4212 13524
rect 8852 13515 8904 13524
rect 8852 13481 8861 13515
rect 8861 13481 8895 13515
rect 8895 13481 8904 13515
rect 8852 13472 8904 13481
rect 9588 13472 9640 13524
rect 1676 13447 1728 13456
rect 1676 13413 1685 13447
rect 1685 13413 1719 13447
rect 1719 13413 1728 13447
rect 1676 13404 1728 13413
rect 4436 13404 4488 13456
rect 5172 13447 5224 13456
rect 5172 13413 5206 13447
rect 5206 13413 5224 13447
rect 5172 13404 5224 13413
rect 8300 13404 8352 13456
rect 8760 13404 8812 13456
rect 9680 13404 9732 13456
rect 6736 13336 6788 13388
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 8208 13336 8260 13388
rect 1676 13268 1728 13320
rect 4620 13268 4672 13320
rect 9588 13268 9640 13320
rect 3884 13200 3936 13252
rect 6736 13200 6788 13252
rect 2504 13132 2556 13184
rect 5816 13132 5868 13184
rect 6092 13132 6144 13184
rect 6828 13132 6880 13184
rect 8852 13132 8904 13184
rect 9404 13132 9456 13184
rect 9956 13132 10008 13184
rect 10784 13132 10836 13184
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 4160 12928 4212 12980
rect 5172 12928 5224 12980
rect 4620 12860 4672 12912
rect 2504 12767 2556 12776
rect 2504 12733 2513 12767
rect 2513 12733 2547 12767
rect 2547 12733 2556 12767
rect 2504 12724 2556 12733
rect 3148 12724 3200 12776
rect 3976 12724 4028 12776
rect 7104 12928 7156 12980
rect 7564 12928 7616 12980
rect 8208 12971 8260 12980
rect 8208 12937 8217 12971
rect 8217 12937 8251 12971
rect 8251 12937 8260 12971
rect 8208 12928 8260 12937
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 10048 12928 10100 12980
rect 10416 12928 10468 12980
rect 6736 12724 6788 12776
rect 10508 12860 10560 12912
rect 11520 12928 11572 12980
rect 9036 12767 9088 12776
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9036 12724 9088 12733
rect 9588 12724 9640 12776
rect 10048 12724 10100 12776
rect 2688 12656 2740 12708
rect 6644 12656 6696 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 7840 12656 7892 12708
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 9680 12588 9732 12640
rect 10140 12588 10192 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 4620 12384 4672 12436
rect 5080 12384 5132 12436
rect 5540 12384 5592 12436
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 4988 12316 5040 12368
rect 6552 12316 6604 12368
rect 6920 12316 6972 12368
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 6828 12291 6880 12300
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 8208 12248 8260 12300
rect 9864 12248 9916 12300
rect 10876 12291 10928 12300
rect 10876 12257 10885 12291
rect 10885 12257 10919 12291
rect 10919 12257 10928 12291
rect 10876 12248 10928 12257
rect 10968 12248 11020 12300
rect 6644 12180 6696 12232
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 6736 12112 6788 12164
rect 8852 12180 8904 12232
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 10508 12180 10560 12232
rect 9036 12112 9088 12164
rect 1768 12044 1820 12096
rect 2504 12087 2556 12096
rect 2504 12053 2513 12087
rect 2513 12053 2547 12087
rect 2547 12053 2556 12087
rect 2504 12044 2556 12053
rect 5172 12044 5224 12096
rect 5724 12044 5776 12096
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 7380 12044 7432 12096
rect 7564 12087 7616 12096
rect 7564 12053 7573 12087
rect 7573 12053 7607 12087
rect 7607 12053 7616 12087
rect 7564 12044 7616 12053
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 10508 12087 10560 12096
rect 10508 12053 10517 12087
rect 10517 12053 10551 12087
rect 10551 12053 10560 12087
rect 10508 12044 10560 12053
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 5080 11840 5132 11892
rect 6736 11840 6788 11892
rect 6828 11840 6880 11892
rect 8208 11840 8260 11892
rect 10048 11883 10100 11892
rect 10048 11849 10057 11883
rect 10057 11849 10091 11883
rect 10091 11849 10100 11883
rect 10048 11840 10100 11849
rect 10876 11840 10928 11892
rect 11520 11840 11572 11892
rect 5816 11772 5868 11824
rect 8300 11772 8352 11824
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 5724 11747 5776 11756
rect 5724 11713 5733 11747
rect 5733 11713 5767 11747
rect 5767 11713 5776 11747
rect 5724 11704 5776 11713
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 8668 11704 8720 11756
rect 8852 11704 8904 11756
rect 5816 11636 5868 11688
rect 6000 11636 6052 11688
rect 8024 11636 8076 11688
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 4988 11543 5040 11552
rect 4988 11509 4997 11543
rect 4997 11509 5031 11543
rect 5031 11509 5040 11543
rect 4988 11500 5040 11509
rect 6828 11568 6880 11620
rect 10508 11636 10560 11688
rect 10968 11704 11020 11756
rect 8760 11500 8812 11552
rect 9404 11500 9456 11552
rect 9588 11543 9640 11552
rect 9588 11509 9597 11543
rect 9597 11509 9631 11543
rect 9631 11509 9640 11543
rect 9588 11500 9640 11509
rect 10048 11500 10100 11552
rect 11428 11500 11480 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 4804 11339 4856 11348
rect 4804 11305 4813 11339
rect 4813 11305 4847 11339
rect 4847 11305 4856 11339
rect 4804 11296 4856 11305
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 7840 11296 7892 11305
rect 8024 11339 8076 11348
rect 8024 11305 8033 11339
rect 8033 11305 8067 11339
rect 8067 11305 8076 11339
rect 8024 11296 8076 11305
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 8852 11296 8904 11348
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 10416 11296 10468 11348
rect 11060 11296 11112 11348
rect 11520 11296 11572 11348
rect 1676 11160 1728 11212
rect 2412 11160 2464 11212
rect 4068 11160 4120 11212
rect 5448 11228 5500 11280
rect 7012 11228 7064 11280
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 4712 11092 4764 11144
rect 5540 11024 5592 11076
rect 9680 11228 9732 11280
rect 11428 11228 11480 11280
rect 6644 11092 6696 11144
rect 11060 11160 11112 11212
rect 11980 11160 12032 11212
rect 12256 11160 12308 11212
rect 2412 10956 2464 11008
rect 7564 10956 7616 11008
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 11152 11024 11204 11076
rect 8852 10956 8904 11008
rect 10784 10956 10836 11008
rect 11336 10956 11388 11008
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 4068 10752 4120 10804
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 5540 10752 5592 10804
rect 6920 10752 6972 10804
rect 8300 10752 8352 10804
rect 9680 10795 9732 10804
rect 9680 10761 9689 10795
rect 9689 10761 9723 10795
rect 9723 10761 9732 10795
rect 9680 10752 9732 10761
rect 10600 10795 10652 10804
rect 10600 10761 10609 10795
rect 10609 10761 10643 10795
rect 10643 10761 10652 10795
rect 10600 10752 10652 10761
rect 10968 10752 11020 10804
rect 11152 10752 11204 10804
rect 8484 10684 8536 10736
rect 2688 10659 2740 10668
rect 2688 10625 2697 10659
rect 2697 10625 2731 10659
rect 2731 10625 2740 10659
rect 2688 10616 2740 10625
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 7012 10616 7064 10668
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 8852 10616 8904 10668
rect 11520 10684 11572 10736
rect 12624 10684 12676 10736
rect 11336 10659 11388 10668
rect 11336 10625 11345 10659
rect 11345 10625 11379 10659
rect 11379 10625 11388 10659
rect 11336 10616 11388 10625
rect 6184 10548 6236 10600
rect 9036 10591 9088 10600
rect 9036 10557 9045 10591
rect 9045 10557 9079 10591
rect 9079 10557 9088 10591
rect 9036 10548 9088 10557
rect 9404 10548 9456 10600
rect 12348 10548 12400 10600
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 15752 10548 15804 10600
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 2136 10412 2188 10421
rect 2412 10480 2464 10532
rect 11336 10480 11388 10532
rect 11612 10480 11664 10532
rect 12440 10480 12492 10532
rect 12900 10523 12952 10532
rect 12900 10489 12909 10523
rect 12909 10489 12943 10523
rect 12943 10489 12952 10523
rect 12900 10480 12952 10489
rect 3424 10412 3476 10464
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 6092 10412 6144 10464
rect 6644 10412 6696 10464
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 8944 10455 8996 10464
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 2688 10208 2740 10260
rect 3424 10208 3476 10260
rect 5540 10208 5592 10260
rect 6828 10208 6880 10260
rect 7012 10208 7064 10260
rect 7196 10208 7248 10260
rect 8116 10251 8168 10260
rect 8116 10217 8125 10251
rect 8125 10217 8159 10251
rect 8159 10217 8168 10251
rect 8116 10208 8168 10217
rect 8852 10208 8904 10260
rect 10968 10208 11020 10260
rect 11428 10208 11480 10260
rect 7564 10140 7616 10192
rect 8300 10140 8352 10192
rect 9036 10140 9088 10192
rect 10784 10140 10836 10192
rect 12992 10140 13044 10192
rect 2044 10115 2096 10124
rect 2044 10081 2078 10115
rect 2078 10081 2096 10115
rect 2044 10072 2096 10081
rect 5448 10072 5500 10124
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 8484 10072 8536 10124
rect 9312 10072 9364 10124
rect 10416 10072 10468 10124
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 7564 10047 7616 10056
rect 4620 10004 4672 10013
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 8852 10004 8904 10056
rect 5080 9936 5132 9988
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 3056 9664 3108 9716
rect 3148 9664 3200 9716
rect 4528 9664 4580 9716
rect 7196 9707 7248 9716
rect 7196 9673 7205 9707
rect 7205 9673 7239 9707
rect 7239 9673 7248 9707
rect 7196 9664 7248 9673
rect 7380 9664 7432 9716
rect 9312 9664 9364 9716
rect 10416 9664 10468 9716
rect 10692 9664 10744 9716
rect 2044 9596 2096 9648
rect 3884 9596 3936 9648
rect 4620 9596 4672 9648
rect 8852 9639 8904 9648
rect 5448 9528 5500 9580
rect 7288 9528 7340 9580
rect 8116 9528 8168 9580
rect 8852 9605 8861 9639
rect 8861 9605 8895 9639
rect 8895 9605 8904 9639
rect 8852 9596 8904 9605
rect 10968 9596 11020 9648
rect 10784 9528 10836 9580
rect 2688 9460 2740 9512
rect 5264 9392 5316 9444
rect 9128 9435 9180 9444
rect 9128 9401 9137 9435
rect 9137 9401 9171 9435
rect 9171 9401 9180 9435
rect 9128 9392 9180 9401
rect 3240 9324 3292 9376
rect 4620 9324 4672 9376
rect 4988 9324 5040 9376
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 9312 9367 9364 9376
rect 9312 9333 9321 9367
rect 9321 9333 9355 9367
rect 9355 9333 9364 9367
rect 9312 9324 9364 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 1768 9163 1820 9172
rect 1768 9129 1777 9163
rect 1777 9129 1811 9163
rect 1811 9129 1820 9163
rect 1768 9120 1820 9129
rect 5540 9120 5592 9172
rect 6000 9120 6052 9172
rect 6184 9120 6236 9172
rect 6920 9163 6972 9172
rect 6920 9129 6929 9163
rect 6929 9129 6963 9163
rect 6963 9129 6972 9163
rect 6920 9120 6972 9129
rect 7564 9120 7616 9172
rect 9956 9120 10008 9172
rect 10232 9120 10284 9172
rect 2504 9052 2556 9104
rect 3332 8984 3384 9036
rect 3884 9027 3936 9036
rect 3884 8993 3893 9027
rect 3893 8993 3927 9027
rect 3927 8993 3936 9027
rect 3884 8984 3936 8993
rect 4988 8984 5040 9036
rect 6000 9027 6052 9036
rect 6000 8993 6009 9027
rect 6009 8993 6043 9027
rect 6043 8993 6052 9027
rect 6000 8984 6052 8993
rect 8208 8984 8260 9036
rect 3240 8916 3292 8968
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 4804 8916 4856 8968
rect 7380 8959 7432 8968
rect 5448 8891 5500 8900
rect 5448 8857 5457 8891
rect 5457 8857 5491 8891
rect 5491 8857 5500 8891
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 9312 8916 9364 8968
rect 9496 8916 9548 8968
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 5448 8848 5500 8857
rect 8852 8848 8904 8900
rect 2780 8780 2832 8832
rect 4528 8780 4580 8832
rect 5908 8780 5960 8832
rect 9496 8780 9548 8832
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 2504 8576 2556 8585
rect 4528 8576 4580 8628
rect 5448 8576 5500 8628
rect 5816 8576 5868 8628
rect 6184 8508 6236 8560
rect 6644 8508 6696 8560
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 1676 8372 1728 8424
rect 2136 8372 2188 8424
rect 2688 8372 2740 8424
rect 5356 8372 5408 8424
rect 7104 8415 7156 8424
rect 3792 8347 3844 8356
rect 3792 8313 3801 8347
rect 3801 8313 3835 8347
rect 3835 8313 3844 8347
rect 3792 8304 3844 8313
rect 4160 8304 4212 8356
rect 4804 8304 4856 8356
rect 5540 8304 5592 8356
rect 6000 8304 6052 8356
rect 7104 8381 7138 8415
rect 7138 8381 7156 8415
rect 7104 8372 7156 8381
rect 7380 8372 7432 8424
rect 2872 8236 2924 8288
rect 3424 8236 3476 8288
rect 9220 8372 9272 8424
rect 9956 8372 10008 8424
rect 7564 8236 7616 8288
rect 8208 8279 8260 8288
rect 8208 8245 8217 8279
rect 8217 8245 8251 8279
rect 8251 8245 8260 8279
rect 8208 8236 8260 8245
rect 8760 8236 8812 8288
rect 8944 8236 8996 8288
rect 11428 8236 11480 8288
rect 11980 8236 12032 8288
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 2412 8075 2464 8084
rect 2412 8041 2421 8075
rect 2421 8041 2455 8075
rect 2455 8041 2464 8075
rect 2412 8032 2464 8041
rect 2780 8032 2832 8084
rect 4068 8032 4120 8084
rect 5540 8032 5592 8084
rect 6828 8032 6880 8084
rect 8208 8032 8260 8084
rect 10232 8075 10284 8084
rect 10232 8041 10241 8075
rect 10241 8041 10275 8075
rect 10275 8041 10284 8075
rect 10232 8032 10284 8041
rect 12072 8032 12124 8084
rect 13268 8032 13320 8084
rect 3240 7964 3292 8016
rect 4988 7964 5040 8016
rect 7564 7964 7616 8016
rect 9220 7964 9272 8016
rect 2872 7896 2924 7948
rect 3148 7896 3200 7948
rect 5448 7896 5500 7948
rect 6092 7896 6144 7948
rect 8852 7896 8904 7948
rect 3332 7828 3384 7880
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 7840 7828 7892 7880
rect 3424 7692 3476 7744
rect 4068 7692 4120 7744
rect 8208 7692 8260 7744
rect 8944 7828 8996 7880
rect 9496 7964 9548 8016
rect 9956 8007 10008 8016
rect 9956 7973 9965 8007
rect 9965 7973 9999 8007
rect 9999 7973 10008 8007
rect 9956 7964 10008 7973
rect 10140 7964 10192 8016
rect 10876 7896 10928 7948
rect 11060 7896 11112 7948
rect 10232 7760 10284 7812
rect 8668 7692 8720 7744
rect 8760 7692 8812 7744
rect 9588 7692 9640 7744
rect 12348 7735 12400 7744
rect 12348 7701 12357 7735
rect 12357 7701 12391 7735
rect 12391 7701 12400 7735
rect 12348 7692 12400 7701
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 3148 7531 3200 7540
rect 2780 7488 2832 7497
rect 3148 7497 3157 7531
rect 3157 7497 3191 7531
rect 3191 7497 3200 7531
rect 3148 7488 3200 7497
rect 3332 7420 3384 7472
rect 5080 7488 5132 7540
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 7840 7531 7892 7540
rect 7840 7497 7849 7531
rect 7849 7497 7883 7531
rect 7883 7497 7892 7531
rect 7840 7488 7892 7497
rect 10876 7488 10928 7540
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 5908 7420 5960 7472
rect 8944 7463 8996 7472
rect 8944 7429 8953 7463
rect 8953 7429 8987 7463
rect 8987 7429 8996 7463
rect 8944 7420 8996 7429
rect 10232 7352 10284 7404
rect 12348 7352 12400 7404
rect 6184 7284 6236 7336
rect 8668 7284 8720 7336
rect 9772 7284 9824 7336
rect 10416 7284 10468 7336
rect 7472 7216 7524 7268
rect 5448 7148 5500 7200
rect 6092 7148 6144 7200
rect 6736 7148 6788 7200
rect 8116 7148 8168 7200
rect 9220 7191 9272 7200
rect 9220 7157 9229 7191
rect 9229 7157 9263 7191
rect 9263 7157 9272 7191
rect 9220 7148 9272 7157
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 10968 7148 11020 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 2044 6944 2096 6996
rect 3424 6944 3476 6996
rect 7840 6944 7892 6996
rect 8852 6944 8904 6996
rect 9404 6944 9456 6996
rect 10232 6987 10284 6996
rect 10232 6953 10241 6987
rect 10241 6953 10275 6987
rect 10275 6953 10284 6987
rect 10232 6944 10284 6953
rect 7472 6876 7524 6928
rect 1584 6808 1636 6860
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 5080 6851 5132 6860
rect 5080 6817 5089 6851
rect 5089 6817 5123 6851
rect 5123 6817 5132 6851
rect 5080 6808 5132 6817
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 8392 6851 8444 6860
rect 8392 6817 8401 6851
rect 8401 6817 8435 6851
rect 8435 6817 8444 6851
rect 8392 6808 8444 6817
rect 8484 6808 8536 6860
rect 8760 6808 8812 6860
rect 7932 6740 7984 6792
rect 8668 6783 8720 6792
rect 8668 6749 8677 6783
rect 8677 6749 8711 6783
rect 8711 6749 8720 6783
rect 8668 6740 8720 6749
rect 572 6672 624 6724
rect 4896 6672 4948 6724
rect 8300 6672 8352 6724
rect 9772 6876 9824 6928
rect 9496 6808 9548 6860
rect 10968 6808 11020 6860
rect 11152 6808 11204 6860
rect 1308 6604 1360 6656
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 5264 6604 5316 6613
rect 5448 6604 5500 6656
rect 5908 6604 5960 6656
rect 8484 6604 8536 6656
rect 9864 6647 9916 6656
rect 9864 6613 9873 6647
rect 9873 6613 9907 6647
rect 9907 6613 9916 6647
rect 9864 6604 9916 6613
rect 11060 6604 11112 6656
rect 11980 6604 12032 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 1400 6332 1452 6384
rect 2504 6400 2556 6452
rect 4988 6400 5040 6452
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 6184 6443 6236 6452
rect 6184 6409 6193 6443
rect 6193 6409 6227 6443
rect 6227 6409 6236 6443
rect 6184 6400 6236 6409
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 5724 6332 5776 6384
rect 6184 6264 6236 6316
rect 2044 6239 2096 6248
rect 2044 6205 2053 6239
rect 2053 6205 2087 6239
rect 2087 6205 2096 6239
rect 2044 6196 2096 6205
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 4712 6196 4764 6248
rect 4988 6196 5040 6248
rect 5540 6196 5592 6248
rect 8024 6400 8076 6452
rect 8392 6400 8444 6452
rect 11152 6400 11204 6452
rect 7932 6375 7984 6384
rect 7932 6341 7941 6375
rect 7941 6341 7975 6375
rect 7975 6341 7984 6375
rect 7932 6332 7984 6341
rect 9496 6332 9548 6384
rect 8668 6307 8720 6316
rect 8300 6196 8352 6248
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10232 6264 10284 6273
rect 8576 6196 8628 6248
rect 9680 6196 9732 6248
rect 11520 6196 11572 6248
rect 5540 6060 5592 6112
rect 7012 6060 7064 6112
rect 7932 6060 7984 6112
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 9496 6103 9548 6112
rect 8484 6060 8536 6069
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 9772 6060 9824 6112
rect 11060 6060 11112 6112
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 9772 5856 9824 5908
rect 10968 5856 11020 5908
rect 11244 5856 11296 5908
rect 8484 5788 8536 5840
rect 8852 5831 8904 5840
rect 8852 5797 8861 5831
rect 8861 5797 8895 5831
rect 8895 5797 8904 5831
rect 8852 5788 8904 5797
rect 3056 5720 3108 5772
rect 5080 5763 5132 5772
rect 5080 5729 5089 5763
rect 5089 5729 5123 5763
rect 5123 5729 5132 5763
rect 5080 5720 5132 5729
rect 6644 5720 6696 5772
rect 9680 5720 9732 5772
rect 5172 5695 5224 5704
rect 5172 5661 5181 5695
rect 5181 5661 5215 5695
rect 5215 5661 5224 5695
rect 5172 5652 5224 5661
rect 6920 5652 6972 5704
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 1768 5516 1820 5568
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 4068 5516 4120 5568
rect 5264 5516 5316 5568
rect 5448 5516 5500 5568
rect 7472 5627 7524 5636
rect 7472 5593 7481 5627
rect 7481 5593 7515 5627
rect 7515 5593 7524 5627
rect 7472 5584 7524 5593
rect 8392 5584 8444 5636
rect 11520 5720 11572 5772
rect 11152 5652 11204 5704
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 5908 5559 5960 5568
rect 5908 5525 5917 5559
rect 5917 5525 5951 5559
rect 5951 5525 5960 5559
rect 5908 5516 5960 5525
rect 7104 5516 7156 5568
rect 8116 5516 8168 5568
rect 8668 5516 8720 5568
rect 8852 5516 8904 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 4804 5355 4856 5364
rect 4804 5321 4813 5355
rect 4813 5321 4847 5355
rect 4847 5321 4856 5355
rect 4804 5312 4856 5321
rect 5264 5312 5316 5364
rect 5632 5312 5684 5364
rect 6644 5312 6696 5364
rect 8116 5312 8168 5364
rect 11980 5312 12032 5364
rect 3056 5244 3108 5296
rect 11060 5244 11112 5296
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 2412 5108 2464 5160
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 5632 5151 5684 5160
rect 5632 5117 5641 5151
rect 5641 5117 5675 5151
rect 5675 5117 5684 5151
rect 5632 5108 5684 5117
rect 5908 5108 5960 5160
rect 6920 5108 6972 5160
rect 7104 5151 7156 5160
rect 7104 5117 7138 5151
rect 7138 5117 7156 5151
rect 7104 5108 7156 5117
rect 11612 5108 11664 5160
rect 3976 5040 4028 5092
rect 9496 5040 9548 5092
rect 11520 5040 11572 5092
rect 5632 4972 5684 5024
rect 6644 4972 6696 5024
rect 7104 4972 7156 5024
rect 8208 5015 8260 5024
rect 8208 4981 8217 5015
rect 8217 4981 8251 5015
rect 8251 4981 8260 5015
rect 8208 4972 8260 4981
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 12716 4972 12768 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 2320 4700 2372 4752
rect 5264 4768 5316 4820
rect 6828 4768 6880 4820
rect 8576 4811 8628 4820
rect 8576 4777 8585 4811
rect 8585 4777 8619 4811
rect 8619 4777 8628 4811
rect 8576 4768 8628 4777
rect 9772 4768 9824 4820
rect 10232 4768 10284 4820
rect 11520 4768 11572 4820
rect 4068 4700 4120 4752
rect 6644 4700 6696 4752
rect 7380 4700 7432 4752
rect 8208 4700 8260 4752
rect 12440 4700 12492 4752
rect 4528 4675 4580 4684
rect 4528 4641 4537 4675
rect 4537 4641 4571 4675
rect 4571 4641 4580 4675
rect 4528 4632 4580 4641
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 12164 4675 12216 4684
rect 12164 4641 12173 4675
rect 12173 4641 12207 4675
rect 12207 4641 12216 4675
rect 12164 4632 12216 4641
rect 2872 4564 2924 4616
rect 3976 4564 4028 4616
rect 6828 4607 6880 4616
rect 3884 4539 3936 4548
rect 3884 4505 3893 4539
rect 3893 4505 3927 4539
rect 3927 4505 3936 4539
rect 3884 4496 3936 4505
rect 3424 4428 3476 4480
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 8300 4496 8352 4548
rect 9588 4496 9640 4548
rect 12900 4632 12952 4684
rect 12624 4564 12676 4616
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 5908 4428 5960 4480
rect 6828 4428 6880 4480
rect 8852 4428 8904 4480
rect 11336 4428 11388 4480
rect 12256 4428 12308 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 2872 4224 2924 4276
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 3332 4224 3384 4276
rect 3976 4224 4028 4276
rect 5172 4267 5224 4276
rect 5172 4233 5181 4267
rect 5181 4233 5215 4267
rect 5215 4233 5224 4267
rect 5172 4224 5224 4233
rect 6184 4267 6236 4276
rect 6184 4233 6193 4267
rect 6193 4233 6227 4267
rect 6227 4233 6236 4267
rect 6184 4224 6236 4233
rect 8392 4267 8444 4276
rect 8392 4233 8401 4267
rect 8401 4233 8435 4267
rect 8435 4233 8444 4267
rect 8392 4224 8444 4233
rect 10876 4224 10928 4276
rect 11152 4224 11204 4276
rect 1492 4020 1544 4072
rect 3056 3952 3108 4004
rect 5264 4156 5316 4208
rect 4528 4088 4580 4140
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 7196 4156 7248 4208
rect 7380 4156 7432 4208
rect 6920 4088 6972 4140
rect 7288 4088 7340 4140
rect 11244 4156 11296 4208
rect 12348 4156 12400 4208
rect 12624 4156 12676 4208
rect 7656 4088 7708 4140
rect 8576 4088 8628 4140
rect 9772 4088 9824 4140
rect 10324 4088 10376 4140
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 12900 4131 12952 4140
rect 10508 4088 10560 4097
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 4528 3952 4580 4004
rect 5448 3952 5500 4004
rect 4988 3884 5040 3936
rect 6184 3884 6236 3936
rect 7288 3927 7340 3936
rect 7288 3893 7297 3927
rect 7297 3893 7331 3927
rect 7331 3893 7340 3927
rect 9312 4020 9364 4072
rect 8760 3995 8812 4004
rect 8760 3961 8769 3995
rect 8769 3961 8803 3995
rect 8803 3961 8812 3995
rect 8760 3952 8812 3961
rect 10048 4020 10100 4072
rect 7288 3884 7340 3893
rect 8392 3884 8444 3936
rect 9312 3884 9364 3936
rect 11060 3952 11112 4004
rect 12624 3952 12676 4004
rect 10232 3884 10284 3936
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 12992 3884 13044 3936
rect 13360 3884 13412 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 1492 3680 1544 3732
rect 2320 3680 2372 3732
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 4988 3680 5040 3732
rect 5080 3680 5132 3732
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 7656 3680 7708 3732
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 8484 3680 8536 3732
rect 10600 3680 10652 3732
rect 10968 3680 11020 3732
rect 11152 3680 11204 3732
rect 2780 3655 2832 3664
rect 2780 3621 2789 3655
rect 2789 3621 2823 3655
rect 2823 3621 2832 3655
rect 2780 3612 2832 3621
rect 3148 3544 3200 3596
rect 4344 3544 4396 3596
rect 6000 3544 6052 3596
rect 6828 3612 6880 3664
rect 9680 3612 9732 3664
rect 12348 3680 12400 3732
rect 2688 3476 2740 3528
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 5816 3519 5868 3528
rect 1952 3408 2004 3460
rect 4436 3408 4488 3460
rect 5816 3485 5825 3519
rect 5825 3485 5859 3519
rect 5859 3485 5868 3519
rect 5816 3476 5868 3485
rect 6276 3476 6328 3528
rect 6920 3544 6972 3596
rect 8116 3476 8168 3528
rect 9956 3544 10008 3596
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 204 3340 256 3392
rect 1308 3340 1360 3392
rect 2412 3340 2464 3392
rect 3424 3340 3476 3392
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 4988 3383 5040 3392
rect 4988 3349 4997 3383
rect 4997 3349 5031 3383
rect 5031 3349 5040 3383
rect 4988 3340 5040 3349
rect 6920 3383 6972 3392
rect 6920 3349 6929 3383
rect 6929 3349 6963 3383
rect 6963 3349 6972 3383
rect 6920 3340 6972 3349
rect 7196 3340 7248 3392
rect 9312 3408 9364 3460
rect 10508 3476 10560 3528
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 2780 3136 2832 3188
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 6828 3136 6880 3188
rect 4436 3111 4488 3120
rect 4436 3077 4445 3111
rect 4445 3077 4479 3111
rect 4479 3077 4488 3111
rect 4436 3068 4488 3077
rect 4712 3111 4764 3120
rect 4712 3077 4721 3111
rect 4721 3077 4755 3111
rect 4755 3077 4764 3111
rect 6000 3111 6052 3120
rect 4712 3068 4764 3077
rect 6000 3077 6009 3111
rect 6009 3077 6043 3111
rect 6043 3077 6052 3111
rect 7840 3136 7892 3188
rect 8852 3136 8904 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 12440 3179 12492 3188
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 6000 3068 6052 3077
rect 8576 3068 8628 3120
rect 9404 3068 9456 3120
rect 1676 2932 1728 2984
rect 2412 2975 2464 2984
rect 2412 2941 2421 2975
rect 2421 2941 2455 2975
rect 2455 2941 2464 2975
rect 2412 2932 2464 2941
rect 5816 3000 5868 3052
rect 4988 2932 5040 2984
rect 7472 2932 7524 2984
rect 7656 2932 7708 2984
rect 8392 2932 8444 2984
rect 11152 3000 11204 3052
rect 13176 3000 13228 3052
rect 2228 2907 2280 2916
rect 2228 2873 2237 2907
rect 2237 2873 2271 2907
rect 2271 2873 2280 2907
rect 2228 2864 2280 2873
rect 7288 2864 7340 2916
rect 8116 2864 8168 2916
rect 7196 2796 7248 2848
rect 7472 2796 7524 2848
rect 9496 2932 9548 2984
rect 12532 2932 12584 2984
rect 9312 2864 9364 2916
rect 9588 2864 9640 2916
rect 13084 2864 13136 2916
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 1676 2635 1728 2644
rect 1676 2601 1685 2635
rect 1685 2601 1719 2635
rect 1719 2601 1728 2635
rect 1676 2592 1728 2601
rect 2412 2635 2464 2644
rect 2412 2601 2421 2635
rect 2421 2601 2455 2635
rect 2455 2601 2464 2635
rect 2412 2592 2464 2601
rect 2872 2592 2924 2644
rect 4344 2635 4396 2644
rect 4344 2601 4353 2635
rect 4353 2601 4387 2635
rect 4387 2601 4396 2635
rect 4344 2592 4396 2601
rect 4620 2635 4672 2644
rect 4620 2601 4629 2635
rect 4629 2601 4663 2635
rect 4663 2601 4672 2635
rect 4620 2592 4672 2601
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 7104 2592 7156 2644
rect 3884 2567 3936 2576
rect 3884 2533 3893 2567
rect 3893 2533 3927 2567
rect 3927 2533 3936 2567
rect 3884 2524 3936 2533
rect 2964 2456 3016 2508
rect 7564 2456 7616 2508
rect 8208 2592 8260 2644
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 10232 2592 10284 2644
rect 10692 2635 10744 2644
rect 10692 2601 10701 2635
rect 10701 2601 10735 2635
rect 10735 2601 10744 2635
rect 10692 2592 10744 2601
rect 11060 2592 11112 2644
rect 12716 2592 12768 2644
rect 13084 2635 13136 2644
rect 13084 2601 13093 2635
rect 13093 2601 13127 2635
rect 13127 2601 13136 2635
rect 13084 2592 13136 2601
rect 13452 2592 13504 2644
rect 10416 2456 10468 2508
rect 12072 2456 12124 2508
rect 13084 2456 13136 2508
rect 2964 2320 3016 2372
rect 5816 2388 5868 2440
rect 7656 2388 7708 2440
rect 11152 2388 11204 2440
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 12164 2320 12216 2372
rect 3332 2252 3384 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 3792 1980 3844 2032
rect 5632 1980 5684 2032
rect 11796 1368 11848 1420
rect 12256 1368 12308 1420
rect 9404 552 9456 604
rect 9496 552 9548 604
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1398 39520 1454 40000
rect 1766 39520 1822 40000
rect 2134 39520 2190 40000
rect 2594 39520 2650 40000
rect 2962 39520 3018 40000
rect 3330 39520 3386 40000
rect 3790 39520 3846 40000
rect 4158 39520 4214 40000
rect 4526 39520 4582 40000
rect 4986 39520 5042 40000
rect 5354 39520 5410 40000
rect 5722 39520 5778 40000
rect 6182 39520 6238 40000
rect 6550 39520 6606 40000
rect 6918 39520 6974 40000
rect 7378 39520 7434 40000
rect 7746 39520 7802 40000
rect 8206 39520 8262 40000
rect 8574 39520 8630 40000
rect 8942 39520 8998 40000
rect 9402 39520 9458 40000
rect 9770 39520 9826 40000
rect 10138 39522 10194 40000
rect 10138 39520 10272 39522
rect 10598 39520 10654 40000
rect 10966 39520 11022 40000
rect 11334 39520 11390 40000
rect 11794 39520 11850 40000
rect 12162 39520 12218 40000
rect 12530 39520 12586 40000
rect 12990 39520 13046 40000
rect 13358 39520 13414 40000
rect 13726 39520 13782 40000
rect 14186 39520 14242 40000
rect 14554 39520 14610 40000
rect 14922 39520 14978 40000
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 34678 244 39520
rect 584 34746 612 39520
rect 572 34740 624 34746
rect 572 34682 624 34688
rect 204 34672 256 34678
rect 204 34614 256 34620
rect 952 34202 980 39520
rect 1412 34678 1440 39520
rect 1490 34912 1546 34921
rect 1490 34847 1546 34856
rect 1308 34672 1360 34678
rect 1308 34614 1360 34620
rect 1400 34672 1452 34678
rect 1400 34614 1452 34620
rect 940 34196 992 34202
rect 940 34138 992 34144
rect 1320 33674 1348 34614
rect 1320 33658 1440 33674
rect 1320 33652 1452 33658
rect 1320 33646 1400 33652
rect 1400 33594 1452 33600
rect 1504 33046 1532 34847
rect 1780 34202 1808 39520
rect 2044 34536 2096 34542
rect 2044 34478 2096 34484
rect 1768 34196 1820 34202
rect 1768 34138 1820 34144
rect 2056 33969 2084 34478
rect 2042 33960 2098 33969
rect 2042 33895 2098 33904
rect 2148 33658 2176 39520
rect 2608 35329 2636 39520
rect 2778 38992 2834 39001
rect 2778 38927 2834 38936
rect 2594 35320 2650 35329
rect 2594 35255 2650 35264
rect 2412 34060 2464 34066
rect 2412 34002 2464 34008
rect 2136 33652 2188 33658
rect 2136 33594 2188 33600
rect 2424 33318 2452 34002
rect 2688 33448 2740 33454
rect 2688 33390 2740 33396
rect 2044 33312 2096 33318
rect 2044 33254 2096 33260
rect 2412 33312 2464 33318
rect 2412 33254 2464 33260
rect 1492 33040 1544 33046
rect 2056 33017 2084 33254
rect 2424 33153 2452 33254
rect 2410 33144 2466 33153
rect 2410 33079 2466 33088
rect 1492 32982 1544 32988
rect 1674 33008 1730 33017
rect 2042 33008 2098 33017
rect 1674 32943 1730 32952
rect 1768 32972 1820 32978
rect 1688 31958 1716 32943
rect 2042 32943 2098 32952
rect 1768 32914 1820 32920
rect 1780 32230 1808 32914
rect 2700 32774 2728 33390
rect 2688 32768 2740 32774
rect 2688 32710 2740 32716
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1676 31952 1728 31958
rect 1676 31894 1728 31900
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1688 31278 1716 31758
rect 1676 31272 1728 31278
rect 1674 31240 1676 31249
rect 1728 31240 1730 31249
rect 1674 31175 1730 31184
rect 1582 30968 1638 30977
rect 1582 30903 1638 30912
rect 1596 30258 1624 30903
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1582 30016 1638 30025
rect 1582 29951 1638 29960
rect 1400 29504 1452 29510
rect 1400 29446 1452 29452
rect 1412 25362 1440 29446
rect 1596 29306 1624 29951
rect 1584 29300 1636 29306
rect 1584 29242 1636 29248
rect 1582 28928 1638 28937
rect 1582 28863 1638 28872
rect 1492 26444 1544 26450
rect 1492 26386 1544 26392
rect 1504 25974 1532 26386
rect 1492 25968 1544 25974
rect 1492 25910 1544 25916
rect 1596 25906 1624 28863
rect 1674 27024 1730 27033
rect 1674 26959 1730 26968
rect 1688 26518 1716 26959
rect 1676 26512 1728 26518
rect 1676 26454 1728 26460
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1400 25356 1452 25362
rect 1400 25298 1452 25304
rect 1412 24954 1440 25298
rect 1584 25288 1636 25294
rect 1584 25230 1636 25236
rect 1596 24993 1624 25230
rect 1582 24984 1638 24993
rect 1400 24948 1452 24954
rect 1582 24919 1638 24928
rect 1400 24890 1452 24896
rect 1780 24177 1808 32166
rect 2226 30696 2282 30705
rect 2226 30631 2282 30640
rect 2240 30326 2268 30631
rect 2228 30320 2280 30326
rect 2228 30262 2280 30268
rect 2042 29200 2098 29209
rect 2042 29135 2044 29144
rect 2096 29135 2098 29144
rect 2044 29106 2096 29112
rect 2056 28218 2084 29106
rect 2044 28212 2096 28218
rect 2044 28154 2096 28160
rect 2056 28014 2084 28154
rect 2596 28144 2648 28150
rect 2596 28086 2648 28092
rect 2044 28008 2096 28014
rect 2044 27950 2096 27956
rect 2504 25696 2556 25702
rect 2504 25638 2556 25644
rect 2516 24857 2544 25638
rect 2502 24848 2558 24857
rect 2502 24783 2558 24792
rect 1766 24168 1822 24177
rect 1766 24103 1822 24112
rect 2412 22976 2464 22982
rect 1582 22944 1638 22953
rect 2412 22918 2464 22924
rect 1582 22879 1638 22888
rect 1596 22642 1624 22879
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 2424 22574 2452 22918
rect 1676 22568 1728 22574
rect 1676 22510 1728 22516
rect 2412 22568 2464 22574
rect 2412 22510 2464 22516
rect 1688 22234 1716 22510
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 1674 21040 1730 21049
rect 1674 20975 1730 20984
rect 1582 19000 1638 19009
rect 1582 18935 1638 18944
rect 1398 18864 1454 18873
rect 1398 18799 1400 18808
rect 1452 18799 1454 18808
rect 1400 18770 1452 18776
rect 1412 17882 1440 18770
rect 1596 18290 1624 18935
rect 1688 18902 1716 20975
rect 1676 18896 1728 18902
rect 1676 18838 1728 18844
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 2226 18184 2282 18193
rect 2226 18119 2228 18128
rect 2280 18119 2282 18128
rect 2228 18090 2280 18096
rect 1400 17876 1452 17882
rect 1400 17818 1452 17824
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1780 17338 1808 17818
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1582 16960 1638 16969
rect 1582 16895 1638 16904
rect 1596 15026 1624 16895
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1674 14920 1730 14929
rect 1674 14855 1730 14864
rect 2226 14920 2282 14929
rect 2226 14855 2228 14864
rect 1688 13462 1716 14855
rect 2280 14855 2282 14864
rect 2228 14826 2280 14832
rect 1676 13456 1728 13462
rect 1676 13398 1728 13404
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1582 13016 1638 13025
rect 1582 12951 1638 12960
rect 1596 11762 1624 12951
rect 1688 12646 1716 13262
rect 1676 12640 1728 12646
rect 1674 12608 1676 12617
rect 1728 12608 1730 12617
rect 1674 12543 1730 12552
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10985 1624 11086
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1688 10266 1716 11154
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1780 10062 1808 12038
rect 2228 11552 2280 11558
rect 2226 11520 2228 11529
rect 2280 11520 2282 11529
rect 2226 11455 2282 11464
rect 2424 11218 2452 17478
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2516 15162 2544 17002
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2516 12782 2544 13126
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2516 12102 2544 12718
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10538 2452 10950
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1780 9178 1808 9998
rect 2056 9654 2084 10066
rect 2044 9648 2096 9654
rect 2042 9616 2044 9625
rect 2096 9616 2098 9625
rect 2042 9551 2098 9560
rect 2056 9525 2084 9551
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8498 1624 8871
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 2148 8430 2176 10406
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 1688 8090 1716 8366
rect 2424 8090 2452 10474
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2516 8634 2544 9046
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2502 7440 2558 7449
rect 2502 7375 2558 7384
rect 2318 7032 2374 7041
rect 2044 6996 2096 7002
rect 2318 6967 2374 6976
rect 2044 6938 2096 6944
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 572 6724 624 6730
rect 572 6666 624 6672
rect 204 3392 256 3398
rect 204 3334 256 3340
rect 216 480 244 3334
rect 584 480 612 6666
rect 1308 6656 1360 6662
rect 1308 6598 1360 6604
rect 1320 3398 1348 6598
rect 1596 6458 1624 6802
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 1308 3392 1360 3398
rect 1308 3334 1360 3340
rect 938 3088 994 3097
rect 938 3023 994 3032
rect 952 480 980 3023
rect 1412 480 1440 6326
rect 2056 6254 2084 6938
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 1490 5808 1546 5817
rect 1490 5743 1546 5752
rect 1504 4078 1532 5743
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1582 4992 1638 5001
rect 1582 4927 1638 4936
rect 1596 4146 1624 4927
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1504 3738 1532 4014
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1688 2650 1716 2926
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1780 480 1808 5510
rect 2332 5234 2360 6967
rect 2516 6866 2544 7375
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2516 6458 2544 6802
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2424 4826 2452 5102
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2320 4752 2372 4758
rect 2320 4694 2372 4700
rect 2332 3738 2360 4694
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1964 3194 1992 3402
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2424 2990 2452 3334
rect 2412 2984 2464 2990
rect 2226 2952 2282 2961
rect 2608 2938 2636 28086
rect 2700 15609 2728 32710
rect 2792 30025 2820 38927
rect 2976 34746 3004 39520
rect 3344 35290 3372 39520
rect 3804 37210 3832 39520
rect 3804 37182 4108 37210
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3422 36952 3478 36961
rect 3622 36944 3918 36964
rect 3422 36887 3478 36896
rect 3436 35737 3464 36887
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3422 35728 3478 35737
rect 3422 35663 3478 35672
rect 3332 35284 3384 35290
rect 3332 35226 3384 35232
rect 3056 35148 3108 35154
rect 3056 35090 3108 35096
rect 2964 34740 3016 34746
rect 2964 34682 3016 34688
rect 3068 34610 3096 35090
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 4080 34626 4108 37182
rect 4172 36825 4200 39520
rect 4158 36816 4214 36825
rect 4158 36751 4214 36760
rect 4250 35320 4306 35329
rect 4250 35255 4252 35264
rect 4304 35255 4306 35264
rect 4252 35226 4304 35232
rect 4252 35148 4304 35154
rect 4252 35090 4304 35096
rect 4264 34785 4292 35090
rect 4250 34776 4306 34785
rect 4250 34711 4252 34720
rect 4304 34711 4306 34720
rect 4252 34682 4304 34688
rect 4540 34649 4568 39520
rect 5000 35834 5028 39520
rect 4988 35828 5040 35834
rect 4988 35770 5040 35776
rect 5172 35148 5224 35154
rect 5172 35090 5224 35096
rect 4526 34640 4582 34649
rect 3056 34604 3108 34610
rect 3056 34546 3108 34552
rect 3332 34604 3384 34610
rect 4080 34598 4200 34626
rect 3332 34546 3384 34552
rect 2964 30592 3016 30598
rect 2964 30534 3016 30540
rect 2976 30190 3004 30534
rect 2964 30184 3016 30190
rect 2964 30126 3016 30132
rect 2778 30016 2834 30025
rect 2778 29951 2834 29960
rect 2780 29844 2832 29850
rect 2780 29786 2832 29792
rect 2792 28762 2820 29786
rect 2872 29708 2924 29714
rect 2872 29650 2924 29656
rect 2884 28966 2912 29650
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 2976 29306 3004 29582
rect 2964 29300 3016 29306
rect 2964 29242 3016 29248
rect 2872 28960 2924 28966
rect 2872 28902 2924 28908
rect 2884 28762 2912 28902
rect 2780 28756 2832 28762
rect 2780 28698 2832 28704
rect 2872 28756 2924 28762
rect 2872 28698 2924 28704
rect 3068 23508 3096 34546
rect 3240 34536 3292 34542
rect 3240 34478 3292 34484
rect 3148 34060 3200 34066
rect 3148 34002 3200 34008
rect 3160 33386 3188 34002
rect 3148 33380 3200 33386
rect 3148 33322 3200 33328
rect 3252 29034 3280 34478
rect 3344 32473 3372 34546
rect 4172 34202 4200 34598
rect 4526 34575 4582 34584
rect 5184 34542 5212 35090
rect 5368 34626 5396 39520
rect 5736 36258 5764 39520
rect 5552 36230 5764 36258
rect 5552 35306 5580 36230
rect 6000 35488 6052 35494
rect 6000 35430 6052 35436
rect 5460 35290 5580 35306
rect 5448 35284 5580 35290
rect 5500 35278 5580 35284
rect 5448 35226 5500 35232
rect 5368 34598 5580 34626
rect 4804 34536 4856 34542
rect 4804 34478 4856 34484
rect 5172 34536 5224 34542
rect 5172 34478 5224 34484
rect 4160 34196 4212 34202
rect 4160 34138 4212 34144
rect 4252 34060 4304 34066
rect 4252 34002 4304 34008
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 4264 33318 4292 34002
rect 4526 33960 4582 33969
rect 4526 33895 4582 33904
rect 4252 33312 4304 33318
rect 4252 33254 4304 33260
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3330 32464 3386 32473
rect 3330 32399 3386 32408
rect 3240 29028 3292 29034
rect 3240 28970 3292 28976
rect 3344 28218 3372 32399
rect 3424 31680 3476 31686
rect 3424 31622 3476 31628
rect 3436 31278 3464 31622
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3424 31272 3476 31278
rect 3424 31214 3476 31220
rect 3436 30190 3464 31214
rect 4160 31136 4212 31142
rect 4160 31078 4212 31084
rect 4068 30592 4120 30598
rect 4068 30534 4120 30540
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3424 30184 3476 30190
rect 3424 30126 3476 30132
rect 3332 28212 3384 28218
rect 3332 28154 3384 28160
rect 3148 24608 3200 24614
rect 3148 24550 3200 24556
rect 3160 24070 3188 24550
rect 3148 24064 3200 24070
rect 3148 24006 3200 24012
rect 3160 23662 3188 24006
rect 3148 23656 3200 23662
rect 3148 23598 3200 23604
rect 3068 23480 3188 23508
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 2780 23248 2832 23254
rect 2780 23190 2832 23196
rect 2792 21962 2820 23190
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 2884 22778 2912 23122
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 2884 22166 2912 22714
rect 2976 22642 3004 23054
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 3068 22574 3096 23258
rect 3056 22568 3108 22574
rect 3056 22510 3108 22516
rect 2964 22432 3016 22438
rect 2964 22374 3016 22380
rect 2976 22234 3004 22374
rect 2964 22228 3016 22234
rect 2964 22170 3016 22176
rect 2872 22160 2924 22166
rect 2872 22102 2924 22108
rect 3160 22114 3188 23480
rect 3344 23338 3372 28154
rect 3436 27130 3464 30126
rect 3516 30116 3568 30122
rect 3516 30058 3568 30064
rect 3528 29510 3556 30058
rect 4080 29850 4108 30534
rect 4068 29844 4120 29850
rect 4068 29786 4120 29792
rect 4172 29646 4200 31078
rect 4160 29640 4212 29646
rect 4160 29582 4212 29588
rect 3516 29504 3568 29510
rect 3516 29446 3568 29452
rect 3528 29170 3556 29446
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 4160 29232 4212 29238
rect 4160 29174 4212 29180
rect 3516 29164 3568 29170
rect 3516 29106 3568 29112
rect 3976 29028 4028 29034
rect 3976 28970 4028 28976
rect 3516 28960 3568 28966
rect 3516 28902 3568 28908
rect 3528 28694 3556 28902
rect 3516 28688 3568 28694
rect 3516 28630 3568 28636
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3700 28076 3752 28082
rect 3700 28018 3752 28024
rect 3712 27674 3740 28018
rect 3700 27668 3752 27674
rect 3700 27610 3752 27616
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3424 27124 3476 27130
rect 3424 27066 3476 27072
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 3516 23588 3568 23594
rect 3516 23530 3568 23536
rect 3344 23310 3464 23338
rect 3436 22681 3464 23310
rect 3422 22672 3478 22681
rect 3528 22642 3556 23530
rect 3896 23186 3924 23598
rect 3884 23180 3936 23186
rect 3884 23122 3936 23128
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3422 22607 3478 22616
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 3252 22234 3280 22510
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3160 22086 3280 22114
rect 2780 21956 2832 21962
rect 2780 21898 2832 21904
rect 3146 20904 3202 20913
rect 2780 20868 2832 20874
rect 3146 20839 3202 20848
rect 2780 20810 2832 20816
rect 2792 19718 2820 20810
rect 2780 19712 2832 19718
rect 2780 19654 2832 19660
rect 2792 19378 2820 19654
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2976 18222 3004 18566
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 3056 18148 3108 18154
rect 3056 18090 3108 18096
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2686 15600 2742 15609
rect 2686 15535 2742 15544
rect 2792 13870 2820 17682
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2884 17338 2912 17614
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2884 16794 2912 17274
rect 2976 17270 3004 17614
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 3068 17202 3096 18090
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13530 2820 13806
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2700 10674 2728 12650
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2700 10266 2728 10610
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2700 8430 2728 9454
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2792 8090 2820 8774
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2792 7546 2820 8026
rect 2884 7954 2912 8230
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2884 4282 2912 4558
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2688 3528 2740 3534
rect 2792 3516 2820 3606
rect 2740 3488 2820 3516
rect 2688 3470 2740 3476
rect 2792 3194 2820 3488
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2412 2926 2464 2932
rect 2226 2887 2228 2896
rect 2280 2887 2282 2896
rect 2516 2910 2636 2938
rect 2228 2858 2280 2864
rect 2410 2680 2466 2689
rect 2410 2615 2412 2624
rect 2464 2615 2466 2624
rect 2412 2586 2464 2592
rect 2134 1456 2190 1465
rect 2134 1391 2190 1400
rect 2148 480 2176 1391
rect 2516 1057 2544 2910
rect 2594 2816 2650 2825
rect 2594 2751 2650 2760
rect 2502 1048 2558 1057
rect 2502 983 2558 992
rect 2608 480 2636 2751
rect 2884 2650 2912 3470
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2976 2514 3004 17070
rect 3068 16794 3096 17138
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 3160 12782 3188 20839
rect 3252 16833 3280 22086
rect 3238 16824 3294 16833
rect 3238 16759 3294 16768
rect 3436 14532 3464 22374
rect 3528 22166 3556 22578
rect 3516 22160 3568 22166
rect 3516 22102 3568 22108
rect 3528 21690 3556 22102
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3988 20913 4016 28970
rect 4172 28762 4200 29174
rect 4160 28756 4212 28762
rect 4160 28698 4212 28704
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 4080 28121 4108 28358
rect 4066 28112 4122 28121
rect 4066 28047 4122 28056
rect 4068 27940 4120 27946
rect 4068 27882 4120 27888
rect 4080 26586 4108 27882
rect 4172 27606 4200 28698
rect 4160 27600 4212 27606
rect 4160 27542 4212 27548
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 4172 26364 4200 26930
rect 4080 26336 4200 26364
rect 4080 25294 4108 26336
rect 4160 25356 4212 25362
rect 4160 25298 4212 25304
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4080 24682 4108 25230
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 4172 24614 4200 25298
rect 4160 24608 4212 24614
rect 4160 24550 4212 24556
rect 4172 23526 4200 24550
rect 4160 23520 4212 23526
rect 4160 23462 4212 23468
rect 4172 23338 4200 23462
rect 4080 23310 4200 23338
rect 4080 23118 4108 23310
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4068 22228 4120 22234
rect 4068 22170 4120 22176
rect 4080 21622 4108 22170
rect 4068 21616 4120 21622
rect 4068 21558 4120 21564
rect 3974 20904 4030 20913
rect 4172 20874 4200 23054
rect 3974 20839 4030 20848
rect 4160 20868 4212 20874
rect 4160 20810 4212 20816
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 4264 19446 4292 33254
rect 4344 31204 4396 31210
rect 4344 31146 4396 31152
rect 4356 30734 4384 31146
rect 4436 30796 4488 30802
rect 4436 30738 4488 30744
rect 4344 30728 4396 30734
rect 4344 30670 4396 30676
rect 4356 30054 4384 30670
rect 4344 30048 4396 30054
rect 4344 29990 4396 29996
rect 4356 29510 4384 29990
rect 4448 29850 4476 30738
rect 4436 29844 4488 29850
rect 4436 29786 4488 29792
rect 4344 29504 4396 29510
rect 4344 29446 4396 29452
rect 4344 29164 4396 29170
rect 4344 29106 4396 29112
rect 4356 28082 4384 29106
rect 4540 28642 4568 33895
rect 4712 33380 4764 33386
rect 4712 33322 4764 33328
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 4448 28614 4568 28642
rect 4344 28076 4396 28082
rect 4344 28018 4396 28024
rect 4448 26382 4476 28614
rect 4632 28558 4660 29446
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 4528 28484 4580 28490
rect 4528 28426 4580 28432
rect 4540 27878 4568 28426
rect 4632 28218 4660 28494
rect 4620 28212 4672 28218
rect 4620 28154 4672 28160
rect 4528 27872 4580 27878
rect 4528 27814 4580 27820
rect 4540 27674 4568 27814
rect 4528 27668 4580 27674
rect 4528 27610 4580 27616
rect 4620 27328 4672 27334
rect 4620 27270 4672 27276
rect 4528 26512 4580 26518
rect 4528 26454 4580 26460
rect 4436 26376 4488 26382
rect 4436 26318 4488 26324
rect 4448 26042 4476 26318
rect 4436 26036 4488 26042
rect 4436 25978 4488 25984
rect 4448 24018 4476 25978
rect 4540 25809 4568 26454
rect 4526 25800 4582 25809
rect 4526 25735 4528 25744
rect 4580 25735 4582 25744
rect 4528 25706 4580 25712
rect 4448 23990 4568 24018
rect 4436 23860 4488 23866
rect 4436 23802 4488 23808
rect 4448 23254 4476 23802
rect 4436 23248 4488 23254
rect 4356 23208 4436 23236
rect 4356 22642 4384 23208
rect 4540 23225 4568 23990
rect 4632 23526 4660 27270
rect 4724 25401 4752 33322
rect 4710 25392 4766 25401
rect 4710 25327 4766 25336
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4436 23190 4488 23196
rect 4526 23216 4582 23225
rect 4526 23151 4582 23160
rect 4724 23066 4752 25327
rect 4816 23322 4844 34478
rect 5552 34202 5580 34598
rect 5724 34536 5776 34542
rect 5724 34478 5776 34484
rect 5540 34196 5592 34202
rect 5540 34138 5592 34144
rect 5172 33312 5224 33318
rect 5172 33254 5224 33260
rect 4986 33144 5042 33153
rect 5184 33114 5212 33254
rect 4986 33079 5042 33088
rect 5172 33108 5224 33114
rect 5000 32570 5028 33079
rect 5172 33050 5224 33056
rect 5184 32570 5212 33050
rect 5540 32904 5592 32910
rect 5540 32846 5592 32852
rect 5448 32768 5500 32774
rect 5448 32710 5500 32716
rect 4988 32564 5040 32570
rect 4988 32506 5040 32512
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 5172 31884 5224 31890
rect 5172 31826 5224 31832
rect 5184 31142 5212 31826
rect 5172 31136 5224 31142
rect 5172 31078 5224 31084
rect 5262 30832 5318 30841
rect 4988 30796 5040 30802
rect 5262 30767 5318 30776
rect 4988 30738 5040 30744
rect 5000 30054 5028 30738
rect 5276 30598 5304 30767
rect 5264 30592 5316 30598
rect 5264 30534 5316 30540
rect 5078 30152 5134 30161
rect 5078 30087 5134 30096
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4988 30048 5040 30054
rect 4988 29990 5040 29996
rect 4908 27334 4936 29990
rect 5000 29782 5028 29990
rect 4988 29776 5040 29782
rect 4988 29718 5040 29724
rect 5092 29646 5120 30087
rect 5276 30054 5304 30534
rect 5356 30252 5408 30258
rect 5356 30194 5408 30200
rect 5264 30048 5316 30054
rect 5264 29990 5316 29996
rect 5172 29776 5224 29782
rect 5172 29718 5224 29724
rect 5080 29640 5132 29646
rect 5080 29582 5132 29588
rect 5092 29306 5120 29582
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 4988 28688 5040 28694
rect 4988 28630 5040 28636
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 4896 26852 4948 26858
rect 4896 26794 4948 26800
rect 4908 26382 4936 26794
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4908 25702 4936 26318
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4908 25498 4936 25638
rect 4896 25492 4948 25498
rect 4896 25434 4948 25440
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4540 23038 4752 23066
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4344 22636 4396 22642
rect 4344 22578 4396 22584
rect 4356 22506 4384 22578
rect 4344 22500 4396 22506
rect 4344 22442 4396 22448
rect 4356 21554 4384 22442
rect 4448 22030 4476 22646
rect 4436 22024 4488 22030
rect 4436 21966 4488 21972
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4448 21146 4476 21966
rect 4436 21140 4488 21146
rect 4436 21082 4488 21088
rect 4540 19496 4568 23038
rect 4816 22964 4844 23258
rect 4724 22936 4844 22964
rect 4896 22976 4948 22982
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4632 21894 4660 22374
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4632 21049 4660 21286
rect 4618 21040 4674 21049
rect 4618 20975 4674 20984
rect 4632 20806 4660 20975
rect 4620 20800 4672 20806
rect 4620 20742 4672 20748
rect 4356 19468 4568 19496
rect 4252 19440 4304 19446
rect 4252 19382 4304 19388
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3988 18222 4016 18702
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3988 17524 4016 18158
rect 4080 18154 4108 19110
rect 4252 18896 4304 18902
rect 4252 18838 4304 18844
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 4172 17898 4200 18294
rect 4264 18086 4292 18838
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4080 17882 4200 17898
rect 4068 17876 4200 17882
rect 4120 17870 4200 17876
rect 4068 17818 4120 17824
rect 4264 17678 4292 18022
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4068 17536 4120 17542
rect 3988 17496 4068 17524
rect 4068 17478 4120 17484
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 4080 16998 4108 17478
rect 4356 17218 4384 19468
rect 4434 19408 4490 19417
rect 4434 19343 4490 19352
rect 4264 17190 4384 17218
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 3620 16794 3648 16934
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3988 16250 4016 16662
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3988 15706 4016 16186
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 4080 15586 4108 16934
rect 4158 16824 4214 16833
rect 4158 16759 4160 16768
rect 4212 16759 4214 16768
rect 4160 16730 4212 16736
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4172 15910 4200 16526
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 3988 15558 4108 15586
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 14822 3556 15302
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3252 14504 3464 14532
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3148 9716 3200 9722
rect 3252 9704 3280 14504
rect 3528 14074 3556 14758
rect 3620 14618 3648 14758
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3884 13864 3936 13870
rect 3988 13852 4016 15558
rect 4172 15178 4200 15846
rect 4264 15570 4292 17190
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4080 15150 4200 15178
rect 4080 15026 4108 15150
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14074 4108 14962
rect 4264 14822 4292 15506
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4172 13870 4200 14282
rect 3936 13824 4016 13852
rect 4160 13864 4212 13870
rect 3884 13806 3936 13812
rect 4160 13806 4212 13812
rect 3896 13258 3924 13806
rect 4172 13530 4200 13806
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 3884 13252 3936 13258
rect 3884 13194 3936 13200
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 4172 12986 4200 13466
rect 4264 13433 4292 14758
rect 4250 13424 4306 13433
rect 4250 13359 4306 13368
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10266 3464 10406
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3200 9676 3280 9704
rect 3148 9658 3200 9664
rect 3068 5896 3096 9658
rect 3884 9648 3936 9654
rect 3882 9616 3884 9625
rect 3936 9616 3938 9625
rect 3882 9551 3938 9560
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 8974 3280 9318
rect 3896 9042 3924 9551
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8498 3280 8910
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3252 8022 3280 8434
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3160 7546 3188 7890
rect 3344 7886 3372 8978
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3988 8401 4016 12718
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4080 10810 4108 11154
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3790 8392 3846 8401
rect 3790 8327 3792 8336
rect 3844 8327 3846 8336
rect 3974 8392 4030 8401
rect 3974 8327 4030 8336
rect 4160 8356 4212 8362
rect 3792 8298 3844 8304
rect 4160 8298 4212 8304
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3344 7478 3372 7822
rect 3436 7750 3464 8230
rect 4068 8084 4120 8090
rect 4172 8072 4200 8298
rect 4120 8044 4200 8072
rect 4068 8026 4120 8032
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3436 7002 3464 7686
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 4080 7313 4108 7686
rect 4066 7304 4122 7313
rect 4066 7239 4122 7248
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3068 5868 3188 5896
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 3068 5302 3096 5714
rect 3056 5296 3108 5302
rect 3054 5264 3056 5273
rect 3108 5264 3110 5273
rect 3054 5199 3110 5208
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 3068 3534 3096 3946
rect 3160 3602 3188 5868
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3436 5166 3464 5510
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3436 4486 3464 5102
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3988 4622 4016 5034
rect 4080 4758 4108 5510
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 3976 4616 4028 4622
rect 3882 4584 3938 4593
rect 3976 4558 4028 4564
rect 3882 4519 3884 4528
rect 3936 4519 3938 4528
rect 3884 4490 3936 4496
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 4298 3464 4422
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3344 4282 3464 4298
rect 3988 4282 4016 4558
rect 4158 4448 4214 4457
rect 4158 4383 4214 4392
rect 3332 4276 3464 4282
rect 3384 4270 3464 4276
rect 3332 4218 3384 4224
rect 3436 3738 3464 4270
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3436 3398 3464 3674
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3884 2576 3936 2582
rect 3882 2544 3884 2553
rect 3936 2544 3938 2553
rect 2964 2508 3016 2514
rect 3882 2479 3938 2488
rect 2964 2450 3016 2456
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2976 480 3004 2314
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3344 480 3372 2246
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3792 2032 3844 2038
rect 3792 1974 3844 1980
rect 3804 480 3832 1974
rect 4172 480 4200 4383
rect 4356 4049 4384 17070
rect 4448 15638 4476 19343
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 17542 4568 19110
rect 4632 17746 4660 20742
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4724 17134 4752 22936
rect 4896 22918 4948 22924
rect 4908 22642 4936 22918
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4908 22166 4936 22578
rect 5000 22506 5028 28630
rect 5092 25702 5120 29242
rect 5184 28762 5212 29718
rect 5172 28756 5224 28762
rect 5172 28698 5224 28704
rect 5276 28642 5304 29990
rect 5368 29594 5396 30194
rect 5460 29714 5488 32710
rect 5552 32502 5580 32846
rect 5540 32496 5592 32502
rect 5540 32438 5592 32444
rect 5552 32026 5580 32438
rect 5630 32328 5686 32337
rect 5630 32263 5686 32272
rect 5644 32230 5672 32263
rect 5632 32224 5684 32230
rect 5632 32166 5684 32172
rect 5540 32020 5592 32026
rect 5540 31962 5592 31968
rect 5632 31952 5684 31958
rect 5632 31894 5684 31900
rect 5644 31482 5672 31894
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 5540 30592 5592 30598
rect 5540 30534 5592 30540
rect 5552 29850 5580 30534
rect 5540 29844 5592 29850
rect 5540 29786 5592 29792
rect 5448 29708 5500 29714
rect 5448 29650 5500 29656
rect 5368 29578 5488 29594
rect 5368 29572 5500 29578
rect 5368 29566 5448 29572
rect 5448 29514 5500 29520
rect 5356 29232 5408 29238
rect 5356 29174 5408 29180
rect 5184 28614 5304 28642
rect 5184 26466 5212 28614
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 5276 27538 5304 28358
rect 5264 27532 5316 27538
rect 5264 27474 5316 27480
rect 5276 27130 5304 27474
rect 5264 27124 5316 27130
rect 5264 27066 5316 27072
rect 5368 26586 5396 29174
rect 5460 29170 5488 29514
rect 5448 29164 5500 29170
rect 5448 29106 5500 29112
rect 5460 28626 5488 29106
rect 5552 29102 5580 29786
rect 5644 29782 5672 30670
rect 5736 30122 5764 34478
rect 5908 32360 5960 32366
rect 5908 32302 5960 32308
rect 5920 32026 5948 32302
rect 5908 32020 5960 32026
rect 5908 31962 5960 31968
rect 5724 30116 5776 30122
rect 5724 30058 5776 30064
rect 5632 29776 5684 29782
rect 5632 29718 5684 29724
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 5644 29170 5672 29582
rect 5816 29504 5868 29510
rect 5816 29446 5868 29452
rect 5828 29170 5856 29446
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 5816 29164 5868 29170
rect 5816 29106 5868 29112
rect 5540 29096 5592 29102
rect 5540 29038 5592 29044
rect 5448 28620 5500 28626
rect 5448 28562 5500 28568
rect 5724 28620 5776 28626
rect 5724 28562 5776 28568
rect 5540 28484 5592 28490
rect 5540 28426 5592 28432
rect 5552 28121 5580 28426
rect 5538 28112 5594 28121
rect 5538 28047 5594 28056
rect 5632 28076 5684 28082
rect 5552 28014 5580 28047
rect 5632 28018 5684 28024
rect 5540 28008 5592 28014
rect 5540 27950 5592 27956
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 5356 26580 5408 26586
rect 5356 26522 5408 26528
rect 5184 26438 5396 26466
rect 5080 25696 5132 25702
rect 5080 25638 5132 25644
rect 5264 24744 5316 24750
rect 5264 24686 5316 24692
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 5092 22234 5120 24550
rect 5184 24410 5212 24550
rect 5172 24404 5224 24410
rect 5172 24346 5224 24352
rect 5184 23730 5212 24346
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5080 22228 5132 22234
rect 5080 22170 5132 22176
rect 4896 22160 4948 22166
rect 5184 22114 5212 23462
rect 4896 22102 4948 22108
rect 5092 22086 5212 22114
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 4816 21690 4844 21830
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4804 19440 4856 19446
rect 4804 19382 4856 19388
rect 4816 18902 4844 19382
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 5000 18970 5028 19110
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 4804 18896 4856 18902
rect 4804 18838 4856 18844
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4632 16561 4660 16730
rect 4618 16552 4674 16561
rect 4528 16516 4580 16522
rect 4618 16487 4674 16496
rect 4528 16458 4580 16464
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 4540 14482 4568 16458
rect 4632 16250 4660 16487
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4712 15632 4764 15638
rect 4712 15574 4764 15580
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4448 14385 4476 14418
rect 4434 14376 4490 14385
rect 4434 14311 4490 14320
rect 4448 13462 4476 14311
rect 4540 13977 4568 14418
rect 4632 14414 4660 15438
rect 4724 14822 4752 15574
rect 4816 15026 4844 18838
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4526 13968 4582 13977
rect 4526 13903 4582 13912
rect 4540 13802 4568 13903
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4436 13456 4488 13462
rect 4436 13398 4488 13404
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4632 12918 4660 13262
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4632 12442 4660 12854
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4724 12322 4752 14758
rect 4908 12481 4936 17614
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 17202 5028 17478
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 5000 16590 5028 17138
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4894 12472 4950 12481
rect 5092 12442 5120 22086
rect 5170 21448 5226 21457
rect 5170 21383 5172 21392
rect 5224 21383 5226 21392
rect 5172 21354 5224 21360
rect 5276 19802 5304 24686
rect 5368 24596 5396 26438
rect 5460 25786 5488 27814
rect 5644 27674 5672 28018
rect 5632 27668 5684 27674
rect 5632 27610 5684 27616
rect 5736 27130 5764 28562
rect 5828 28082 5856 29106
rect 6012 29034 6040 35430
rect 6196 34746 6224 39520
rect 6564 37754 6592 39520
rect 6564 37726 6684 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6656 35290 6684 37726
rect 6932 35834 6960 39520
rect 7286 36816 7342 36825
rect 7286 36751 7342 36760
rect 7300 36378 7328 36751
rect 7288 36372 7340 36378
rect 7288 36314 7340 36320
rect 7196 36236 7248 36242
rect 7196 36178 7248 36184
rect 6920 35828 6972 35834
rect 6920 35770 6972 35776
rect 7208 35494 7236 36178
rect 7288 35624 7340 35630
rect 7288 35566 7340 35572
rect 7196 35488 7248 35494
rect 7196 35430 7248 35436
rect 6644 35284 6696 35290
rect 6644 35226 6696 35232
rect 6828 35148 6880 35154
rect 6828 35090 6880 35096
rect 6184 34740 6236 34746
rect 6184 34682 6236 34688
rect 6840 34542 6868 35090
rect 7300 34950 7328 35566
rect 7392 35290 7420 39520
rect 7380 35284 7432 35290
rect 7380 35226 7432 35232
rect 7472 35148 7524 35154
rect 7472 35090 7524 35096
rect 7288 34944 7340 34950
rect 7288 34886 7340 34892
rect 7102 34776 7158 34785
rect 7102 34711 7158 34720
rect 6828 34536 6880 34542
rect 6828 34478 6880 34484
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6092 34060 6144 34066
rect 6092 34002 6144 34008
rect 6104 33318 6132 34002
rect 6092 33312 6144 33318
rect 6092 33254 6144 33260
rect 6000 29028 6052 29034
rect 6000 28970 6052 28976
rect 5908 28620 5960 28626
rect 5908 28562 5960 28568
rect 5816 28076 5868 28082
rect 5816 28018 5868 28024
rect 5920 27130 5948 28562
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 5908 27124 5960 27130
rect 5908 27066 5960 27072
rect 6012 27010 6040 28970
rect 5920 26982 6040 27010
rect 5920 26976 5948 26982
rect 5736 26948 5948 26976
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5552 25906 5580 26318
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 5644 25838 5672 26522
rect 5632 25832 5684 25838
rect 5460 25770 5580 25786
rect 5632 25774 5684 25780
rect 5460 25764 5592 25770
rect 5460 25758 5540 25764
rect 5540 25706 5592 25712
rect 5552 25498 5580 25706
rect 5632 25696 5684 25702
rect 5632 25638 5684 25644
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5448 24744 5500 24750
rect 5446 24712 5448 24721
rect 5500 24712 5502 24721
rect 5446 24647 5502 24656
rect 5368 24568 5488 24596
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 5368 22778 5396 24006
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5354 22128 5410 22137
rect 5460 22114 5488 24568
rect 5644 23662 5672 25638
rect 5632 23656 5684 23662
rect 5632 23598 5684 23604
rect 5736 23508 5764 26948
rect 6000 26920 6052 26926
rect 6000 26862 6052 26868
rect 6104 26874 6132 33254
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6550 33008 6606 33017
rect 6550 32943 6606 32952
rect 6564 32570 6592 32943
rect 6644 32904 6696 32910
rect 6644 32846 6696 32852
rect 6184 32564 6236 32570
rect 6184 32506 6236 32512
rect 6552 32564 6604 32570
rect 6552 32506 6604 32512
rect 6196 26994 6224 32506
rect 6564 32298 6592 32506
rect 6552 32292 6604 32298
rect 6552 32234 6604 32240
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6656 31906 6684 32846
rect 6736 32292 6788 32298
rect 6736 32234 6788 32240
rect 6564 31890 6684 31906
rect 6552 31884 6684 31890
rect 6604 31878 6684 31884
rect 6552 31826 6604 31832
rect 6564 31482 6592 31826
rect 6552 31476 6604 31482
rect 6552 31418 6604 31424
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6644 30592 6696 30598
rect 6644 30534 6696 30540
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6656 29850 6684 30534
rect 6644 29844 6696 29850
rect 6644 29786 6696 29792
rect 6276 29708 6328 29714
rect 6276 29650 6328 29656
rect 6288 29034 6316 29650
rect 6276 29028 6328 29034
rect 6276 28970 6328 28976
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6656 28762 6684 29786
rect 6748 29073 6776 32234
rect 6734 29064 6790 29073
rect 6734 28999 6790 29008
rect 6644 28756 6696 28762
rect 6644 28698 6696 28704
rect 6748 28234 6776 28999
rect 6656 28206 6776 28234
rect 6840 28218 6868 34478
rect 6920 32972 6972 32978
rect 6920 32914 6972 32920
rect 6932 32502 6960 32914
rect 7012 32768 7064 32774
rect 7012 32710 7064 32716
rect 6920 32496 6972 32502
rect 6920 32438 6972 32444
rect 6920 32360 6972 32366
rect 6920 32302 6972 32308
rect 6932 32026 6960 32302
rect 6920 32020 6972 32026
rect 6920 31962 6972 31968
rect 6920 31136 6972 31142
rect 6920 31078 6972 31084
rect 6932 30705 6960 31078
rect 6918 30696 6974 30705
rect 6918 30631 6974 30640
rect 7024 29646 7052 32710
rect 7116 30802 7144 34711
rect 7196 31952 7248 31958
rect 7196 31894 7248 31900
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 7208 30734 7236 31894
rect 7300 31362 7328 34886
rect 7484 34746 7512 35090
rect 7472 34740 7524 34746
rect 7472 34682 7524 34688
rect 7378 34640 7434 34649
rect 7378 34575 7434 34584
rect 7392 33658 7420 34575
rect 7760 34202 7788 39520
rect 8220 35578 8248 39520
rect 7944 35550 8248 35578
rect 7838 34640 7894 34649
rect 7838 34575 7894 34584
rect 7852 34542 7880 34575
rect 7840 34536 7892 34542
rect 7840 34478 7892 34484
rect 7748 34196 7800 34202
rect 7748 34138 7800 34144
rect 7840 34060 7892 34066
rect 7840 34002 7892 34008
rect 7852 33658 7880 34002
rect 7380 33652 7432 33658
rect 7380 33594 7432 33600
rect 7840 33652 7892 33658
rect 7840 33594 7892 33600
rect 7852 33561 7880 33594
rect 7838 33552 7894 33561
rect 7838 33487 7894 33496
rect 7748 33448 7800 33454
rect 7748 33390 7800 33396
rect 7760 33289 7788 33390
rect 7746 33280 7802 33289
rect 7746 33215 7802 33224
rect 7944 32366 7972 35550
rect 8208 35488 8260 35494
rect 8208 35430 8260 35436
rect 8116 34944 8168 34950
rect 8116 34886 8168 34892
rect 8220 34898 8248 35430
rect 8128 34542 8156 34886
rect 8220 34870 8432 34898
rect 8208 34740 8260 34746
rect 8208 34682 8260 34688
rect 8220 34626 8248 34682
rect 8220 34598 8340 34626
rect 8116 34536 8168 34542
rect 8116 34478 8168 34484
rect 8024 34468 8076 34474
rect 8024 34410 8076 34416
rect 7932 32360 7984 32366
rect 7932 32302 7984 32308
rect 7380 32224 7432 32230
rect 7380 32166 7432 32172
rect 7392 31890 7420 32166
rect 7472 31952 7524 31958
rect 7472 31894 7524 31900
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 7484 31482 7512 31894
rect 7472 31476 7524 31482
rect 7472 31418 7524 31424
rect 7300 31334 7604 31362
rect 7286 30968 7342 30977
rect 7286 30903 7288 30912
rect 7340 30903 7342 30912
rect 7288 30874 7340 30880
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 7208 30394 7236 30670
rect 7196 30388 7248 30394
rect 7196 30330 7248 30336
rect 7300 30258 7328 30874
rect 7380 30796 7432 30802
rect 7380 30738 7432 30744
rect 7104 30252 7156 30258
rect 7104 30194 7156 30200
rect 7288 30252 7340 30258
rect 7288 30194 7340 30200
rect 7012 29640 7064 29646
rect 7012 29582 7064 29588
rect 7024 29306 7052 29582
rect 7012 29300 7064 29306
rect 7012 29242 7064 29248
rect 6920 28960 6972 28966
rect 6920 28902 6972 28908
rect 6932 28422 6960 28902
rect 7024 28762 7052 29242
rect 7012 28756 7064 28762
rect 7012 28698 7064 28704
rect 7024 28558 7052 28698
rect 7116 28694 7144 30194
rect 7392 30054 7420 30738
rect 7380 30048 7432 30054
rect 7380 29990 7432 29996
rect 7104 28688 7156 28694
rect 7104 28630 7156 28636
rect 7012 28552 7064 28558
rect 7012 28494 7064 28500
rect 6920 28416 6972 28422
rect 6920 28358 6972 28364
rect 6828 28212 6880 28218
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6656 27554 6684 28206
rect 6828 28154 6880 28160
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 6564 27526 6684 27554
rect 6184 26988 6236 26994
rect 6184 26930 6236 26936
rect 5816 26852 5868 26858
rect 5816 26794 5868 26800
rect 5828 23746 5856 26794
rect 5908 26376 5960 26382
rect 5908 26318 5960 26324
rect 5920 25158 5948 26318
rect 5908 25152 5960 25158
rect 5908 25094 5960 25100
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5920 24206 5948 24754
rect 6012 24410 6040 26862
rect 6104 26846 6224 26874
rect 6564 26858 6592 27526
rect 6748 27334 6776 28018
rect 7024 27962 7052 28494
rect 6840 27934 7052 27962
rect 6840 27538 6868 27934
rect 7104 27668 7156 27674
rect 7104 27610 7156 27616
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6736 27328 6788 27334
rect 6736 27270 6788 27276
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6000 24404 6052 24410
rect 6000 24346 6052 24352
rect 6012 24313 6040 24346
rect 5998 24304 6054 24313
rect 5998 24239 6054 24248
rect 6092 24268 6144 24274
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 5920 23866 5948 24142
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 6012 23798 6040 24239
rect 6092 24210 6144 24216
rect 6000 23792 6052 23798
rect 5828 23718 5948 23746
rect 6000 23734 6052 23740
rect 5644 23480 5764 23508
rect 5644 22114 5672 23480
rect 5410 22086 5488 22114
rect 5552 22086 5672 22114
rect 5816 22092 5868 22098
rect 5354 22063 5410 22072
rect 5184 19774 5304 19802
rect 5184 19242 5212 19774
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 5184 17678 5212 19178
rect 5276 19174 5304 19654
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5276 17882 5304 19110
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5170 17232 5226 17241
rect 5368 17218 5396 22063
rect 5552 22012 5580 22086
rect 5816 22034 5868 22040
rect 5724 22024 5776 22030
rect 5552 21984 5672 22012
rect 5446 21584 5502 21593
rect 5446 21519 5448 21528
rect 5500 21519 5502 21528
rect 5448 21490 5500 21496
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5552 20942 5580 21422
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5460 18222 5488 18906
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5460 17746 5488 18022
rect 5552 17814 5580 18566
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5460 17338 5488 17682
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5170 17167 5226 17176
rect 5276 17190 5396 17218
rect 5184 17134 5212 17167
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5184 15706 5212 15982
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 14618 5212 14758
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5184 13462 5212 14418
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 5184 12986 5212 13398
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4894 12407 4950 12416
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4988 12368 5040 12374
rect 4448 12294 4752 12322
rect 4894 12336 4950 12345
rect 4448 6440 4476 12294
rect 4988 12310 5040 12316
rect 4894 12271 4950 12280
rect 4802 11520 4858 11529
rect 4802 11455 4858 11464
rect 4816 11354 4844 11455
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4724 10810 4752 11086
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4540 9722 4568 9998
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4632 9654 4660 9998
rect 4724 9761 4752 10746
rect 4710 9752 4766 9761
rect 4710 9687 4766 9696
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8838 4568 8910
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 8634 4568 8774
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4448 6412 4568 6440
rect 4436 6248 4488 6254
rect 4434 6216 4436 6225
rect 4488 6216 4490 6225
rect 4434 6151 4490 6160
rect 4540 5273 4568 6412
rect 4526 5264 4582 5273
rect 4526 5199 4582 5208
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4540 4146 4568 4626
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4342 4040 4398 4049
rect 4342 3975 4398 3984
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4264 2825 4292 3334
rect 4250 2816 4306 2825
rect 4250 2751 4306 2760
rect 4356 2650 4384 3538
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4448 3126 4476 3402
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4540 480 4568 3946
rect 4632 2972 4660 9318
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8362 4844 8910
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4724 3126 4752 6190
rect 4816 5370 4844 8298
rect 4908 6848 4936 12271
rect 5000 11558 5028 12310
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5092 11898 5120 12242
rect 5184 12102 5212 12922
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5000 9382 5028 11494
rect 5092 9994 5120 11834
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8022 5028 8978
rect 4988 8016 5040 8022
rect 4986 7984 4988 7993
rect 5040 7984 5042 7993
rect 4986 7919 5042 7928
rect 5000 7449 5028 7919
rect 5092 7546 5120 9930
rect 5276 9450 5304 17190
rect 5552 16998 5580 17750
rect 5644 17649 5672 21984
rect 5724 21966 5776 21972
rect 5736 20874 5764 21966
rect 5828 21332 5856 22034
rect 5920 21486 5948 23718
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 5908 21480 5960 21486
rect 5908 21422 5960 21428
rect 5908 21344 5960 21350
rect 5828 21304 5908 21332
rect 5908 21286 5960 21292
rect 5724 20868 5776 20874
rect 5724 20810 5776 20816
rect 5920 20602 5948 21286
rect 5908 20596 5960 20602
rect 5908 20538 5960 20544
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5630 17640 5686 17649
rect 5630 17575 5686 17584
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5552 16266 5580 16934
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5368 16238 5580 16266
rect 5368 15978 5396 16238
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5368 15434 5396 15914
rect 5644 15910 5672 16390
rect 5736 16114 5764 16730
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5460 15314 5488 15846
rect 5632 15360 5684 15366
rect 5460 15286 5580 15314
rect 5632 15302 5684 15308
rect 5552 14550 5580 15286
rect 5644 14822 5672 15302
rect 5736 15026 5764 16050
rect 5828 15858 5856 20266
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5920 16590 5948 20198
rect 6012 17218 6040 23598
rect 6104 23594 6132 24210
rect 6092 23588 6144 23594
rect 6092 23530 6144 23536
rect 6104 21146 6132 23530
rect 6196 23236 6224 26846
rect 6552 26852 6604 26858
rect 6552 26794 6604 26800
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6276 26512 6328 26518
rect 6276 26454 6328 26460
rect 6288 26042 6316 26454
rect 6656 26042 6684 27066
rect 6748 26518 6776 27270
rect 6840 27130 6868 27474
rect 6828 27124 6880 27130
rect 6828 27066 6880 27072
rect 6826 27024 6882 27033
rect 6826 26959 6882 26968
rect 6840 26926 6868 26959
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6736 26512 6788 26518
rect 6736 26454 6788 26460
rect 7116 26042 7144 27610
rect 7196 27532 7248 27538
rect 7196 27474 7248 27480
rect 7208 26246 7236 27474
rect 7288 26784 7340 26790
rect 7288 26726 7340 26732
rect 7300 26314 7328 26726
rect 7288 26308 7340 26314
rect 7288 26250 7340 26256
rect 7196 26240 7248 26246
rect 7196 26182 7248 26188
rect 6276 26036 6328 26042
rect 6276 25978 6328 25984
rect 6644 26036 6696 26042
rect 6644 25978 6696 25984
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6656 25362 6684 25978
rect 6644 25356 6696 25362
rect 6644 25298 6696 25304
rect 6656 24954 6684 25298
rect 7208 25158 7236 26182
rect 7288 26036 7340 26042
rect 7288 25978 7340 25984
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 6644 24948 6696 24954
rect 6644 24890 6696 24896
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6748 24070 6776 25094
rect 7208 24886 7236 25094
rect 7196 24880 7248 24886
rect 7102 24848 7158 24857
rect 7196 24822 7248 24828
rect 7102 24783 7158 24792
rect 6920 24744 6972 24750
rect 6840 24692 6920 24698
rect 6840 24686 6972 24692
rect 6840 24670 6960 24686
rect 7012 24676 7064 24682
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6644 23656 6696 23662
rect 6644 23598 6696 23604
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6196 23208 6316 23236
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6196 22778 6224 23054
rect 6184 22772 6236 22778
rect 6184 22714 6236 22720
rect 6182 22672 6238 22681
rect 6288 22658 6316 23208
rect 6656 23050 6684 23598
rect 6644 23044 6696 23050
rect 6644 22986 6696 22992
rect 6656 22778 6684 22986
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6288 22630 6684 22658
rect 6182 22607 6238 22616
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 6104 20262 6132 20878
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6012 17190 6132 17218
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5920 16046 5948 16390
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 6000 15904 6052 15910
rect 5828 15830 5948 15858
rect 6000 15846 6052 15852
rect 5920 15745 5948 15830
rect 5906 15736 5962 15745
rect 5816 15700 5868 15706
rect 5906 15671 5962 15680
rect 5816 15642 5868 15648
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5736 14482 5764 14962
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5828 14414 5856 15642
rect 5908 15632 5960 15638
rect 5906 15600 5908 15609
rect 5960 15600 5962 15609
rect 5906 15535 5962 15544
rect 5920 15094 5948 15535
rect 6012 15162 6040 15846
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 5908 15088 5960 15094
rect 5908 15030 5960 15036
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5538 12608 5594 12617
rect 5538 12543 5594 12552
rect 5552 12442 5580 12543
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5644 11370 5672 14214
rect 5828 13841 5856 14350
rect 5814 13832 5870 13841
rect 5814 13767 5870 13776
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5828 13190 5856 13670
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5814 12200 5870 12209
rect 5814 12135 5870 12144
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5736 11762 5764 12038
rect 5828 11830 5856 12135
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5460 11342 5672 11370
rect 5460 11286 5488 11342
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10810 5580 11018
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5736 10674 5764 11698
rect 5828 11694 5856 11766
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 10266 5580 10406
rect 5540 10260 5592 10266
rect 5828 10248 5856 11630
rect 5540 10202 5592 10208
rect 5644 10220 5856 10248
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5460 10010 5488 10066
rect 5460 9982 5580 10010
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5368 8945 5396 9318
rect 5354 8936 5410 8945
rect 5460 8906 5488 9522
rect 5552 9178 5580 9982
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5354 8871 5410 8880
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5460 8634 5488 8842
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5368 7886 5396 8366
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5552 8090 5580 8298
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 4986 7440 5042 7449
rect 4986 7375 5042 7384
rect 5368 7290 5396 7822
rect 5460 7546 5488 7890
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5368 7262 5488 7290
rect 5460 7206 5488 7262
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5080 6860 5132 6866
rect 4908 6820 5028 6848
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4802 4040 4858 4049
rect 4802 3975 4858 3984
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4632 2944 4752 2972
rect 4618 2816 4674 2825
rect 4618 2751 4674 2760
rect 4632 2650 4660 2751
rect 4724 2689 4752 2944
rect 4816 2825 4844 3975
rect 4802 2816 4858 2825
rect 4908 2802 4936 6666
rect 5000 6458 5028 6820
rect 5080 6802 5132 6808
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 5000 6254 5028 6394
rect 4988 6248 5040 6254
rect 5092 6225 5120 6802
rect 5460 6662 5488 7142
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5538 6624 5594 6633
rect 4988 6190 5040 6196
rect 5078 6216 5134 6225
rect 5078 6151 5134 6160
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5092 4593 5120 5714
rect 5172 5704 5224 5710
rect 5276 5681 5304 6598
rect 5538 6559 5594 6568
rect 5552 6458 5580 6559
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5552 6254 5580 6394
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5172 5646 5224 5652
rect 5262 5672 5318 5681
rect 5078 4584 5134 4593
rect 5078 4519 5134 4528
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5000 3738 5028 3878
rect 5092 3738 5120 4519
rect 5184 4282 5212 5646
rect 5552 5658 5580 6054
rect 5262 5607 5318 5616
rect 5368 5630 5580 5658
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5276 5370 5304 5510
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5276 4826 5304 5306
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5276 4214 5304 4762
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 2990 5028 3334
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4908 2774 5028 2802
rect 4802 2751 4858 2760
rect 4710 2680 4766 2689
rect 4620 2644 4672 2650
rect 4710 2615 4766 2624
rect 4620 2586 4672 2592
rect 5000 480 5028 2774
rect 5368 480 5396 5630
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 4010 5488 5510
rect 5644 5370 5672 10220
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5828 9489 5856 10066
rect 5814 9480 5870 9489
rect 5814 9415 5870 9424
rect 5828 8634 5856 9415
rect 5920 8838 5948 14826
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 14074 6040 14758
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6104 13546 6132 17190
rect 6196 16726 6224 22607
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6656 21729 6684 22630
rect 6748 22166 6776 24006
rect 6840 23322 6868 24670
rect 7012 24618 7064 24624
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6932 23594 6960 24006
rect 7024 23866 7052 24618
rect 7116 24614 7144 24783
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 7208 23662 7236 24210
rect 7196 23656 7248 23662
rect 7196 23598 7248 23604
rect 6920 23588 6972 23594
rect 6920 23530 6972 23536
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 6840 22574 6868 23122
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6932 22522 6960 23054
rect 7208 22710 7236 23054
rect 7196 22704 7248 22710
rect 7194 22672 7196 22681
rect 7248 22672 7250 22681
rect 7194 22607 7250 22616
rect 6840 22386 6868 22510
rect 6932 22494 7052 22522
rect 6840 22358 6960 22386
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6642 21720 6698 21729
rect 6932 21690 6960 22358
rect 6642 21655 6698 21664
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6472 20330 6500 20946
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6748 20602 6776 20878
rect 7024 20874 7052 22494
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7116 21593 7144 21830
rect 7102 21584 7158 21593
rect 7102 21519 7158 21528
rect 6828 20868 6880 20874
rect 6828 20810 6880 20816
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6840 20466 6868 20810
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6460 20324 6512 20330
rect 6460 20266 6512 20272
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6840 20058 6868 20402
rect 6920 20324 6972 20330
rect 6920 20266 6972 20272
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6932 19718 6960 20266
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6748 18873 6776 18906
rect 6734 18864 6790 18873
rect 6734 18799 6790 18808
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6656 18426 6684 18634
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6840 18222 6868 19110
rect 6932 18698 6960 19654
rect 7300 19281 7328 25978
rect 7392 24596 7420 29990
rect 7472 28960 7524 28966
rect 7472 28902 7524 28908
rect 7484 28694 7512 28902
rect 7576 28801 7604 31334
rect 7840 30592 7892 30598
rect 7840 30534 7892 30540
rect 7748 30116 7800 30122
rect 7748 30058 7800 30064
rect 7760 29850 7788 30058
rect 7852 30054 7880 30534
rect 7840 30048 7892 30054
rect 7840 29990 7892 29996
rect 7748 29844 7800 29850
rect 7748 29786 7800 29792
rect 7562 28792 7618 28801
rect 7562 28727 7618 28736
rect 7472 28688 7524 28694
rect 7472 28630 7524 28636
rect 7562 28656 7618 28665
rect 7484 28218 7512 28630
rect 7562 28591 7564 28600
rect 7616 28591 7618 28600
rect 7564 28562 7616 28568
rect 7472 28212 7524 28218
rect 7472 28154 7524 28160
rect 7470 28112 7526 28121
rect 7470 28047 7472 28056
rect 7524 28047 7526 28056
rect 7472 28018 7524 28024
rect 7484 27674 7512 28018
rect 7576 27946 7604 28562
rect 7748 28552 7800 28558
rect 7748 28494 7800 28500
rect 7760 28082 7788 28494
rect 7748 28076 7800 28082
rect 7748 28018 7800 28024
rect 7564 27940 7616 27946
rect 7564 27882 7616 27888
rect 7472 27668 7524 27674
rect 7472 27610 7524 27616
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7484 26450 7512 26862
rect 7472 26444 7524 26450
rect 7472 26386 7524 26392
rect 7576 26042 7604 27270
rect 7852 26489 7880 29990
rect 7944 28558 7972 32302
rect 8036 31346 8064 34410
rect 8128 33300 8156 34478
rect 8128 33272 8248 33300
rect 8220 32042 8248 33272
rect 8312 32570 8340 34598
rect 8300 32564 8352 32570
rect 8300 32506 8352 32512
rect 8220 32026 8340 32042
rect 8220 32020 8352 32026
rect 8220 32014 8300 32020
rect 8024 31340 8076 31346
rect 8024 31282 8076 31288
rect 8024 31204 8076 31210
rect 8024 31146 8076 31152
rect 8036 29850 8064 31146
rect 8116 31136 8168 31142
rect 8116 31078 8168 31084
rect 8128 30938 8156 31078
rect 8116 30932 8168 30938
rect 8116 30874 8168 30880
rect 8128 30394 8156 30874
rect 8116 30388 8168 30394
rect 8116 30330 8168 30336
rect 8220 30258 8248 32014
rect 8300 31962 8352 31968
rect 8404 30258 8432 34870
rect 8588 33658 8616 39520
rect 8956 37210 8984 39520
rect 8772 37182 8984 37210
rect 8576 33652 8628 33658
rect 8576 33594 8628 33600
rect 8588 33538 8616 33594
rect 8496 33510 8616 33538
rect 8208 30252 8260 30258
rect 8208 30194 8260 30200
rect 8392 30252 8444 30258
rect 8392 30194 8444 30200
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 8220 29646 8248 30194
rect 8300 29844 8352 29850
rect 8300 29786 8352 29792
rect 8208 29640 8260 29646
rect 8208 29582 8260 29588
rect 8220 29306 8248 29582
rect 8208 29300 8260 29306
rect 8208 29242 8260 29248
rect 8312 28914 8340 29786
rect 8220 28886 8340 28914
rect 8392 28960 8444 28966
rect 8392 28902 8444 28908
rect 8220 28762 8248 28886
rect 8208 28756 8260 28762
rect 8208 28698 8260 28704
rect 7932 28552 7984 28558
rect 7932 28494 7984 28500
rect 7838 26480 7894 26489
rect 7838 26415 7894 26424
rect 7564 26036 7616 26042
rect 7564 25978 7616 25984
rect 7576 25673 7604 25978
rect 7656 25696 7708 25702
rect 7562 25664 7618 25673
rect 7656 25638 7708 25644
rect 7562 25599 7618 25608
rect 7472 25152 7524 25158
rect 7472 25094 7524 25100
rect 7484 24750 7512 25094
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7392 24568 7512 24596
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7392 22166 7420 22510
rect 7380 22160 7432 22166
rect 7380 22102 7432 22108
rect 7380 21480 7432 21486
rect 7484 21457 7512 24568
rect 7562 23352 7618 23361
rect 7562 23287 7564 23296
rect 7616 23287 7618 23296
rect 7564 23258 7616 23264
rect 7576 22506 7604 23258
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7576 21554 7604 22442
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7380 21422 7432 21428
rect 7470 21448 7526 21457
rect 7392 21146 7420 21422
rect 7470 21383 7526 21392
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7286 19272 7342 19281
rect 7286 19207 7342 19216
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6748 16794 6776 17478
rect 6840 17066 6868 18158
rect 7116 17882 7144 18770
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7208 18426 7236 18702
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7104 17604 7156 17610
rect 7104 17546 7156 17552
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6828 17060 6880 17066
rect 6828 17002 6880 17008
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6196 16250 6224 16662
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6182 16008 6238 16017
rect 6288 15978 6316 16594
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6182 15943 6238 15952
rect 6276 15972 6328 15978
rect 6196 15706 6224 15943
rect 6276 15914 6328 15920
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6182 15600 6238 15609
rect 6182 15535 6238 15544
rect 6196 14521 6224 15535
rect 6656 15502 6684 16526
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6368 14544 6420 14550
rect 6182 14512 6238 14521
rect 6368 14486 6420 14492
rect 6182 14447 6238 14456
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13734 6224 14350
rect 6380 14074 6408 14486
rect 6748 14414 6776 16186
rect 6826 15872 6882 15881
rect 6826 15807 6882 15816
rect 6840 15706 6868 15807
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6828 15496 6880 15502
rect 6880 15444 6960 15450
rect 6828 15438 6960 15444
rect 6840 15422 6960 15438
rect 6932 15026 6960 15422
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6734 13696 6790 13705
rect 6289 13628 6585 13648
rect 6734 13631 6790 13640
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6104 13518 6224 13546
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11694 6040 12038
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5998 11112 6054 11121
rect 5998 11047 6054 11056
rect 6012 9178 6040 11047
rect 6104 10470 6132 13126
rect 6196 10606 6224 13518
rect 6748 13394 6776 13631
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6840 13274 6868 14962
rect 7024 14770 7052 17070
rect 7116 16946 7144 17546
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17066 7236 17478
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7116 16918 7236 16946
rect 7208 15978 7236 16918
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15638 7144 15846
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7208 15065 7236 15914
rect 7300 15502 7328 19207
rect 7484 16640 7512 21383
rect 7576 21078 7604 21490
rect 7564 21072 7616 21078
rect 7564 21014 7616 21020
rect 7668 19417 7696 25638
rect 7944 25106 7972 28494
rect 8116 28416 8168 28422
rect 8116 28358 8168 28364
rect 8128 28150 8156 28358
rect 8116 28144 8168 28150
rect 8116 28086 8168 28092
rect 7852 25078 7972 25106
rect 7748 21344 7800 21350
rect 7746 21312 7748 21321
rect 7800 21312 7802 21321
rect 7746 21247 7802 21256
rect 7852 21146 7880 25078
rect 7932 23792 7984 23798
rect 7932 23734 7984 23740
rect 7944 23254 7972 23734
rect 8024 23588 8076 23594
rect 8024 23530 8076 23536
rect 8036 23322 8064 23530
rect 8024 23316 8076 23322
rect 8024 23258 8076 23264
rect 7932 23248 7984 23254
rect 7932 23190 7984 23196
rect 8022 23216 8078 23225
rect 8022 23151 8078 23160
rect 8128 23168 8156 28086
rect 8404 28014 8432 28902
rect 8208 28008 8260 28014
rect 8206 27976 8208 27985
rect 8392 28008 8444 28014
rect 8260 27976 8262 27985
rect 8392 27950 8444 27956
rect 8206 27911 8262 27920
rect 8496 25809 8524 33510
rect 8576 32428 8628 32434
rect 8576 32370 8628 32376
rect 8588 31958 8616 32370
rect 8772 32337 8800 37182
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 9310 33960 9366 33969
rect 9310 33895 9366 33904
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9324 33658 9352 33895
rect 9416 33810 9444 39520
rect 9680 34060 9732 34066
rect 9680 34002 9732 34008
rect 9416 33782 9628 33810
rect 9312 33652 9364 33658
rect 9312 33594 9364 33600
rect 9324 33386 9352 33594
rect 9312 33380 9364 33386
rect 9312 33322 9364 33328
rect 9496 33312 9548 33318
rect 9496 33254 9548 33260
rect 9402 33144 9458 33153
rect 9508 33114 9536 33254
rect 9402 33079 9458 33088
rect 9496 33108 9548 33114
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 9324 32366 9352 32710
rect 9312 32360 9364 32366
rect 8758 32328 8814 32337
rect 8668 32292 8720 32298
rect 8758 32263 8814 32272
rect 9310 32328 9312 32337
rect 9364 32328 9366 32337
rect 9310 32263 9366 32272
rect 8668 32234 8720 32240
rect 8576 31952 8628 31958
rect 8576 31894 8628 31900
rect 8588 30326 8616 31894
rect 8576 30320 8628 30326
rect 8576 30262 8628 30268
rect 8576 29776 8628 29782
rect 8576 29718 8628 29724
rect 8588 28762 8616 29718
rect 8576 28756 8628 28762
rect 8576 28698 8628 28704
rect 8482 25800 8538 25809
rect 8482 25735 8538 25744
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8312 24410 8340 24754
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8208 23724 8260 23730
rect 8260 23684 8340 23712
rect 8208 23666 8260 23672
rect 8208 23180 8260 23186
rect 8036 22574 8064 23151
rect 8128 23140 8208 23168
rect 8208 23122 8260 23128
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7654 19408 7710 19417
rect 7654 19343 7710 19352
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7576 19145 7604 19178
rect 7562 19136 7618 19145
rect 7562 19071 7618 19080
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7392 16612 7512 16640
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7194 15056 7250 15065
rect 7194 14991 7250 15000
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7194 14784 7250 14793
rect 7024 14742 7144 14770
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7024 14074 7052 14554
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7116 13394 7144 14742
rect 7194 14719 7250 14728
rect 7208 13802 7236 14719
rect 7300 14618 7328 14962
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7392 13954 7420 16612
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 7484 16046 7512 16458
rect 7654 16144 7710 16153
rect 7760 16114 7788 17002
rect 7852 16794 7880 18362
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7944 17066 7972 17682
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7654 16079 7656 16088
rect 7708 16079 7710 16088
rect 7748 16108 7800 16114
rect 7656 16050 7708 16056
rect 7748 16050 7800 16056
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7484 14958 7512 15982
rect 7576 15570 7604 15982
rect 7668 15706 7696 16050
rect 7944 15706 7972 17002
rect 8036 16046 8064 22510
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8128 21486 8156 21966
rect 8220 21894 8248 23122
rect 8312 22778 8340 23684
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8206 21448 8262 21457
rect 8206 21383 8262 21392
rect 8220 21146 8248 21383
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8114 21040 8170 21049
rect 8114 20975 8170 20984
rect 8128 20942 8156 20975
rect 8116 20936 8168 20942
rect 8116 20878 8168 20884
rect 8128 20618 8156 20878
rect 8220 20754 8248 21082
rect 8312 21026 8340 22442
rect 8404 21690 8432 23598
rect 8496 22506 8524 25735
rect 8680 24449 8708 32234
rect 8772 30598 8800 32263
rect 8852 32224 8904 32230
rect 8852 32166 8904 32172
rect 8760 30592 8812 30598
rect 8760 30534 8812 30540
rect 8864 29850 8892 32166
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 9324 30190 9352 30534
rect 9312 30184 9364 30190
rect 9312 30126 9364 30132
rect 8852 29844 8904 29850
rect 8852 29786 8904 29792
rect 8760 29572 8812 29578
rect 8760 29514 8812 29520
rect 8772 28150 8800 29514
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8852 29096 8904 29102
rect 8852 29038 8904 29044
rect 8942 29064 8998 29073
rect 8760 28144 8812 28150
rect 8760 28086 8812 28092
rect 8760 27872 8812 27878
rect 8758 27840 8760 27849
rect 8812 27840 8814 27849
rect 8758 27775 8814 27784
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8666 24440 8722 24449
rect 8666 24375 8722 24384
rect 8668 24064 8720 24070
rect 8668 24006 8720 24012
rect 8680 23730 8708 24006
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 8680 22778 8708 23666
rect 8772 23118 8800 26726
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 8772 22234 8800 23054
rect 8760 22228 8812 22234
rect 8760 22170 8812 22176
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8496 21146 8524 21830
rect 8574 21720 8630 21729
rect 8574 21655 8630 21664
rect 8588 21350 8616 21655
rect 8576 21344 8628 21350
rect 8864 21332 8892 29038
rect 8942 28999 8944 29008
rect 8996 28999 8998 29008
rect 8944 28970 8996 28976
rect 9220 28960 9272 28966
rect 9220 28902 9272 28908
rect 9232 28558 9260 28902
rect 9220 28552 9272 28558
rect 9220 28494 9272 28500
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 9324 28132 9352 30126
rect 9140 28104 9352 28132
rect 9140 27538 9168 28104
rect 9220 27872 9272 27878
rect 9272 27820 9352 27826
rect 9220 27814 9352 27820
rect 9232 27798 9352 27814
rect 9128 27532 9180 27538
rect 9128 27474 9180 27480
rect 9324 27334 9352 27798
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9324 27033 9352 27270
rect 9310 27024 9366 27033
rect 9310 26959 9366 26968
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 9048 24177 9076 24550
rect 9324 24177 9352 24686
rect 9034 24168 9090 24177
rect 9034 24103 9090 24112
rect 9310 24168 9366 24177
rect 9310 24103 9366 24112
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 9232 23361 9260 23666
rect 9218 23352 9274 23361
rect 9218 23287 9274 23296
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 9324 21554 9352 21830
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 8576 21286 8628 21292
rect 8772 21304 8892 21332
rect 9310 21312 9366 21321
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8312 20998 8524 21026
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8220 20726 8340 20754
rect 8128 20590 8248 20618
rect 8312 20602 8340 20726
rect 8220 19718 8248 20590
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8404 20058 8432 20878
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8208 19712 8260 19718
rect 8260 19660 8340 19666
rect 8208 19654 8340 19660
rect 8220 19638 8340 19654
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8220 18358 8248 18702
rect 8208 18352 8260 18358
rect 8208 18294 8260 18300
rect 8312 18222 8340 19638
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8116 18148 8168 18154
rect 8116 18090 8168 18096
rect 8128 17678 8156 18090
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8128 17338 8156 17614
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 8128 16726 8156 17274
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8220 15910 8248 16594
rect 8024 15904 8076 15910
rect 8208 15904 8260 15910
rect 8024 15846 8076 15852
rect 8206 15872 8208 15881
rect 8260 15872 8262 15881
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7484 14618 7512 14894
rect 7576 14890 7604 15506
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7576 14074 7604 14826
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7392 13926 7788 13954
rect 7470 13832 7526 13841
rect 7196 13796 7248 13802
rect 7470 13767 7526 13776
rect 7196 13738 7248 13744
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6736 13252 6788 13258
rect 6840 13246 6960 13274
rect 6736 13194 6788 13200
rect 6748 12782 6776 13194
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6644 12708 6696 12714
rect 6644 12650 6696 12656
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6564 11778 6592 12310
rect 6656 12238 6684 12650
rect 6734 12608 6790 12617
rect 6734 12543 6790 12552
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6748 12170 6776 12543
rect 6840 12306 6868 13126
rect 6932 12374 6960 13246
rect 7116 12986 7144 13330
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6748 11898 6776 12106
rect 6840 11898 6868 12242
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6564 11750 6776 11778
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5814 8392 5870 8401
rect 5814 8327 5870 8336
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5644 5166 5672 5306
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5644 2038 5672 4966
rect 5632 2032 5684 2038
rect 5632 1974 5684 1980
rect 5736 480 5764 6326
rect 5828 5137 5856 8327
rect 5920 7478 5948 8774
rect 6012 8362 6040 8978
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 6104 7954 6132 10406
rect 6196 9178 6224 10542
rect 6656 10470 6684 11086
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6196 8566 6224 9114
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6196 7546 6224 8502
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6656 7546 6684 8502
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 6196 7342 6224 7482
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6748 7206 6776 11750
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6840 11354 6868 11562
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6840 10266 6868 11290
rect 6932 10810 6960 12174
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7024 10674 7052 11222
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7024 10266 7052 10610
rect 7208 10266 7236 13738
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11762 7420 12038
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 6918 9752 6974 9761
rect 7208 9722 7236 10202
rect 7392 9722 7420 10406
rect 6918 9687 6974 9696
rect 7196 9716 7248 9722
rect 6932 9178 6960 9687
rect 7196 9658 7248 9664
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6932 8514 6960 9114
rect 6840 8486 7144 8514
rect 6840 8090 6868 8486
rect 7116 8430 7144 8486
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 5574 5948 6598
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5920 5166 5948 5510
rect 5908 5160 5960 5166
rect 5814 5128 5870 5137
rect 5908 5102 5960 5108
rect 5814 5063 5870 5072
rect 5920 4486 5948 5102
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5828 3534 5856 4082
rect 6104 3618 6132 7142
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6182 6896 6238 6905
rect 6182 6831 6184 6840
rect 6236 6831 6238 6840
rect 6184 6802 6236 6808
rect 6196 6458 6224 6802
rect 6642 6488 6698 6497
rect 6184 6452 6236 6458
rect 6642 6423 6644 6432
rect 6184 6394 6236 6400
rect 6696 6423 6698 6432
rect 6644 6394 6696 6400
rect 6642 6352 6698 6361
rect 6184 6316 6236 6322
rect 6642 6287 6698 6296
rect 6184 6258 6236 6264
rect 6196 4282 6224 6258
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6656 5778 6684 6287
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6656 5370 6684 5714
rect 6920 5704 6972 5710
rect 6734 5672 6790 5681
rect 6734 5607 6790 5616
rect 6840 5652 6920 5658
rect 6840 5646 6972 5652
rect 6840 5630 6960 5646
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6656 5030 6684 5306
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6196 4049 6224 4218
rect 6182 4040 6238 4049
rect 6182 3975 6238 3984
rect 6196 3942 6224 3975
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6656 3738 6684 4694
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6000 3596 6052 3602
rect 6104 3590 6224 3618
rect 6000 3538 6052 3544
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5828 3058 5856 3470
rect 6012 3126 6040 3538
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5828 2650 5856 2994
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5828 2446 5856 2586
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6196 480 6224 3590
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6288 3194 6316 3470
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6748 1306 6776 5607
rect 6840 4826 6868 5630
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6932 4706 6960 5102
rect 6840 4678 6960 4706
rect 6840 4622 6868 4678
rect 6828 4616 6880 4622
rect 6826 4584 6828 4593
rect 6880 4584 6882 4593
rect 6826 4519 6882 4528
rect 6828 4480 6880 4486
rect 7024 4457 7052 6054
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7116 5166 7144 5510
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6828 4422 6880 4428
rect 7010 4448 7066 4457
rect 6840 3670 6868 4422
rect 7010 4383 7066 4392
rect 7010 4176 7066 4185
rect 6920 4140 6972 4146
rect 7010 4111 7066 4120
rect 6920 4082 6972 4088
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6932 3602 6960 4082
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6932 3482 6960 3538
rect 6840 3454 6960 3482
rect 6840 3369 6868 3454
rect 6920 3392 6972 3398
rect 6826 3360 6882 3369
rect 6920 3334 6972 3340
rect 6826 3295 6882 3304
rect 6840 3194 6868 3295
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6932 3097 6960 3334
rect 6918 3088 6974 3097
rect 6918 3023 6974 3032
rect 6564 1278 6776 1306
rect 6564 480 6592 1278
rect 7024 1034 7052 4111
rect 7116 2650 7144 4966
rect 7208 4214 7236 9658
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7208 3777 7236 4150
rect 7300 4146 7328 9522
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7392 8430 7420 8910
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7484 7274 7512 13767
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7576 12102 7604 12922
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7576 11762 7604 12038
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 11014 7604 11698
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10674 7604 10950
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10198 7604 10610
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7576 9178 7604 9998
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7562 8664 7618 8673
rect 7562 8599 7618 8608
rect 7576 8294 7604 8599
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7576 8022 7604 8230
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7484 6934 7512 7210
rect 7472 6928 7524 6934
rect 7524 6876 7604 6882
rect 7472 6870 7604 6876
rect 7484 6854 7604 6870
rect 7470 5808 7526 5817
rect 7470 5743 7526 5752
rect 7484 5642 7512 5743
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7470 4720 7526 4729
rect 7392 4214 7420 4694
rect 7470 4655 7526 4664
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7484 4026 7512 4655
rect 7392 3998 7512 4026
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7194 3768 7250 3777
rect 7194 3703 7250 3712
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7208 2854 7236 3334
rect 7300 2922 7328 3878
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1465 7144 2246
rect 7102 1456 7158 1465
rect 7102 1391 7158 1400
rect 6932 1006 7052 1034
rect 6932 480 6960 1006
rect 7392 480 7420 3998
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7484 2854 7512 2926
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7484 2553 7512 2790
rect 7470 2544 7526 2553
rect 7576 2514 7604 6854
rect 7760 5930 7788 13926
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7852 11354 7880 12650
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7852 7546 7880 7822
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7852 7002 7880 7482
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7944 6905 7972 15438
rect 8036 12889 8064 15846
rect 8206 15807 8262 15816
rect 8312 15722 8340 17070
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8220 15706 8340 15722
rect 8404 15706 8432 16526
rect 8496 16522 8524 20998
rect 8588 18306 8616 21286
rect 8772 19174 8800 21304
rect 9310 21247 9366 21256
rect 8944 21140 8996 21146
rect 8864 21100 8944 21128
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8588 18278 8708 18306
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8588 17542 8616 18158
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8208 15700 8340 15706
rect 8260 15694 8340 15700
rect 8208 15642 8260 15648
rect 8206 15600 8262 15609
rect 8206 15535 8208 15544
rect 8260 15535 8262 15544
rect 8208 15506 8260 15512
rect 8220 15094 8248 15506
rect 8312 15162 8340 15694
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8208 15088 8260 15094
rect 8404 15042 8432 15506
rect 8496 15502 8524 16050
rect 8588 15570 8616 17478
rect 8680 16794 8708 18278
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8208 15030 8260 15036
rect 8312 15014 8432 15042
rect 8114 13696 8170 13705
rect 8114 13631 8170 13640
rect 8022 12880 8078 12889
rect 8022 12815 8078 12824
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11801 8064 12038
rect 8022 11792 8078 11801
rect 8022 11727 8078 11736
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8036 11354 8064 11630
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 8128 10266 8156 13631
rect 8312 13462 8340 15014
rect 8496 14482 8524 15438
rect 8680 15162 8708 16594
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8772 15042 8800 19110
rect 8864 17678 8892 21100
rect 8944 21082 8996 21088
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9324 18329 9352 21247
rect 9310 18320 9366 18329
rect 9310 18255 9366 18264
rect 8944 18080 8996 18086
rect 9312 18080 9364 18086
rect 8944 18022 8996 18028
rect 9310 18048 9312 18057
rect 9364 18048 9366 18057
rect 8956 17746 8984 18022
rect 9310 17983 9366 17992
rect 9310 17912 9366 17921
rect 9310 17847 9366 17856
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8956 17524 8984 17682
rect 8864 17496 8984 17524
rect 8864 17338 8892 17496
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 8864 15978 8892 16730
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 9324 16114 9352 17847
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8588 15014 8800 15042
rect 8864 15026 8892 15574
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 9324 15026 9352 16050
rect 8852 15020 8904 15026
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8220 12986 8248 13330
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 11898 8248 12242
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8220 11121 8248 11834
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 8206 11112 8262 11121
rect 8206 11047 8262 11056
rect 8312 10810 8340 11766
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8128 9586 8156 10202
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8128 9081 8156 9318
rect 8114 9072 8170 9081
rect 8114 9007 8170 9016
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8220 8294 8248 8978
rect 8208 8288 8260 8294
rect 8206 8256 8208 8265
rect 8260 8256 8262 8265
rect 8206 8191 8262 8200
rect 8220 8090 8248 8191
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8312 7970 8340 10134
rect 8404 7993 8432 13806
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 12986 8524 13670
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8496 12442 8524 12922
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8482 11656 8538 11665
rect 8482 11591 8538 11600
rect 8496 11354 8524 11591
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8496 10742 8524 11290
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8496 10305 8524 10678
rect 8482 10296 8538 10305
rect 8482 10231 8538 10240
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8036 7942 8340 7970
rect 8390 7984 8446 7993
rect 7930 6896 7986 6905
rect 7930 6831 7986 6840
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7944 6390 7972 6734
rect 8036 6458 8064 7942
rect 8390 7919 8446 7928
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8116 7200 8168 7206
rect 8114 7168 8116 7177
rect 8168 7168 8170 7177
rect 8114 7103 8170 7112
rect 8220 6497 8248 7686
rect 8404 7018 8432 7919
rect 8312 6990 8432 7018
rect 8312 6730 8340 6990
rect 8496 6866 8524 10066
rect 8588 8673 8616 15014
rect 8852 14962 8904 14968
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9416 14958 9444 33079
rect 9496 33050 9548 33056
rect 9508 32026 9536 33050
rect 9496 32020 9548 32026
rect 9496 31962 9548 31968
rect 9600 31958 9628 33782
rect 9692 32978 9720 34002
rect 9784 33538 9812 39520
rect 10152 39494 10272 39520
rect 10048 34944 10100 34950
rect 10048 34886 10100 34892
rect 10060 34649 10088 34886
rect 10046 34640 10102 34649
rect 10046 34575 10102 34584
rect 10060 34542 10088 34575
rect 10048 34536 10100 34542
rect 10048 34478 10100 34484
rect 10060 34202 10088 34478
rect 10048 34196 10100 34202
rect 10048 34138 10100 34144
rect 10048 34060 10100 34066
rect 10048 34002 10100 34008
rect 9784 33510 9904 33538
rect 10060 33522 10088 34002
rect 9680 32972 9732 32978
rect 9680 32914 9732 32920
rect 9588 31952 9640 31958
rect 9588 31894 9640 31900
rect 9600 29578 9628 31894
rect 9692 30802 9720 32914
rect 9680 30796 9732 30802
rect 9680 30738 9732 30744
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 9496 29504 9548 29510
rect 9496 29446 9548 29452
rect 9508 29170 9536 29446
rect 9588 29232 9640 29238
rect 9588 29174 9640 29180
rect 9496 29164 9548 29170
rect 9496 29106 9548 29112
rect 9508 27946 9536 29106
rect 9496 27940 9548 27946
rect 9496 27882 9548 27888
rect 9508 27674 9536 27882
rect 9496 27668 9548 27674
rect 9496 27610 9548 27616
rect 9600 26602 9628 29174
rect 9680 29028 9732 29034
rect 9680 28970 9732 28976
rect 9692 28558 9720 28970
rect 9876 28948 9904 33510
rect 10048 33516 10100 33522
rect 10048 33458 10100 33464
rect 10048 32972 10100 32978
rect 10048 32914 10100 32920
rect 10060 32570 10088 32914
rect 10048 32564 10100 32570
rect 10048 32506 10100 32512
rect 10060 32473 10088 32506
rect 10046 32464 10102 32473
rect 10046 32399 10102 32408
rect 9956 31816 10008 31822
rect 9956 31758 10008 31764
rect 9968 30326 9996 31758
rect 10138 31240 10194 31249
rect 10138 31175 10194 31184
rect 10152 31142 10180 31175
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 10244 30920 10272 39494
rect 10414 33416 10470 33425
rect 10414 33351 10470 33360
rect 10322 33144 10378 33153
rect 10322 33079 10378 33088
rect 10336 32570 10364 33079
rect 10324 32564 10376 32570
rect 10324 32506 10376 32512
rect 10336 32366 10364 32506
rect 10324 32360 10376 32366
rect 10324 32302 10376 32308
rect 10244 30892 10364 30920
rect 10232 30796 10284 30802
rect 10232 30738 10284 30744
rect 9956 30320 10008 30326
rect 9956 30262 10008 30268
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 10048 29028 10100 29034
rect 10048 28970 10100 28976
rect 9784 28920 9904 28948
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 9784 27690 9812 28920
rect 9692 27662 9812 27690
rect 9692 26761 9720 27662
rect 9772 27532 9824 27538
rect 9772 27474 9824 27480
rect 9784 26790 9812 27474
rect 10060 27033 10088 28970
rect 10046 27024 10102 27033
rect 10046 26959 10102 26968
rect 9772 26784 9824 26790
rect 9678 26752 9734 26761
rect 9772 26726 9824 26732
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 9678 26687 9734 26696
rect 9600 26586 9720 26602
rect 9600 26580 9732 26586
rect 9600 26574 9680 26580
rect 9496 26376 9548 26382
rect 9496 26318 9548 26324
rect 9508 25974 9536 26318
rect 9496 25968 9548 25974
rect 9496 25910 9548 25916
rect 9600 25498 9628 26574
rect 9680 26522 9732 26528
rect 9678 26480 9734 26489
rect 9678 26415 9734 26424
rect 9692 26314 9720 26415
rect 9680 26308 9732 26314
rect 9680 26250 9732 26256
rect 9680 25968 9732 25974
rect 9680 25910 9732 25916
rect 9692 25702 9720 25910
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9496 25220 9548 25226
rect 9496 25162 9548 25168
rect 9508 24818 9536 25162
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9508 24410 9536 24754
rect 9600 24614 9628 25094
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9600 23633 9628 24550
rect 9692 24313 9720 25638
rect 9678 24304 9734 24313
rect 9678 24239 9734 24248
rect 9692 23769 9720 24239
rect 9678 23760 9734 23769
rect 9678 23695 9734 23704
rect 9586 23624 9642 23633
rect 9586 23559 9642 23568
rect 9680 23588 9732 23594
rect 9680 23530 9732 23536
rect 9692 23118 9720 23530
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9680 22976 9732 22982
rect 9680 22918 9732 22924
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9508 21078 9536 21490
rect 9496 21072 9548 21078
rect 9496 21014 9548 21020
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 8680 11762 8708 14894
rect 8852 14816 8904 14822
rect 9508 14770 9536 20538
rect 9586 19408 9642 19417
rect 9586 19343 9642 19352
rect 9600 18873 9628 19343
rect 9586 18864 9642 18873
rect 9586 18799 9642 18808
rect 9692 18766 9720 22918
rect 9784 21185 9812 26726
rect 10060 26450 10088 26726
rect 10048 26444 10100 26450
rect 10048 26386 10100 26392
rect 10060 25974 10088 26386
rect 10048 25968 10100 25974
rect 10048 25910 10100 25916
rect 10152 25786 10180 29990
rect 10244 29850 10272 30738
rect 10232 29844 10284 29850
rect 10232 29786 10284 29792
rect 10244 28762 10272 29786
rect 10336 29034 10364 30892
rect 10324 29028 10376 29034
rect 10324 28970 10376 28976
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 10244 28014 10272 28698
rect 10324 28416 10376 28422
rect 10324 28358 10376 28364
rect 10232 28008 10284 28014
rect 10232 27950 10284 27956
rect 10336 27674 10364 28358
rect 10324 27668 10376 27674
rect 10324 27610 10376 27616
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10244 26790 10272 27406
rect 10428 26874 10456 33351
rect 10508 31680 10560 31686
rect 10508 31622 10560 31628
rect 10520 31278 10548 31622
rect 10508 31272 10560 31278
rect 10508 31214 10560 31220
rect 10612 30977 10640 39520
rect 10980 35714 11008 39520
rect 11348 37874 11376 39520
rect 11336 37868 11388 37874
rect 11336 37810 11388 37816
rect 11808 37754 11836 39520
rect 10704 35686 11008 35714
rect 11348 37726 11836 37754
rect 10598 30968 10654 30977
rect 10598 30903 10654 30912
rect 10704 30841 10732 35686
rect 11152 35148 11204 35154
rect 11152 35090 11204 35096
rect 11060 34672 11112 34678
rect 11060 34614 11112 34620
rect 10784 33924 10836 33930
rect 10784 33866 10836 33872
rect 10796 31278 10824 33866
rect 11072 33674 11100 34614
rect 11164 34202 11192 35090
rect 11152 34196 11204 34202
rect 11152 34138 11204 34144
rect 11244 34196 11296 34202
rect 11244 34138 11296 34144
rect 11152 34060 11204 34066
rect 11152 34002 11204 34008
rect 10980 33658 11100 33674
rect 10968 33652 11100 33658
rect 11020 33646 11100 33652
rect 10968 33594 11020 33600
rect 10874 33552 10930 33561
rect 11164 33538 11192 34002
rect 11256 33658 11284 34138
rect 11244 33652 11296 33658
rect 11244 33594 11296 33600
rect 10874 33487 10930 33496
rect 10980 33510 11192 33538
rect 10888 33114 10916 33487
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 10784 31272 10836 31278
rect 10784 31214 10836 31220
rect 10796 30938 10824 31214
rect 10784 30932 10836 30938
rect 10784 30874 10836 30880
rect 10690 30832 10746 30841
rect 10690 30767 10746 30776
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10508 30048 10560 30054
rect 10508 29990 10560 29996
rect 10520 29782 10548 29990
rect 10508 29776 10560 29782
rect 10508 29718 10560 29724
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10520 29034 10548 29582
rect 10508 29028 10560 29034
rect 10508 28970 10560 28976
rect 10520 27849 10548 28970
rect 10612 28218 10640 30194
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 10796 28218 10824 28494
rect 10600 28212 10652 28218
rect 10600 28154 10652 28160
rect 10784 28212 10836 28218
rect 10784 28154 10836 28160
rect 10506 27840 10562 27849
rect 10506 27775 10562 27784
rect 10336 26846 10456 26874
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 10230 26616 10286 26625
rect 10230 26551 10286 26560
rect 10244 26042 10272 26551
rect 10232 26036 10284 26042
rect 10232 25978 10284 25984
rect 10152 25758 10272 25786
rect 9864 25696 9916 25702
rect 9862 25664 9864 25673
rect 10140 25696 10192 25702
rect 9916 25664 9918 25673
rect 10140 25638 10192 25644
rect 9862 25599 9918 25608
rect 10048 25424 10100 25430
rect 10046 25392 10048 25401
rect 10100 25392 10102 25401
rect 10046 25327 10102 25336
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9876 23866 9904 24550
rect 10060 24410 10088 25230
rect 10152 24818 10180 25638
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 10152 24410 10180 24754
rect 10244 24750 10272 25758
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9862 23760 9918 23769
rect 9862 23695 9918 23704
rect 9876 22982 9904 23695
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 10244 22642 10272 23122
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10046 22128 10102 22137
rect 10046 22063 10048 22072
rect 10100 22063 10102 22072
rect 10048 22034 10100 22040
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9876 21350 9904 21966
rect 10060 21690 10088 22034
rect 10244 22030 10272 22578
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9770 21176 9826 21185
rect 9770 21111 9826 21120
rect 9876 20913 9904 21286
rect 10244 21146 10272 21966
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 10140 20936 10192 20942
rect 9862 20904 9918 20913
rect 10140 20878 10192 20884
rect 9862 20839 9918 20848
rect 10048 20800 10100 20806
rect 9770 20768 9826 20777
rect 10048 20742 10100 20748
rect 9770 20703 9826 20712
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9600 18290 9628 18634
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9600 17921 9628 18226
rect 9586 17912 9642 17921
rect 9586 17847 9642 17856
rect 9692 16810 9720 18566
rect 9784 17898 9812 20703
rect 10060 20398 10088 20742
rect 10152 20602 10180 20878
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9954 19952 10010 19961
rect 9954 19887 9956 19896
rect 10008 19887 10010 19896
rect 9956 19858 10008 19864
rect 9968 19310 9996 19858
rect 10060 19514 10088 20334
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 10048 19168 10100 19174
rect 10336 19122 10364 26846
rect 10416 26784 10468 26790
rect 10416 26726 10468 26732
rect 10428 25294 10456 26726
rect 10520 25838 10548 27775
rect 10612 26382 10640 28154
rect 10784 27668 10836 27674
rect 10784 27610 10836 27616
rect 10692 27328 10744 27334
rect 10692 27270 10744 27276
rect 10704 26858 10732 27270
rect 10796 26994 10824 27610
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10692 26852 10744 26858
rect 10692 26794 10744 26800
rect 10704 26586 10732 26794
rect 10692 26580 10744 26586
rect 10692 26522 10744 26528
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 10690 25664 10746 25673
rect 10612 25498 10640 25638
rect 10690 25599 10746 25608
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 10416 25288 10468 25294
rect 10416 25230 10468 25236
rect 10612 24954 10640 25298
rect 10600 24948 10652 24954
rect 10600 24890 10652 24896
rect 10416 24744 10468 24750
rect 10416 24686 10468 24692
rect 10048 19110 10100 19116
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9876 18086 9904 18702
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9784 17870 9904 17898
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9784 17270 9812 17682
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9600 16794 9720 16810
rect 9588 16788 9720 16794
rect 9640 16782 9720 16788
rect 9588 16730 9640 16736
rect 9600 16046 9628 16730
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9692 14793 9720 15098
rect 8852 14758 8904 14764
rect 8864 14618 8892 14758
rect 9324 14742 9536 14770
rect 9678 14784 9734 14793
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8772 13870 8800 14554
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8864 13530 8892 14554
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8956 13870 8984 13942
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8772 11642 8800 13398
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8864 12646 8892 13126
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8852 12640 8904 12646
rect 8850 12608 8852 12617
rect 8904 12608 8906 12617
rect 8850 12543 8906 12552
rect 8850 12336 8906 12345
rect 8850 12271 8906 12280
rect 8864 12238 8892 12271
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8864 11762 8892 12174
rect 9048 12170 9076 12718
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8680 11614 8800 11642
rect 8574 8664 8630 8673
rect 8574 8599 8630 8608
rect 8680 7970 8708 11614
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8772 8786 8800 11494
rect 8864 11354 8892 11698
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8864 10674 8892 10950
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8864 10266 8892 10610
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8864 10062 8892 10202
rect 8956 10169 8984 10406
rect 9048 10198 9076 10542
rect 9036 10192 9088 10198
rect 8942 10160 8998 10169
rect 9036 10134 9088 10140
rect 9324 10130 9352 14742
rect 9678 14719 9734 14728
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 13938 9536 14214
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9494 13832 9550 13841
rect 9494 13767 9550 13776
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 11558 9444 13126
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9402 10840 9458 10849
rect 9402 10775 9458 10784
rect 9416 10606 9444 10775
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9402 10296 9458 10305
rect 9402 10231 9458 10240
rect 8942 10095 8998 10104
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8864 9654 8892 9998
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 9324 9722 9352 9862
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 9310 9616 9366 9625
rect 8864 8906 8892 9590
rect 9310 9551 9366 9560
rect 9126 9480 9182 9489
rect 9126 9415 9128 9424
rect 9180 9415 9182 9424
rect 9128 9386 9180 9392
rect 9324 9382 9352 9551
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9416 9092 9444 10231
rect 9407 9064 9444 9092
rect 9312 8968 9364 8974
rect 9407 8956 9435 9064
rect 9508 8974 9536 13767
rect 9600 13530 9628 14486
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 14074 9720 14350
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9692 13462 9720 13806
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9600 12782 9628 13262
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9692 12646 9720 13398
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9496 8968 9548 8974
rect 9407 8928 9444 8956
rect 9312 8910 9364 8916
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8772 8758 8892 8786
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8588 7942 8708 7970
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8206 6488 8262 6497
rect 8024 6452 8076 6458
rect 8404 6458 8432 6802
rect 8484 6656 8536 6662
rect 8588 6633 8616 7942
rect 8772 7750 8800 8230
rect 8864 7954 8892 8758
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8680 7342 8708 7686
rect 8864 7426 8892 7890
rect 8956 7886 8984 8230
rect 9232 8022 9260 8366
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8944 7472 8996 7478
rect 8942 7440 8944 7449
rect 8996 7440 8998 7449
rect 8864 7398 8942 7426
rect 8942 7375 8998 7384
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 6798 8708 7278
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8484 6598 8536 6604
rect 8574 6624 8630 6633
rect 8206 6423 8262 6432
rect 8392 6452 8444 6458
rect 8024 6394 8076 6400
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 8036 6225 8064 6394
rect 8220 6338 8248 6423
rect 8392 6394 8444 6400
rect 8220 6310 8340 6338
rect 8312 6254 8340 6310
rect 8300 6248 8352 6254
rect 8022 6216 8078 6225
rect 8300 6190 8352 6196
rect 8022 6151 8078 6160
rect 8496 6118 8524 6598
rect 8574 6559 8630 6568
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 7760 5902 7880 5930
rect 7746 5808 7802 5817
rect 7746 5743 7802 5752
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7668 3738 7696 4082
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7668 2990 7696 3674
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7470 2479 7526 2488
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7668 2446 7696 2926
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7760 480 7788 5743
rect 7852 3641 7880 5902
rect 7944 5710 7972 6054
rect 8496 5846 8524 6054
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5574 8156 5646
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8128 5370 8156 5510
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8220 4758 8248 4966
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8312 4434 8340 4490
rect 8220 4406 8340 4434
rect 8022 3904 8078 3913
rect 8022 3839 8078 3848
rect 8036 3738 8064 3839
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7838 3632 7894 3641
rect 7838 3567 7894 3576
rect 7852 3194 7880 3567
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 8128 2922 8156 3470
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 8128 2530 8156 2858
rect 8220 2650 8248 4406
rect 8404 4282 8432 5578
rect 8588 4826 8616 6190
rect 8680 5574 8708 6258
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8482 4584 8538 4593
rect 8482 4519 8538 4528
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8390 4040 8446 4049
rect 8390 3975 8446 3984
rect 8404 3942 8432 3975
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8404 3738 8432 3878
rect 8496 3738 8524 4519
rect 8588 4146 8616 4762
rect 8772 4162 8800 6802
rect 8864 5846 8892 6938
rect 9232 6905 9260 7142
rect 9218 6896 9274 6905
rect 9218 6831 9274 6840
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8864 5030 8892 5510
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9324 5137 9352 8910
rect 9416 7290 9444 8928
rect 9496 8910 9548 8916
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9508 8022 9536 8774
rect 9600 8242 9628 11494
rect 9692 11286 9720 12174
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9692 10810 9720 11222
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9784 9081 9812 17070
rect 9876 16017 9904 17870
rect 9968 17814 9996 18634
rect 10060 18193 10088 19110
rect 10244 19094 10364 19122
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 10152 18426 10180 18838
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10244 18306 10272 19094
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10152 18278 10272 18306
rect 10336 18290 10364 18906
rect 10324 18284 10376 18290
rect 10046 18184 10102 18193
rect 10046 18119 10102 18128
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9956 17808 10008 17814
rect 9956 17750 10008 17756
rect 9968 17338 9996 17750
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9968 16153 9996 17274
rect 9954 16144 10010 16153
rect 9954 16079 10010 16088
rect 9862 16008 9918 16017
rect 9862 15943 9918 15952
rect 9862 15056 9918 15065
rect 9862 14991 9918 15000
rect 9876 14618 9904 14991
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9876 14226 9904 14554
rect 9968 14550 9996 16079
rect 10060 15502 10088 18022
rect 10152 15609 10180 18278
rect 10324 18226 10376 18232
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10244 16794 10272 18090
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10336 16998 10364 17138
rect 10428 17134 10456 24686
rect 10704 24274 10732 25599
rect 10784 25220 10836 25226
rect 10784 25162 10836 25168
rect 10796 24682 10824 25162
rect 10784 24676 10836 24682
rect 10784 24618 10836 24624
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10704 23594 10732 24210
rect 10692 23588 10744 23594
rect 10692 23530 10744 23536
rect 10704 23254 10732 23530
rect 10692 23248 10744 23254
rect 10692 23190 10744 23196
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10520 20058 10548 20946
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10520 19802 10548 19994
rect 10520 19774 10640 19802
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10520 19378 10548 19654
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10520 18426 10548 19314
rect 10612 18970 10640 19774
rect 10888 19360 10916 33050
rect 10980 32570 11008 33510
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 10968 32564 11020 32570
rect 10968 32506 11020 32512
rect 11072 32434 11100 32846
rect 11256 32842 11284 33594
rect 11244 32836 11296 32842
rect 11244 32778 11296 32784
rect 11060 32428 11112 32434
rect 11060 32370 11112 32376
rect 10968 32224 11020 32230
rect 10968 32166 11020 32172
rect 10980 31958 11008 32166
rect 11072 32026 11100 32370
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 10968 31952 11020 31958
rect 10968 31894 11020 31900
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 11256 30870 11284 31078
rect 11244 30864 11296 30870
rect 11244 30806 11296 30812
rect 11256 30394 11284 30806
rect 11244 30388 11296 30394
rect 11244 30330 11296 30336
rect 11150 30288 11206 30297
rect 11150 30223 11206 30232
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10980 29866 11008 29990
rect 11164 29866 11192 30223
rect 10980 29838 11192 29866
rect 10968 29776 11020 29782
rect 10968 29718 11020 29724
rect 10980 29306 11008 29718
rect 10968 29300 11020 29306
rect 10968 29242 11020 29248
rect 11060 28620 11112 28626
rect 11060 28562 11112 28568
rect 11072 28218 11100 28562
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10980 26518 11008 26930
rect 10968 26512 11020 26518
rect 10968 26454 11020 26460
rect 10980 24750 11008 26454
rect 10968 24744 11020 24750
rect 10968 24686 11020 24692
rect 10980 24410 11008 24686
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 11058 23352 11114 23361
rect 11058 23287 11060 23296
rect 11112 23287 11114 23296
rect 11060 23258 11112 23264
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 10980 20602 11008 22714
rect 11164 22234 11192 29838
rect 11244 29844 11296 29850
rect 11244 29786 11296 29792
rect 11256 29306 11284 29786
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11348 22658 11376 37726
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 12176 34490 12204 39520
rect 12256 37868 12308 37874
rect 12256 37810 12308 37816
rect 11992 34462 12204 34490
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11428 33312 11480 33318
rect 11428 33254 11480 33260
rect 11440 31754 11468 33254
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11612 33040 11664 33046
rect 11992 32994 12020 34462
rect 12072 34400 12124 34406
rect 12072 34342 12124 34348
rect 12084 34134 12112 34342
rect 12072 34128 12124 34134
rect 12072 34070 12124 34076
rect 12084 33522 12112 34070
rect 12072 33516 12124 33522
rect 12072 33458 12124 33464
rect 12084 33318 12112 33458
rect 12162 33416 12218 33425
rect 12162 33351 12164 33360
rect 12216 33351 12218 33360
rect 12164 33322 12216 33328
rect 12072 33312 12124 33318
rect 12072 33254 12124 33260
rect 11612 32982 11664 32988
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 11532 32026 11560 32710
rect 11624 32570 11652 32982
rect 11900 32966 12020 32994
rect 11612 32564 11664 32570
rect 11612 32506 11664 32512
rect 11900 32337 11928 32966
rect 12084 32910 12112 33254
rect 11980 32904 12032 32910
rect 11980 32846 12032 32852
rect 12072 32904 12124 32910
rect 12072 32846 12124 32852
rect 11992 32570 12020 32846
rect 11980 32564 12032 32570
rect 11980 32506 12032 32512
rect 11886 32328 11942 32337
rect 11886 32263 11942 32272
rect 11992 32230 12020 32506
rect 12070 32328 12126 32337
rect 12070 32263 12126 32272
rect 11980 32224 12032 32230
rect 11980 32166 12032 32172
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 11428 31748 11480 31754
rect 11428 31690 11480 31696
rect 11440 31142 11468 31690
rect 11532 31482 11560 31962
rect 11520 31476 11572 31482
rect 11520 31418 11572 31424
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 11428 31136 11480 31142
rect 11428 31078 11480 31084
rect 11532 30938 11560 31282
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11520 30932 11572 30938
rect 11520 30874 11572 30880
rect 11532 29782 11560 30874
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11520 29776 11572 29782
rect 11520 29718 11572 29724
rect 11520 29504 11572 29510
rect 11520 29446 11572 29452
rect 11532 28558 11560 29446
rect 12084 29034 12112 32263
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 12072 29028 12124 29034
rect 12072 28970 12124 28976
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11532 28218 11560 28494
rect 11520 28212 11572 28218
rect 11520 28154 11572 28160
rect 11532 27606 11560 28154
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11520 27600 11572 27606
rect 11520 27542 11572 27548
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 11440 26790 11468 27406
rect 11532 27130 11560 27542
rect 11520 27124 11572 27130
rect 11520 27066 11572 27072
rect 11428 26784 11480 26790
rect 11428 26726 11480 26732
rect 11440 25673 11468 26726
rect 11532 26042 11560 27066
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 11426 25664 11482 25673
rect 11426 25599 11482 25608
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11992 24614 12020 28970
rect 12268 28914 12296 37810
rect 12544 35034 12572 39520
rect 12544 35006 12664 35034
rect 12532 34944 12584 34950
rect 12532 34886 12584 34892
rect 12544 33998 12572 34886
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12544 33674 12572 33934
rect 12360 33646 12572 33674
rect 12360 33454 12388 33646
rect 12348 33448 12400 33454
rect 12348 33390 12400 33396
rect 12440 33312 12492 33318
rect 12440 33254 12492 33260
rect 12348 31884 12400 31890
rect 12348 31826 12400 31832
rect 12360 31770 12388 31826
rect 12452 31770 12480 33254
rect 12636 32230 12664 35006
rect 12898 33552 12954 33561
rect 12898 33487 12954 33496
rect 12912 33386 12940 33487
rect 12900 33380 12952 33386
rect 12900 33322 12952 33328
rect 12808 33312 12860 33318
rect 12808 33254 12860 33260
rect 12820 33114 12848 33254
rect 12808 33108 12860 33114
rect 12808 33050 12860 33056
rect 12820 32434 12848 33050
rect 12808 32428 12860 32434
rect 12808 32370 12860 32376
rect 12624 32224 12676 32230
rect 12624 32166 12676 32172
rect 12360 31742 12480 31770
rect 12360 31482 12388 31742
rect 12348 31476 12400 31482
rect 12348 31418 12400 31424
rect 12438 30152 12494 30161
rect 12438 30087 12494 30096
rect 12452 29889 12480 30087
rect 12438 29880 12494 29889
rect 12438 29815 12494 29824
rect 12084 28886 12296 28914
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11518 24168 11574 24177
rect 11518 24103 11574 24112
rect 11532 23866 11560 24103
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11440 22778 11468 23190
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11348 22630 11468 22658
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11152 22092 11204 22098
rect 11440 22080 11468 22630
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11440 22052 11560 22080
rect 11152 22034 11204 22040
rect 11164 21944 11192 22034
rect 11164 21916 11376 21944
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11164 20398 11192 20538
rect 11152 20392 11204 20398
rect 11152 20334 11204 20340
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10796 19332 10916 19360
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10612 18306 10640 18770
rect 10520 18278 10640 18306
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10520 18086 10548 18278
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10336 16590 10364 16934
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10414 16552 10470 16561
rect 10336 15638 10364 16526
rect 10414 16487 10470 16496
rect 10428 15910 10456 16487
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10324 15632 10376 15638
rect 10138 15600 10194 15609
rect 10324 15574 10376 15580
rect 10414 15600 10470 15609
rect 10138 15535 10194 15544
rect 10414 15535 10470 15544
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10060 15162 10088 15438
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10324 14952 10376 14958
rect 10046 14920 10102 14929
rect 10324 14894 10376 14900
rect 10428 14906 10456 15535
rect 10520 15042 10548 18022
rect 10598 17640 10654 17649
rect 10598 17575 10654 17584
rect 10612 17338 10640 17575
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10612 17134 10640 17274
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10704 16810 10732 18294
rect 10796 18057 10824 19332
rect 10874 19136 10930 19145
rect 10874 19071 10930 19080
rect 10782 18048 10838 18057
rect 10782 17983 10838 17992
rect 10796 17066 10824 17983
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10704 16782 10824 16810
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10612 15706 10640 16594
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10704 15162 10732 16594
rect 10796 15201 10824 16782
rect 10782 15192 10838 15201
rect 10692 15156 10744 15162
rect 10782 15127 10838 15136
rect 10692 15098 10744 15104
rect 10520 15014 10732 15042
rect 10046 14855 10102 14864
rect 9956 14544 10008 14550
rect 9956 14486 10008 14492
rect 9876 14198 9996 14226
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 12306 9904 14010
rect 9968 13190 9996 14198
rect 10060 14074 10088 14855
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10138 14376 10194 14385
rect 10138 14311 10194 14320
rect 10152 14278 10180 14311
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 10060 12986 10088 13874
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10152 12866 10180 14214
rect 10244 13977 10272 14758
rect 10230 13968 10286 13977
rect 10230 13903 10286 13912
rect 9968 12838 10180 12866
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9770 9072 9826 9081
rect 9770 9007 9826 9016
rect 9600 8214 9720 8242
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9416 7262 9536 7290
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9416 7002 9444 7142
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9402 6896 9458 6905
rect 9508 6866 9536 7262
rect 9402 6831 9458 6840
rect 9496 6860 9548 6866
rect 9310 5128 9366 5137
rect 9310 5063 9366 5072
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8864 4486 8892 4966
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8680 4134 8800 4162
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8404 2990 8432 3674
rect 8680 3618 8708 4134
rect 8758 4040 8814 4049
rect 8758 3975 8760 3984
rect 8812 3975 8814 3984
rect 8760 3946 8812 3952
rect 8758 3768 8814 3777
rect 8758 3703 8814 3712
rect 8496 3590 8708 3618
rect 8496 3097 8524 3590
rect 8576 3120 8628 3126
rect 8482 3088 8538 3097
rect 8576 3062 8628 3068
rect 8482 3023 8538 3032
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8496 2650 8524 3023
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8128 2502 8248 2530
rect 8220 480 8248 2502
rect 8588 480 8616 3062
rect 8772 1306 8800 3703
rect 8864 3194 8892 4422
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 9324 4078 9352 5063
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3466 9352 3878
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 9324 2922 9352 3402
rect 9416 3126 9444 6831
rect 9496 6802 9548 6808
rect 9508 6390 9536 6802
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9496 6112 9548 6118
rect 9494 6080 9496 6089
rect 9548 6080 9550 6089
rect 9494 6015 9550 6024
rect 9600 5930 9628 7686
rect 9692 7313 9720 8214
rect 9784 7342 9812 9007
rect 9772 7336 9824 7342
rect 9678 7304 9734 7313
rect 9772 7278 9824 7284
rect 9678 7239 9734 7248
rect 9692 6254 9720 7239
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6934 9812 7142
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9876 6746 9904 12242
rect 9968 9178 9996 12838
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10060 11898 10088 12718
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10152 12442 10180 12582
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10046 11792 10102 11801
rect 10046 11727 10102 11736
rect 10060 11558 10088 11727
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11354 10088 11494
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10244 9178 10272 13903
rect 10336 13705 10364 14894
rect 10428 14878 10640 14906
rect 10416 13728 10468 13734
rect 10322 13696 10378 13705
rect 10416 13670 10468 13676
rect 10322 13631 10378 13640
rect 10322 13424 10378 13433
rect 10322 13359 10378 13368
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 9968 8430 9996 9114
rect 10244 9058 10272 9114
rect 10152 9030 10272 9058
rect 9956 8424 10008 8430
rect 10008 8384 10088 8412
rect 9956 8366 10008 8372
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9784 6718 9904 6746
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9784 6118 9812 6718
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9600 5914 9812 5930
rect 9600 5908 9824 5914
rect 9600 5902 9772 5908
rect 9600 5794 9628 5902
rect 9772 5850 9824 5856
rect 9508 5766 9628 5794
rect 9680 5772 9732 5778
rect 9508 5098 9536 5766
rect 9680 5714 9732 5720
rect 9692 5658 9720 5714
rect 9600 5630 9720 5658
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9508 3398 9536 5034
rect 9600 4554 9628 5630
rect 9770 5264 9826 5273
rect 9770 5199 9826 5208
rect 9784 4826 9812 5199
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9876 4729 9904 6598
rect 9862 4720 9918 4729
rect 9862 4655 9918 4664
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9678 3768 9734 3777
rect 9678 3703 9734 3712
rect 9692 3670 9720 3703
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9508 2990 9536 3334
rect 9692 3194 9720 3606
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9494 2816 9550 2825
rect 9494 2751 9550 2760
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8772 1278 8984 1306
rect 8956 480 8984 1278
rect 9508 610 9536 2751
rect 9600 2650 9628 2858
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9404 604 9456 610
rect 9404 546 9456 552
rect 9496 604 9548 610
rect 9496 546 9548 552
rect 9416 480 9444 546
rect 9784 480 9812 4082
rect 9968 3602 9996 7958
rect 10060 4078 10088 8384
rect 10152 8022 10180 9030
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8265 10272 8910
rect 10230 8256 10286 8265
rect 10230 8191 10286 8200
rect 10244 8090 10272 8191
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 10244 7410 10272 7754
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10138 7168 10194 7177
rect 10138 7103 10194 7112
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 10152 480 10180 7103
rect 10244 7002 10272 7346
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10244 6322 10272 6938
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10244 3942 10272 4762
rect 10336 4146 10364 13359
rect 10428 12986 10456 13670
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10428 11354 10456 12922
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10520 12238 10548 12854
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11694 10548 12038
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10612 10810 10640 14878
rect 10704 12209 10732 15014
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14278 10824 14758
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10888 13433 10916 19071
rect 10980 18766 11008 20198
rect 11164 19854 11192 20334
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11072 18873 11100 19246
rect 11164 18970 11192 19790
rect 11256 19378 11284 19858
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11256 19174 11284 19314
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11058 18864 11114 18873
rect 11058 18799 11114 18808
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11072 18154 11100 18566
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 17338 11008 18022
rect 11058 17912 11114 17921
rect 11058 17847 11060 17856
rect 11112 17847 11114 17856
rect 11060 17818 11112 17824
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11256 17202 11284 19110
rect 11348 18902 11376 21916
rect 11336 18896 11388 18902
rect 11336 18838 11388 18844
rect 11532 18834 11560 22052
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11794 19272 11850 19281
rect 11794 19207 11796 19216
rect 11848 19207 11850 19216
rect 11796 19178 11848 19184
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11900 18154 11928 18838
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11348 17338 11376 17478
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11334 17232 11390 17241
rect 11244 17196 11296 17202
rect 11334 17167 11390 17176
rect 11244 17138 11296 17144
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11256 16794 11284 16934
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11256 16250 11284 16730
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 10980 15026 11008 15574
rect 11164 15502 11192 16050
rect 11348 15978 11376 17167
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11164 15162 11192 15438
rect 11334 15192 11390 15201
rect 11152 15156 11204 15162
rect 11334 15127 11390 15136
rect 11152 15098 11204 15104
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 11164 14618 11192 15098
rect 11244 14884 11296 14890
rect 11244 14826 11296 14832
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 10980 14074 11008 14554
rect 11256 14498 11284 14826
rect 11164 14470 11284 14498
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10874 13424 10930 13433
rect 10874 13359 10930 13368
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 12345 10824 13126
rect 11058 12472 11114 12481
rect 11058 12407 11114 12416
rect 10782 12336 10838 12345
rect 10782 12271 10838 12280
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10690 12200 10746 12209
rect 10690 12135 10746 12144
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10428 9722 10456 10066
rect 10704 9722 10732 12038
rect 10888 11898 10916 12242
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10198 10824 10950
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10796 9586 10824 10134
rect 10888 9625 10916 11834
rect 10980 11762 11008 12242
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11072 11354 11100 12407
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11164 11268 11192 14470
rect 11348 12481 11376 15127
rect 11334 12472 11390 12481
rect 11334 12407 11390 12416
rect 11334 12336 11390 12345
rect 11334 12271 11390 12280
rect 11164 11240 11284 11268
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10968 10804 11020 10810
rect 11072 10792 11100 11154
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11164 10810 11192 11018
rect 11020 10764 11100 10792
rect 11152 10804 11204 10810
rect 10968 10746 11020 10752
rect 11152 10746 11204 10752
rect 10980 10266 11008 10746
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11164 10146 11192 10746
rect 10980 10118 11192 10146
rect 10980 9654 11008 10118
rect 10968 9648 11020 9654
rect 10874 9616 10930 9625
rect 10784 9580 10836 9586
rect 10968 9590 11020 9596
rect 10874 9551 10930 9560
rect 10784 9522 10836 9528
rect 10888 7954 10916 9551
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10888 7546 10916 7890
rect 11072 7546 11100 7890
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10244 3505 10272 3538
rect 10230 3496 10286 3505
rect 10230 3431 10286 3440
rect 10244 2650 10272 3431
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10428 2514 10456 7278
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 6866 11008 7142
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 5914 11008 6802
rect 11072 6662 11100 7482
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11164 6458 11192 6802
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11072 5817 11100 6054
rect 11058 5808 11114 5817
rect 11164 5794 11192 6394
rect 11256 5914 11284 11240
rect 11348 11014 11376 12271
rect 11440 11665 11468 18022
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11520 17264 11572 17270
rect 11520 17206 11572 17212
rect 11532 16658 11560 17206
rect 11900 17202 11928 17478
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11532 16250 11560 16594
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11532 14482 11560 16186
rect 11900 16114 11928 16594
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11532 14074 11560 14418
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11532 12986 11560 14010
rect 11808 13870 11836 14418
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11532 11898 11560 12922
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11426 11656 11482 11665
rect 11426 11591 11482 11600
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11440 11286 11468 11494
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11520 11348 11572 11354
rect 11992 11336 12020 24550
rect 12084 24154 12112 28886
rect 12636 28744 12664 32166
rect 12268 28716 12664 28744
rect 12162 27976 12218 27985
rect 12162 27911 12218 27920
rect 12176 24682 12204 27911
rect 12164 24676 12216 24682
rect 12164 24618 12216 24624
rect 12084 24126 12204 24154
rect 12072 20324 12124 20330
rect 12072 20266 12124 20272
rect 12084 18970 12112 20266
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12176 17241 12204 24126
rect 12268 23322 12296 28716
rect 12622 28656 12678 28665
rect 12622 28591 12678 28600
rect 12636 25498 12664 28591
rect 13004 28121 13032 39520
rect 12990 28112 13046 28121
rect 12990 28047 13046 28056
rect 12900 27328 12952 27334
rect 12900 27270 12952 27276
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12636 25378 12664 25434
rect 12532 25356 12584 25362
rect 12636 25350 12756 25378
rect 12532 25298 12584 25304
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12360 24698 12388 25094
rect 12544 24954 12572 25298
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 12360 24670 12480 24698
rect 12452 24070 12480 24670
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12360 23594 12388 24006
rect 12532 23860 12584 23866
rect 12532 23802 12584 23808
rect 12438 23760 12494 23769
rect 12438 23695 12440 23704
rect 12492 23695 12494 23704
rect 12440 23666 12492 23672
rect 12438 23624 12494 23633
rect 12348 23588 12400 23594
rect 12438 23559 12494 23568
rect 12348 23530 12400 23536
rect 12452 23526 12480 23559
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 12544 23254 12572 23802
rect 12636 23662 12664 24550
rect 12728 24410 12756 25350
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12728 23594 12756 24006
rect 12716 23588 12768 23594
rect 12716 23530 12768 23536
rect 12624 23520 12676 23526
rect 12676 23468 12756 23474
rect 12624 23462 12756 23468
rect 12636 23446 12756 23462
rect 12532 23248 12584 23254
rect 12532 23190 12584 23196
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22778 12480 23122
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12544 22710 12572 23190
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12440 21344 12492 21350
rect 12268 21292 12440 21298
rect 12268 21286 12492 21292
rect 12268 21270 12480 21286
rect 12268 18222 12296 21270
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12544 20466 12572 20742
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12360 20262 12388 20334
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12360 20058 12388 20198
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12452 19961 12480 20198
rect 12438 19952 12494 19961
rect 12438 19887 12494 19896
rect 12544 19514 12572 20402
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12360 18290 12388 18770
rect 12544 18766 12572 19314
rect 12622 19272 12678 19281
rect 12622 19207 12624 19216
rect 12676 19207 12678 19216
rect 12624 19178 12676 19184
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12162 17232 12218 17241
rect 12072 17196 12124 17202
rect 12728 17218 12756 23446
rect 12820 21049 12848 26862
rect 12912 25498 12940 27270
rect 13372 26926 13400 39520
rect 13634 36680 13690 36689
rect 13634 36615 13690 36624
rect 13450 35728 13506 35737
rect 13450 35663 13506 35672
rect 13464 34542 13492 35663
rect 13648 34746 13676 36615
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 13452 34536 13504 34542
rect 13452 34478 13504 34484
rect 13452 34060 13504 34066
rect 13452 34002 13504 34008
rect 13464 33658 13492 34002
rect 13452 33652 13504 33658
rect 13452 33594 13504 33600
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 12912 25294 12940 25434
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 12912 24886 12940 25230
rect 13176 24948 13228 24954
rect 13176 24890 13228 24896
rect 12900 24880 12952 24886
rect 12900 24822 12952 24828
rect 12912 24410 12940 24822
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 12912 23798 12940 24346
rect 12900 23792 12952 23798
rect 12900 23734 12952 23740
rect 13004 23644 13032 24550
rect 13188 24410 13216 24890
rect 13740 24721 13768 39520
rect 13912 37188 13964 37194
rect 13912 37130 13964 37136
rect 13924 28665 13952 37130
rect 14200 29889 14228 39520
rect 14568 37194 14596 39520
rect 14556 37188 14608 37194
rect 14556 37130 14608 37136
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14936 31822 14964 39520
rect 14924 31816 14976 31822
rect 14924 31758 14976 31764
rect 14740 31748 14792 31754
rect 14740 31690 14792 31696
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14186 29880 14242 29889
rect 14186 29815 14242 29824
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 13910 28656 13966 28665
rect 13910 28591 13966 28600
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 13726 24712 13782 24721
rect 13726 24647 13782 24656
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13004 23616 13124 23644
rect 12900 23316 12952 23322
rect 12900 23258 12952 23264
rect 12806 21040 12862 21049
rect 12806 20975 12862 20984
rect 12162 17167 12218 17176
rect 12544 17190 12756 17218
rect 12072 17138 12124 17144
rect 12084 16794 12112 17138
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12176 16674 12204 17070
rect 11520 11290 11572 11296
rect 11900 11308 12020 11336
rect 12084 16646 12204 16674
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11532 11234 11560 11290
rect 11440 11150 11468 11222
rect 11532 11206 11652 11234
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11348 10674 11376 10950
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11164 5766 11284 5794
rect 11058 5743 11114 5752
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10782 4856 10838 4865
rect 10782 4791 10838 4800
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10520 3534 10548 4082
rect 10612 3738 10640 4626
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10704 3913 10732 4558
rect 10690 3904 10746 3913
rect 10690 3839 10746 3848
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10690 3632 10746 3641
rect 10796 3618 10824 4791
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4282 10916 4558
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10888 3720 10916 4218
rect 11072 4185 11100 5238
rect 11164 5030 11192 5646
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11164 4282 11192 4966
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11256 4214 11284 5766
rect 11348 4486 11376 10474
rect 11440 10266 11468 11086
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11244 4208 11296 4214
rect 11058 4176 11114 4185
rect 11244 4150 11296 4156
rect 11058 4111 11114 4120
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10968 3732 11020 3738
rect 10888 3692 10968 3720
rect 10968 3674 11020 3680
rect 10796 3590 10916 3618
rect 10690 3567 10746 3576
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10598 3496 10654 3505
rect 10598 3431 10654 3440
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10612 480 10640 3431
rect 10704 2650 10732 3567
rect 10888 2666 10916 3590
rect 10692 2644 10744 2650
rect 10888 2638 11008 2666
rect 11072 2650 11100 3946
rect 11336 3936 11388 3942
rect 11334 3904 11336 3913
rect 11388 3904 11390 3913
rect 11334 3839 11390 3848
rect 11440 3754 11468 8230
rect 11532 6254 11560 10678
rect 11624 10538 11652 11206
rect 11900 10849 11928 11308
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11886 10840 11942 10849
rect 11886 10775 11942 10784
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11992 8294 12020 11154
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 12084 8090 12112 16646
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12162 13424 12218 13433
rect 12162 13359 12218 13368
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 7970 12204 13359
rect 12268 11218 12296 15846
rect 12348 13864 12400 13870
rect 12400 13812 12480 13818
rect 12348 13806 12480 13812
rect 12360 13790 12480 13806
rect 12452 12442 12480 13790
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12360 10606 12388 11086
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12440 10532 12492 10538
rect 12440 10474 12492 10480
rect 12452 9926 12480 10474
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12084 7942 12204 7970
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11532 5098 11560 5714
rect 11992 5710 12020 6598
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5370 12020 5646
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11612 5160 11664 5166
rect 11610 5128 11612 5137
rect 11664 5128 11666 5137
rect 11520 5092 11572 5098
rect 11610 5063 11666 5072
rect 11520 5034 11572 5040
rect 11532 4826 11560 5034
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11348 3726 11468 3754
rect 11164 3194 11192 3674
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11164 3058 11192 3130
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 10692 2586 10744 2592
rect 10980 480 11008 2638
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11164 2446 11192 2994
rect 11348 2802 11376 3726
rect 12084 3505 12112 7942
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12360 7410 12388 7686
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12452 6361 12480 9862
rect 12438 6352 12494 6361
rect 12438 6287 12494 6296
rect 12254 6216 12310 6225
rect 12254 6151 12310 6160
rect 12268 4842 12296 6151
rect 12544 5681 12572 17190
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12636 10742 12664 17002
rect 12714 13288 12770 13297
rect 12714 13223 12770 13232
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12728 7562 12756 13223
rect 12912 10538 12940 23258
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13004 19378 13032 19654
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 13004 10198 13032 10610
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 12728 7534 13032 7562
rect 12806 7440 12862 7449
rect 12806 7375 12862 7384
rect 12530 5672 12586 5681
rect 12530 5607 12586 5616
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12268 4814 12572 4842
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12070 3496 12126 3505
rect 12070 3431 12126 3440
rect 11328 2774 11376 2802
rect 11328 2666 11356 2774
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11328 2638 11376 2666
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11348 480 11376 2638
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 12084 2258 12112 2450
rect 12176 2378 12204 4626
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 12084 2230 12204 2258
rect 11796 1420 11848 1426
rect 11796 1362 11848 1368
rect 11808 480 11836 1362
rect 12176 480 12204 2230
rect 12268 1426 12296 4422
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12360 3738 12388 4150
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12452 3194 12480 4694
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12544 2990 12572 4814
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12636 4214 12664 4558
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12636 3641 12664 3946
rect 12622 3632 12678 3641
rect 12622 3567 12678 3576
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12530 2816 12586 2825
rect 12530 2751 12586 2760
rect 12256 1420 12308 1426
rect 12256 1362 12308 1368
rect 12544 480 12572 2751
rect 12728 2650 12756 4966
rect 12820 4026 12848 7375
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12912 4146 12940 4626
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12820 3998 12940 4026
rect 12912 2825 12940 3998
rect 13004 3942 13032 7534
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13096 2922 13124 23616
rect 13188 23526 13216 24210
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 13266 23760 13322 23769
rect 13266 23695 13268 23704
rect 13320 23695 13322 23704
rect 13268 23666 13320 23672
rect 13176 23520 13228 23526
rect 13176 23462 13228 23468
rect 13634 23352 13690 23361
rect 13634 23287 13690 23296
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13464 22098 13492 22918
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13464 21350 13492 22034
rect 13648 21962 13676 23287
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14752 22001 14780 31690
rect 15396 30297 15424 39520
rect 15764 33561 15792 39520
rect 15750 33552 15806 33561
rect 15750 33487 15806 33496
rect 15382 30288 15438 30297
rect 15382 30223 15438 30232
rect 14738 21992 14794 22001
rect 13636 21956 13688 21962
rect 14738 21927 14794 21936
rect 13636 21898 13688 21904
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13542 16688 13598 16697
rect 13542 16623 13598 16632
rect 13556 15026 13584 16623
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13924 10033 13952 18158
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15382 10160 15438 10169
rect 15382 10095 15438 10104
rect 13910 10024 13966 10033
rect 13910 9959 13966 9968
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14186 8936 14242 8945
rect 14186 8871 14242 8880
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13084 2916 13136 2922
rect 13084 2858 13136 2864
rect 13096 2825 13124 2858
rect 12898 2816 12954 2825
rect 12898 2751 12954 2760
rect 13082 2816 13138 2825
rect 13082 2751 13138 2760
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 13096 2514 13124 2586
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 13188 2446 13216 2994
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13280 2258 13308 8026
rect 13450 5672 13506 5681
rect 13450 5607 13506 5616
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13372 4049 13400 4558
rect 13358 4040 13414 4049
rect 13358 3975 13414 3984
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13004 2230 13308 2258
rect 13004 480 13032 2230
rect 13372 480 13400 3878
rect 13464 2650 13492 5607
rect 13726 2952 13782 2961
rect 13726 2887 13782 2896
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13740 480 13768 2887
rect 14200 480 14228 8871
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14922 3088 14978 3097
rect 14922 3023 14978 3032
rect 14646 2816 14702 2825
rect 14646 2751 14702 2760
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14660 1986 14688 2751
rect 14568 1958 14688 1986
rect 14568 480 14596 1958
rect 14936 480 14964 3023
rect 15396 480 15424 10095
rect 15764 480 15792 10542
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 1490 34856 1546 34912
rect 2042 33904 2098 33960
rect 2778 38936 2834 38992
rect 2594 35264 2650 35320
rect 2410 33088 2466 33144
rect 1674 32952 1730 33008
rect 2042 32952 2098 33008
rect 1674 31220 1676 31240
rect 1676 31220 1728 31240
rect 1728 31220 1730 31240
rect 1674 31184 1730 31220
rect 1582 30912 1638 30968
rect 1582 29960 1638 30016
rect 1582 28872 1638 28928
rect 1674 26968 1730 27024
rect 1582 24928 1638 24984
rect 2226 30640 2282 30696
rect 2042 29164 2098 29200
rect 2042 29144 2044 29164
rect 2044 29144 2096 29164
rect 2096 29144 2098 29164
rect 2502 24792 2558 24848
rect 1766 24112 1822 24168
rect 1582 22888 1638 22944
rect 1674 20984 1730 21040
rect 1582 18944 1638 19000
rect 1398 18828 1454 18864
rect 1398 18808 1400 18828
rect 1400 18808 1452 18828
rect 1452 18808 1454 18828
rect 2226 18148 2282 18184
rect 2226 18128 2228 18148
rect 2228 18128 2280 18148
rect 2280 18128 2282 18148
rect 1582 16904 1638 16960
rect 1674 14864 1730 14920
rect 2226 14884 2282 14920
rect 2226 14864 2228 14884
rect 2228 14864 2280 14884
rect 2280 14864 2282 14884
rect 1582 12960 1638 13016
rect 1674 12588 1676 12608
rect 1676 12588 1728 12608
rect 1728 12588 1730 12608
rect 1674 12552 1730 12588
rect 1582 10920 1638 10976
rect 2226 11500 2228 11520
rect 2228 11500 2280 11520
rect 2280 11500 2282 11520
rect 2226 11464 2282 11500
rect 2042 9596 2044 9616
rect 2044 9596 2096 9616
rect 2096 9596 2098 9616
rect 2042 9560 2098 9596
rect 1582 8880 1638 8936
rect 2502 7384 2558 7440
rect 2318 6976 2374 7032
rect 938 3032 994 3088
rect 1490 5752 1546 5808
rect 1582 4936 1638 4992
rect 2226 2916 2282 2952
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3422 36896 3478 36952
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3422 35672 3478 35728
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 4158 36760 4214 36816
rect 4250 35284 4306 35320
rect 4250 35264 4252 35284
rect 4252 35264 4304 35284
rect 4304 35264 4306 35284
rect 4250 34740 4306 34776
rect 4250 34720 4252 34740
rect 4252 34720 4304 34740
rect 4304 34720 4306 34740
rect 2778 29960 2834 30016
rect 4526 34584 4582 34640
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 4526 33904 4582 33960
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3330 32408 3386 32464
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3422 22616 3478 22672
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3146 20848 3202 20904
rect 2686 15544 2742 15600
rect 2226 2896 2228 2916
rect 2228 2896 2280 2916
rect 2280 2896 2282 2916
rect 2410 2644 2466 2680
rect 2410 2624 2412 2644
rect 2412 2624 2464 2644
rect 2464 2624 2466 2644
rect 2134 1400 2190 1456
rect 2594 2760 2650 2816
rect 2502 992 2558 1048
rect 3238 16768 3294 16824
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 4066 28056 4122 28112
rect 3974 20848 4030 20904
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 4526 25764 4582 25800
rect 4526 25744 4528 25764
rect 4528 25744 4580 25764
rect 4580 25744 4582 25764
rect 4710 25336 4766 25392
rect 4526 23160 4582 23216
rect 4986 33088 5042 33144
rect 5262 30776 5318 30832
rect 5078 30096 5134 30152
rect 4618 20984 4674 21040
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 4434 19352 4490 19408
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 4158 16788 4214 16824
rect 4158 16768 4160 16788
rect 4160 16768 4212 16788
rect 4212 16768 4214 16788
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 4250 13368 4306 13424
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3882 9596 3884 9616
rect 3884 9596 3936 9616
rect 3936 9596 3938 9616
rect 3882 9560 3938 9596
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3790 8356 3846 8392
rect 3790 8336 3792 8356
rect 3792 8336 3844 8356
rect 3844 8336 3846 8356
rect 3974 8336 4030 8392
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 4066 7248 4122 7304
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3054 5244 3056 5264
rect 3056 5244 3108 5264
rect 3108 5244 3110 5264
rect 3054 5208 3110 5244
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3882 4548 3938 4584
rect 3882 4528 3884 4548
rect 3884 4528 3936 4548
rect 3936 4528 3938 4548
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 4158 4392 4214 4448
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3882 2524 3884 2544
rect 3884 2524 3936 2544
rect 3936 2524 3938 2544
rect 3882 2488 3938 2524
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 5630 32272 5686 32328
rect 5538 28056 5594 28112
rect 4618 16496 4674 16552
rect 4434 14320 4490 14376
rect 4526 13912 4582 13968
rect 4894 12416 4950 12472
rect 5170 21412 5226 21448
rect 5170 21392 5172 21412
rect 5172 21392 5224 21412
rect 5224 21392 5226 21412
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 7286 36760 7342 36816
rect 7102 34720 7158 34776
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 5446 24692 5448 24712
rect 5448 24692 5500 24712
rect 5500 24692 5502 24712
rect 5446 24656 5502 24692
rect 5354 22072 5410 22128
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6550 32952 6606 33008
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6734 29008 6790 29064
rect 6918 30640 6974 30696
rect 7378 34584 7434 34640
rect 7838 34584 7894 34640
rect 7838 33496 7894 33552
rect 7746 33224 7802 33280
rect 7286 30932 7342 30968
rect 7286 30912 7288 30932
rect 7288 30912 7340 30932
rect 7340 30912 7342 30932
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 5998 24248 6054 24304
rect 5170 17176 5226 17232
rect 5446 21548 5502 21584
rect 5446 21528 5448 21548
rect 5448 21528 5500 21548
rect 5500 21528 5502 21548
rect 4894 12280 4950 12336
rect 4802 11464 4858 11520
rect 4710 9696 4766 9752
rect 4434 6196 4436 6216
rect 4436 6196 4488 6216
rect 4488 6196 4490 6216
rect 4434 6160 4490 6196
rect 4526 5208 4582 5264
rect 4342 3984 4398 4040
rect 4250 2760 4306 2816
rect 4986 7964 4988 7984
rect 4988 7964 5040 7984
rect 5040 7964 5042 7984
rect 4986 7928 5042 7964
rect 5630 17584 5686 17640
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6826 26968 6882 27024
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 7102 24792 7158 24848
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6182 22616 6238 22672
rect 5906 15680 5962 15736
rect 5906 15580 5908 15600
rect 5908 15580 5960 15600
rect 5960 15580 5962 15600
rect 5906 15544 5962 15580
rect 5538 12552 5594 12608
rect 5814 13776 5870 13832
rect 5814 12144 5870 12200
rect 5354 8880 5410 8936
rect 4986 7384 5042 7440
rect 4802 3984 4858 4040
rect 4618 2760 4674 2816
rect 4802 2760 4858 2816
rect 5078 6160 5134 6216
rect 5538 6568 5594 6624
rect 5078 4528 5134 4584
rect 5262 5616 5318 5672
rect 4710 2624 4766 2680
rect 5814 9424 5870 9480
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 7194 22652 7196 22672
rect 7196 22652 7248 22672
rect 7248 22652 7250 22672
rect 7194 22616 7250 22652
rect 6642 21664 6698 21720
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 7102 21528 7158 21584
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6734 18808 6790 18864
rect 7562 28736 7618 28792
rect 7562 28620 7618 28656
rect 7562 28600 7564 28620
rect 7564 28600 7616 28620
rect 7616 28600 7618 28620
rect 7470 28076 7526 28112
rect 7470 28056 7472 28076
rect 7472 28056 7524 28076
rect 7524 28056 7526 28076
rect 7838 26424 7894 26480
rect 7562 25608 7618 25664
rect 7562 23316 7618 23352
rect 7562 23296 7564 23316
rect 7564 23296 7616 23316
rect 7616 23296 7618 23316
rect 7470 21392 7526 21448
rect 7286 19216 7342 19272
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6182 15952 6238 16008
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6182 15544 6238 15600
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6182 14456 6238 14512
rect 6826 15816 6882 15872
rect 6734 13640 6790 13696
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 5998 11056 6054 11112
rect 7746 21292 7748 21312
rect 7748 21292 7800 21312
rect 7800 21292 7802 21312
rect 7746 21256 7802 21292
rect 8022 23160 8078 23216
rect 8206 27956 8208 27976
rect 8208 27956 8260 27976
rect 8260 27956 8262 27976
rect 8206 27920 8262 27956
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 9310 33904 9366 33960
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 9402 33088 9458 33144
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8758 32272 8814 32328
rect 9310 32308 9312 32328
rect 9312 32308 9364 32328
rect 9364 32308 9366 32328
rect 9310 32272 9366 32308
rect 8482 25744 8538 25800
rect 7654 19352 7710 19408
rect 7562 19080 7618 19136
rect 7194 15000 7250 15056
rect 7194 14728 7250 14784
rect 7654 16108 7710 16144
rect 7654 16088 7656 16108
rect 7656 16088 7708 16108
rect 7708 16088 7710 16108
rect 8206 21392 8262 21448
rect 8114 20984 8170 21040
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8758 27820 8760 27840
rect 8760 27820 8812 27840
rect 8812 27820 8814 27840
rect 8758 27784 8814 27820
rect 8666 24384 8722 24440
rect 8574 21664 8630 21720
rect 8942 29028 8998 29064
rect 8942 29008 8944 29028
rect 8944 29008 8996 29028
rect 8996 29008 8998 29028
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 9310 26968 9366 27024
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 9034 24112 9090 24168
rect 9310 24112 9366 24168
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 9218 23296 9274 23352
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8206 15852 8208 15872
rect 8208 15852 8260 15872
rect 8260 15852 8262 15872
rect 7470 13776 7526 13832
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6734 12552 6790 12608
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 5814 8336 5870 8392
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6918 9696 6974 9752
rect 5814 5072 5870 5128
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6182 6860 6238 6896
rect 6182 6840 6184 6860
rect 6184 6840 6236 6860
rect 6236 6840 6238 6860
rect 6642 6452 6698 6488
rect 6642 6432 6644 6452
rect 6644 6432 6696 6452
rect 6696 6432 6698 6452
rect 6642 6296 6698 6352
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6734 5616 6790 5672
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6182 3984 6238 4040
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 6826 4564 6828 4584
rect 6828 4564 6880 4584
rect 6880 4564 6882 4584
rect 6826 4528 6882 4564
rect 7010 4392 7066 4448
rect 7010 4120 7066 4176
rect 6826 3304 6882 3360
rect 6918 3032 6974 3088
rect 7562 8608 7618 8664
rect 7470 5752 7526 5808
rect 7470 4664 7526 4720
rect 7194 3712 7250 3768
rect 7102 1400 7158 1456
rect 7470 2488 7526 2544
rect 8206 15816 8262 15852
rect 9310 21256 9366 21312
rect 8206 15564 8262 15600
rect 8206 15544 8208 15564
rect 8208 15544 8260 15564
rect 8260 15544 8262 15564
rect 8114 13640 8170 13696
rect 8022 12824 8078 12880
rect 8022 11736 8078 11792
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 9310 18264 9366 18320
rect 9310 18028 9312 18048
rect 9312 18028 9364 18048
rect 9364 18028 9366 18048
rect 9310 17992 9366 18028
rect 9310 17856 9366 17912
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8206 11056 8262 11112
rect 8114 9016 8170 9072
rect 8206 8236 8208 8256
rect 8208 8236 8260 8256
rect 8260 8236 8262 8256
rect 8206 8200 8262 8236
rect 8482 11600 8538 11656
rect 8482 10240 8538 10296
rect 7930 6840 7986 6896
rect 8390 7928 8446 7984
rect 8114 7148 8116 7168
rect 8116 7148 8168 7168
rect 8168 7148 8170 7168
rect 8114 7112 8170 7148
rect 10046 34584 10102 34640
rect 10046 32408 10102 32464
rect 10138 31184 10194 31240
rect 10414 33360 10470 33416
rect 10322 33088 10378 33144
rect 10046 26968 10102 27024
rect 9678 26696 9734 26752
rect 9678 26424 9734 26480
rect 9678 24248 9734 24304
rect 9678 23704 9734 23760
rect 9586 23568 9642 23624
rect 9586 19352 9642 19408
rect 9586 18808 9642 18864
rect 10598 30912 10654 30968
rect 10874 33496 10930 33552
rect 10690 30776 10746 30832
rect 10506 27784 10562 27840
rect 10230 26560 10286 26616
rect 9862 25644 9864 25664
rect 9864 25644 9916 25664
rect 9916 25644 9918 25664
rect 9862 25608 9918 25644
rect 10046 25372 10048 25392
rect 10048 25372 10100 25392
rect 10100 25372 10102 25392
rect 10046 25336 10102 25372
rect 9862 23704 9918 23760
rect 10046 22092 10102 22128
rect 10046 22072 10048 22092
rect 10048 22072 10100 22092
rect 10100 22072 10102 22092
rect 9770 21120 9826 21176
rect 9862 20848 9918 20904
rect 9770 20712 9826 20768
rect 9586 17856 9642 17912
rect 9954 19916 10010 19952
rect 9954 19896 9956 19916
rect 9956 19896 10008 19916
rect 10008 19896 10010 19916
rect 10690 25608 10746 25664
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8850 12588 8852 12608
rect 8852 12588 8904 12608
rect 8904 12588 8906 12608
rect 8850 12552 8906 12588
rect 8850 12280 8906 12336
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8574 8608 8630 8664
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8942 10104 8998 10160
rect 9678 14728 9734 14784
rect 9494 13776 9550 13832
rect 9402 10784 9458 10840
rect 9402 10240 9458 10296
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 9310 9560 9366 9616
rect 9126 9444 9182 9480
rect 9126 9424 9128 9444
rect 9128 9424 9180 9444
rect 9180 9424 9182 9444
rect 8206 6432 8262 6488
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8942 7420 8944 7440
rect 8944 7420 8996 7440
rect 8996 7420 8998 7440
rect 8942 7384 8998 7420
rect 8022 6160 8078 6216
rect 8574 6568 8630 6624
rect 7746 5752 7802 5808
rect 8022 3848 8078 3904
rect 7838 3576 7894 3632
rect 8482 4528 8538 4584
rect 8390 3984 8446 4040
rect 9218 6840 9274 6896
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 10046 18128 10102 18184
rect 9954 16088 10010 16144
rect 9862 15952 9918 16008
rect 9862 15000 9918 15056
rect 11150 30232 11206 30288
rect 11058 23316 11114 23352
rect 11058 23296 11060 23316
rect 11060 23296 11112 23316
rect 11112 23296 11114 23316
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 12162 33380 12218 33416
rect 12162 33360 12164 33380
rect 12164 33360 12216 33380
rect 12216 33360 12218 33380
rect 11886 32272 11942 32328
rect 12070 32272 12126 32328
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11426 25608 11482 25664
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 12898 33496 12954 33552
rect 12438 30096 12494 30152
rect 12438 29824 12494 29880
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11518 24112 11574 24168
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 10414 16496 10470 16552
rect 10138 15544 10194 15600
rect 10414 15544 10470 15600
rect 10046 14864 10102 14920
rect 10598 17584 10654 17640
rect 10874 19080 10930 19136
rect 10782 17992 10838 18048
rect 10782 15136 10838 15192
rect 10138 14320 10194 14376
rect 10230 13912 10286 13968
rect 9770 9016 9826 9072
rect 9402 6840 9458 6896
rect 9310 5072 9366 5128
rect 8758 4004 8814 4040
rect 8758 3984 8760 4004
rect 8760 3984 8812 4004
rect 8812 3984 8814 4004
rect 8758 3712 8814 3768
rect 8482 3032 8538 3088
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 9494 6060 9496 6080
rect 9496 6060 9548 6080
rect 9548 6060 9550 6080
rect 9494 6024 9550 6060
rect 9678 7248 9734 7304
rect 10046 11736 10102 11792
rect 10322 13640 10378 13696
rect 10322 13368 10378 13424
rect 9770 5208 9826 5264
rect 9862 4664 9918 4720
rect 9678 3712 9734 3768
rect 9494 2760 9550 2816
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 10230 8200 10286 8256
rect 10138 7112 10194 7168
rect 11058 18808 11114 18864
rect 11058 17876 11114 17912
rect 11058 17856 11060 17876
rect 11060 17856 11112 17876
rect 11112 17856 11114 17876
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11794 19236 11850 19272
rect 11794 19216 11796 19236
rect 11796 19216 11848 19236
rect 11848 19216 11850 19236
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11334 17176 11390 17232
rect 11334 15136 11390 15192
rect 10874 13368 10930 13424
rect 11058 12416 11114 12472
rect 10782 12280 10838 12336
rect 10690 12144 10746 12200
rect 11334 12416 11390 12472
rect 11334 12280 11390 12336
rect 10874 9560 10930 9616
rect 10230 3440 10286 3496
rect 11058 5752 11114 5808
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11426 11600 11482 11656
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 12162 27920 12218 27976
rect 12622 28600 12678 28656
rect 12990 28056 13046 28112
rect 12438 23724 12494 23760
rect 12438 23704 12440 23724
rect 12440 23704 12492 23724
rect 12492 23704 12494 23724
rect 12438 23568 12494 23624
rect 12438 19896 12494 19952
rect 12622 19236 12678 19272
rect 12622 19216 12624 19236
rect 12624 19216 12676 19236
rect 12676 19216 12678 19236
rect 12162 17176 12218 17232
rect 13634 36624 13690 36680
rect 13450 35672 13506 35728
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14186 29824 14242 29880
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 13910 28600 13966 28656
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 13726 24656 13782 24712
rect 12806 20984 12862 21040
rect 10782 4800 10838 4856
rect 10690 3848 10746 3904
rect 10690 3576 10746 3632
rect 11058 4120 11114 4176
rect 10598 3440 10654 3496
rect 11334 3884 11336 3904
rect 11336 3884 11388 3904
rect 11388 3884 11390 3904
rect 11334 3848 11390 3884
rect 11886 10784 11942 10840
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 12162 13368 12218 13424
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11610 5108 11612 5128
rect 11612 5108 11664 5128
rect 11664 5108 11666 5128
rect 11610 5072 11666 5108
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 12438 6296 12494 6352
rect 12254 6160 12310 6216
rect 12714 13232 12770 13288
rect 12806 7384 12862 7440
rect 12530 5616 12586 5672
rect 12070 3440 12126 3496
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12622 3576 12678 3632
rect 12530 2760 12586 2816
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 13266 23724 13322 23760
rect 13266 23704 13268 23724
rect 13268 23704 13320 23724
rect 13320 23704 13322 23724
rect 13634 23296 13690 23352
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 15750 33496 15806 33552
rect 15382 30232 15438 30288
rect 14738 21936 14794 21992
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 13542 16632 13598 16688
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 15382 10104 15438 10160
rect 13910 9968 13966 10024
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14186 8880 14242 8936
rect 12898 2760 12954 2816
rect 13082 2760 13138 2816
rect 13450 5616 13506 5672
rect 13358 3984 13414 4040
rect 13726 2896 13782 2952
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14922 3032 14978 3088
rect 14646 2760 14702 2816
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
<< metal3 >>
rect 0 38994 480 39024
rect 2773 38994 2839 38997
rect 0 38992 2839 38994
rect 0 38936 2778 38992
rect 2834 38936 2839 38992
rect 0 38934 2839 38936
rect 0 38904 480 38934
rect 2773 38931 2839 38934
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 0 36954 480 36984
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 3417 36954 3483 36957
rect 0 36952 3483 36954
rect 0 36896 3422 36952
rect 3478 36896 3483 36952
rect 0 36894 3483 36896
rect 0 36864 480 36894
rect 3417 36891 3483 36894
rect 4153 36818 4219 36821
rect 7281 36818 7347 36821
rect 4153 36816 7347 36818
rect 4153 36760 4158 36816
rect 4214 36760 7286 36816
rect 7342 36760 7347 36816
rect 4153 36758 7347 36760
rect 4153 36755 4219 36758
rect 7281 36755 7347 36758
rect 13629 36682 13695 36685
rect 15520 36682 16000 36712
rect 13629 36680 16000 36682
rect 13629 36624 13634 36680
rect 13690 36624 16000 36680
rect 13629 36622 16000 36624
rect 13629 36619 13695 36622
rect 15520 36592 16000 36622
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 3417 35730 3483 35733
rect 13445 35730 13511 35733
rect 3417 35728 13511 35730
rect 3417 35672 3422 35728
rect 3478 35672 13450 35728
rect 13506 35672 13511 35728
rect 3417 35670 13511 35672
rect 3417 35667 3483 35670
rect 13445 35667 13511 35670
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 2589 35322 2655 35325
rect 4245 35322 4311 35325
rect 2589 35320 4311 35322
rect 2589 35264 2594 35320
rect 2650 35264 4250 35320
rect 4306 35264 4311 35320
rect 2589 35262 4311 35264
rect 2589 35259 2655 35262
rect 4245 35259 4311 35262
rect 0 34914 480 34944
rect 1485 34914 1551 34917
rect 0 34912 1551 34914
rect 0 34856 1490 34912
rect 1546 34856 1551 34912
rect 0 34854 1551 34856
rect 0 34824 480 34854
rect 1485 34851 1551 34854
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 4245 34778 4311 34781
rect 7097 34778 7163 34781
rect 4245 34776 7163 34778
rect 4245 34720 4250 34776
rect 4306 34720 7102 34776
rect 7158 34720 7163 34776
rect 4245 34718 7163 34720
rect 4245 34715 4311 34718
rect 7097 34715 7163 34718
rect 4521 34642 4587 34645
rect 7373 34642 7439 34645
rect 4521 34640 7439 34642
rect 4521 34584 4526 34640
rect 4582 34584 7378 34640
rect 7434 34584 7439 34640
rect 4521 34582 7439 34584
rect 4521 34579 4587 34582
rect 7373 34579 7439 34582
rect 7833 34642 7899 34645
rect 10041 34642 10107 34645
rect 7833 34640 10107 34642
rect 7833 34584 7838 34640
rect 7894 34584 10046 34640
rect 10102 34584 10107 34640
rect 7833 34582 10107 34584
rect 7833 34579 7899 34582
rect 10041 34579 10107 34582
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 2037 33962 2103 33965
rect 4521 33962 4587 33965
rect 9305 33962 9371 33965
rect 2037 33960 9371 33962
rect 2037 33904 2042 33960
rect 2098 33904 4526 33960
rect 4582 33904 9310 33960
rect 9366 33904 9371 33960
rect 2037 33902 9371 33904
rect 2037 33899 2103 33902
rect 4521 33899 4587 33902
rect 9305 33899 9371 33902
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 7833 33554 7899 33557
rect 10869 33554 10935 33557
rect 7833 33552 10935 33554
rect 7833 33496 7838 33552
rect 7894 33496 10874 33552
rect 10930 33496 10935 33552
rect 7833 33494 10935 33496
rect 7833 33491 7899 33494
rect 10869 33491 10935 33494
rect 12893 33554 12959 33557
rect 15745 33554 15811 33557
rect 12893 33552 15811 33554
rect 12893 33496 12898 33552
rect 12954 33496 15750 33552
rect 15806 33496 15811 33552
rect 12893 33494 15811 33496
rect 12893 33491 12959 33494
rect 15745 33491 15811 33494
rect 10409 33418 10475 33421
rect 12157 33418 12223 33421
rect 10409 33416 12223 33418
rect 10409 33360 10414 33416
rect 10470 33360 12162 33416
rect 12218 33360 12223 33416
rect 10409 33358 12223 33360
rect 10409 33355 10475 33358
rect 12157 33355 12223 33358
rect 7741 33282 7807 33285
rect 7741 33280 9506 33282
rect 7741 33224 7746 33280
rect 7802 33224 9506 33280
rect 7741 33222 9506 33224
rect 7741 33219 7807 33222
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 9446 33149 9506 33222
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 2405 33146 2471 33149
rect 4981 33146 5047 33149
rect 9397 33146 9506 33149
rect 10317 33146 10383 33149
rect 2405 33144 5047 33146
rect 2405 33088 2410 33144
rect 2466 33088 4986 33144
rect 5042 33088 5047 33144
rect 2405 33086 5047 33088
rect 9316 33144 10383 33146
rect 9316 33088 9402 33144
rect 9458 33088 10322 33144
rect 10378 33088 10383 33144
rect 9316 33086 10383 33088
rect 2405 33083 2471 33086
rect 4981 33083 5047 33086
rect 9397 33083 9463 33086
rect 10317 33083 10383 33086
rect 0 33010 480 33040
rect 1669 33010 1735 33013
rect 0 33008 1735 33010
rect 0 32952 1674 33008
rect 1730 32952 1735 33008
rect 0 32950 1735 32952
rect 0 32920 480 32950
rect 1669 32947 1735 32950
rect 2037 33010 2103 33013
rect 6545 33010 6611 33013
rect 2037 33008 6611 33010
rect 2037 32952 2042 33008
rect 2098 32952 6550 33008
rect 6606 32952 6611 33008
rect 2037 32950 6611 32952
rect 2037 32947 2103 32950
rect 6545 32947 6611 32950
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 3325 32466 3391 32469
rect 10041 32466 10107 32469
rect 3325 32464 10107 32466
rect 3325 32408 3330 32464
rect 3386 32408 10046 32464
rect 10102 32408 10107 32464
rect 3325 32406 10107 32408
rect 3325 32403 3391 32406
rect 10041 32403 10107 32406
rect 5625 32330 5691 32333
rect 8753 32330 8819 32333
rect 5625 32328 8819 32330
rect 5625 32272 5630 32328
rect 5686 32272 8758 32328
rect 8814 32272 8819 32328
rect 5625 32270 8819 32272
rect 5625 32267 5691 32270
rect 8753 32267 8819 32270
rect 9305 32330 9371 32333
rect 11881 32330 11947 32333
rect 12065 32330 12131 32333
rect 9305 32328 12131 32330
rect 9305 32272 9310 32328
rect 9366 32272 11886 32328
rect 11942 32272 12070 32328
rect 12126 32272 12131 32328
rect 9305 32270 12131 32272
rect 9305 32267 9371 32270
rect 11881 32267 11947 32270
rect 12065 32267 12131 32270
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 1669 31242 1735 31245
rect 10133 31242 10199 31245
rect 1669 31240 10199 31242
rect 1669 31184 1674 31240
rect 1730 31184 10138 31240
rect 10194 31184 10199 31240
rect 1669 31182 10199 31184
rect 1669 31179 1735 31182
rect 10133 31179 10199 31182
rect 6277 31040 6597 31041
rect 0 30970 480 31000
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 1577 30970 1643 30973
rect 0 30968 1643 30970
rect 0 30912 1582 30968
rect 1638 30912 1643 30968
rect 0 30910 1643 30912
rect 0 30880 480 30910
rect 1577 30907 1643 30910
rect 7281 30970 7347 30973
rect 10593 30970 10659 30973
rect 7281 30968 10659 30970
rect 7281 30912 7286 30968
rect 7342 30912 10598 30968
rect 10654 30912 10659 30968
rect 7281 30910 10659 30912
rect 7281 30907 7347 30910
rect 10593 30907 10659 30910
rect 5257 30834 5323 30837
rect 10685 30834 10751 30837
rect 5257 30832 10751 30834
rect 5257 30776 5262 30832
rect 5318 30776 10690 30832
rect 10746 30776 10751 30832
rect 5257 30774 10751 30776
rect 5257 30771 5323 30774
rect 10685 30771 10751 30774
rect 2221 30698 2287 30701
rect 6913 30698 6979 30701
rect 2221 30696 6979 30698
rect 2221 30640 2226 30696
rect 2282 30640 6918 30696
rect 6974 30640 6979 30696
rect 2221 30638 6979 30640
rect 2221 30635 2287 30638
rect 6913 30635 6979 30638
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 11145 30290 11211 30293
rect 15377 30290 15443 30293
rect 11145 30288 15443 30290
rect 11145 30232 11150 30288
rect 11206 30232 15382 30288
rect 15438 30232 15443 30288
rect 11145 30230 15443 30232
rect 11145 30227 11211 30230
rect 15377 30227 15443 30230
rect 5073 30154 5139 30157
rect 12433 30154 12499 30157
rect 5073 30152 12499 30154
rect 5073 30096 5078 30152
rect 5134 30096 12438 30152
rect 12494 30096 12499 30152
rect 5073 30094 12499 30096
rect 5073 30091 5139 30094
rect 12433 30091 12499 30094
rect 1577 30018 1643 30021
rect 2773 30018 2839 30021
rect 15520 30018 16000 30048
rect 1577 30016 2839 30018
rect 1577 29960 1582 30016
rect 1638 29960 2778 30016
rect 2834 29960 2839 30016
rect 1577 29958 2839 29960
rect 1577 29955 1643 29958
rect 2773 29955 2839 29958
rect 12022 29958 16000 30018
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 2037 29202 2103 29205
rect 12022 29202 12082 29958
rect 15520 29928 16000 29958
rect 12433 29882 12499 29885
rect 14181 29882 14247 29885
rect 12433 29880 14247 29882
rect 12433 29824 12438 29880
rect 12494 29824 14186 29880
rect 14242 29824 14247 29880
rect 12433 29822 14247 29824
rect 12433 29819 12499 29822
rect 14181 29819 14247 29822
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 2037 29200 12082 29202
rect 2037 29144 2042 29200
rect 2098 29144 12082 29200
rect 2037 29142 12082 29144
rect 2037 29139 2103 29142
rect 6729 29066 6795 29069
rect 8937 29066 9003 29069
rect 6729 29064 9003 29066
rect 6729 29008 6734 29064
rect 6790 29008 8942 29064
rect 8998 29008 9003 29064
rect 6729 29006 9003 29008
rect 6729 29003 6795 29006
rect 8937 29003 9003 29006
rect 0 28930 480 28960
rect 1577 28930 1643 28933
rect 0 28928 1643 28930
rect 0 28872 1582 28928
rect 1638 28872 1643 28928
rect 0 28870 1643 28872
rect 0 28840 480 28870
rect 1577 28867 1643 28870
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 7557 28794 7623 28797
rect 8150 28794 8156 28796
rect 7557 28792 8156 28794
rect 7557 28736 7562 28792
rect 7618 28736 8156 28792
rect 7557 28734 8156 28736
rect 7557 28731 7623 28734
rect 8150 28732 8156 28734
rect 8220 28732 8226 28796
rect 7557 28658 7623 28661
rect 12617 28658 12683 28661
rect 13905 28658 13971 28661
rect 7557 28656 13971 28658
rect 7557 28600 7562 28656
rect 7618 28600 12622 28656
rect 12678 28600 13910 28656
rect 13966 28600 13971 28656
rect 7557 28598 13971 28600
rect 7557 28595 7623 28598
rect 12617 28595 12683 28598
rect 13905 28595 13971 28598
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 4061 28114 4127 28117
rect 5533 28114 5599 28117
rect 4061 28112 5599 28114
rect 4061 28056 4066 28112
rect 4122 28056 5538 28112
rect 5594 28056 5599 28112
rect 4061 28054 5599 28056
rect 4061 28051 4127 28054
rect 5533 28051 5599 28054
rect 7465 28114 7531 28117
rect 12985 28114 13051 28117
rect 7465 28112 13051 28114
rect 7465 28056 7470 28112
rect 7526 28056 12990 28112
rect 13046 28056 13051 28112
rect 7465 28054 13051 28056
rect 7465 28051 7531 28054
rect 12985 28051 13051 28054
rect 8201 27978 8267 27981
rect 12157 27978 12223 27981
rect 8201 27976 12223 27978
rect 8201 27920 8206 27976
rect 8262 27920 12162 27976
rect 12218 27920 12223 27976
rect 8201 27918 12223 27920
rect 8201 27915 8267 27918
rect 12157 27915 12223 27918
rect 8753 27842 8819 27845
rect 10501 27842 10567 27845
rect 8753 27840 10567 27842
rect 8753 27784 8758 27840
rect 8814 27784 10506 27840
rect 10562 27784 10567 27840
rect 8753 27782 10567 27784
rect 8753 27779 8819 27782
rect 10501 27779 10567 27782
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 0 27026 480 27056
rect 1669 27026 1735 27029
rect 0 27024 1735 27026
rect 0 26968 1674 27024
rect 1730 26968 1735 27024
rect 0 26966 1735 26968
rect 0 26936 480 26966
rect 1669 26963 1735 26966
rect 6821 27026 6887 27029
rect 9305 27026 9371 27029
rect 6821 27024 9371 27026
rect 6821 26968 6826 27024
rect 6882 26968 9310 27024
rect 9366 26968 9371 27024
rect 6821 26966 9371 26968
rect 6821 26963 6887 26966
rect 9305 26963 9371 26966
rect 9806 26964 9812 27028
rect 9876 27026 9882 27028
rect 10041 27026 10107 27029
rect 9876 27024 10107 27026
rect 9876 26968 10046 27024
rect 10102 26968 10107 27024
rect 9876 26966 10107 26968
rect 9876 26964 9882 26966
rect 10041 26963 10107 26966
rect 9673 26754 9739 26757
rect 9673 26752 10242 26754
rect 9673 26696 9678 26752
rect 9734 26696 10242 26752
rect 9673 26694 10242 26696
rect 9673 26691 9739 26694
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 10182 26621 10242 26694
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 10182 26616 10291 26621
rect 10182 26560 10230 26616
rect 10286 26560 10291 26616
rect 10182 26558 10291 26560
rect 10225 26555 10291 26558
rect 7833 26482 7899 26485
rect 9673 26482 9739 26485
rect 7833 26480 9739 26482
rect 7833 26424 7838 26480
rect 7894 26424 9678 26480
rect 9734 26424 9739 26480
rect 7833 26422 9739 26424
rect 7833 26419 7899 26422
rect 9673 26419 9739 26422
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 4521 25802 4587 25805
rect 8477 25802 8543 25805
rect 4521 25800 8543 25802
rect 4521 25744 4526 25800
rect 4582 25744 8482 25800
rect 8538 25744 8543 25800
rect 4521 25742 8543 25744
rect 4521 25739 4587 25742
rect 8477 25739 8543 25742
rect 7557 25666 7623 25669
rect 9857 25666 9923 25669
rect 10685 25666 10751 25669
rect 11421 25666 11487 25669
rect 7557 25664 11487 25666
rect 7557 25608 7562 25664
rect 7618 25608 9862 25664
rect 9918 25608 10690 25664
rect 10746 25608 11426 25664
rect 11482 25608 11487 25664
rect 7557 25606 11487 25608
rect 7557 25603 7623 25606
rect 9857 25603 9923 25606
rect 10685 25603 10751 25606
rect 11421 25603 11487 25606
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 4705 25394 4771 25397
rect 10041 25394 10107 25397
rect 4705 25392 10107 25394
rect 4705 25336 4710 25392
rect 4766 25336 10046 25392
rect 10102 25336 10107 25392
rect 4705 25334 10107 25336
rect 4705 25331 4771 25334
rect 10041 25331 10107 25334
rect 3610 25056 3930 25057
rect 0 24986 480 25016
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 1577 24986 1643 24989
rect 0 24984 1643 24986
rect 0 24928 1582 24984
rect 1638 24928 1643 24984
rect 0 24926 1643 24928
rect 0 24896 480 24926
rect 1577 24923 1643 24926
rect 2497 24850 2563 24853
rect 7097 24850 7163 24853
rect 2497 24848 7163 24850
rect 2497 24792 2502 24848
rect 2558 24792 7102 24848
rect 7158 24792 7163 24848
rect 2497 24790 7163 24792
rect 2497 24787 2563 24790
rect 7097 24787 7163 24790
rect 5441 24714 5507 24717
rect 13721 24714 13787 24717
rect 5441 24712 13787 24714
rect 5441 24656 5446 24712
rect 5502 24656 13726 24712
rect 13782 24656 13787 24712
rect 5441 24654 13787 24656
rect 5441 24651 5507 24654
rect 13721 24651 13787 24654
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 8661 24442 8727 24445
rect 9438 24442 9444 24444
rect 8661 24440 9444 24442
rect 8661 24384 8666 24440
rect 8722 24384 9444 24440
rect 8661 24382 9444 24384
rect 8661 24379 8727 24382
rect 9438 24380 9444 24382
rect 9508 24380 9514 24444
rect 5993 24306 6059 24309
rect 9673 24306 9739 24309
rect 5993 24304 9739 24306
rect 5993 24248 5998 24304
rect 6054 24248 9678 24304
rect 9734 24248 9739 24304
rect 5993 24246 9739 24248
rect 5993 24243 6059 24246
rect 9673 24243 9739 24246
rect 1761 24170 1827 24173
rect 9029 24170 9095 24173
rect 1761 24168 9095 24170
rect 1761 24112 1766 24168
rect 1822 24112 9034 24168
rect 9090 24112 9095 24168
rect 1761 24110 9095 24112
rect 1761 24107 1827 24110
rect 9029 24107 9095 24110
rect 9305 24170 9371 24173
rect 11513 24170 11579 24173
rect 9305 24168 11579 24170
rect 9305 24112 9310 24168
rect 9366 24112 11518 24168
rect 11574 24112 11579 24168
rect 9305 24110 11579 24112
rect 9305 24107 9371 24110
rect 11513 24107 11579 24110
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 9673 23762 9739 23765
rect 9857 23762 9923 23765
rect 9673 23760 9923 23762
rect 9673 23704 9678 23760
rect 9734 23704 9862 23760
rect 9918 23704 9923 23760
rect 9673 23702 9923 23704
rect 9673 23699 9739 23702
rect 9857 23699 9923 23702
rect 12433 23762 12499 23765
rect 13261 23762 13327 23765
rect 12433 23760 13327 23762
rect 12433 23704 12438 23760
rect 12494 23704 13266 23760
rect 13322 23704 13327 23760
rect 12433 23702 13327 23704
rect 12433 23699 12499 23702
rect 13261 23699 13327 23702
rect 9581 23626 9647 23629
rect 12433 23626 12499 23629
rect 9581 23624 12499 23626
rect 9581 23568 9586 23624
rect 9642 23568 12438 23624
rect 12494 23568 12499 23624
rect 9581 23566 12499 23568
rect 9581 23563 9647 23566
rect 12433 23563 12499 23566
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 7557 23354 7623 23357
rect 9213 23354 9279 23357
rect 11053 23354 11119 23357
rect 7557 23352 11119 23354
rect 7557 23296 7562 23352
rect 7618 23296 9218 23352
rect 9274 23296 11058 23352
rect 11114 23296 11119 23352
rect 7557 23294 11119 23296
rect 7557 23291 7623 23294
rect 9213 23291 9279 23294
rect 11053 23291 11119 23294
rect 13629 23354 13695 23357
rect 15520 23354 16000 23384
rect 13629 23352 16000 23354
rect 13629 23296 13634 23352
rect 13690 23296 16000 23352
rect 13629 23294 16000 23296
rect 13629 23291 13695 23294
rect 15520 23264 16000 23294
rect 4521 23218 4587 23221
rect 8017 23218 8083 23221
rect 4521 23216 8083 23218
rect 4521 23160 4526 23216
rect 4582 23160 8022 23216
rect 8078 23160 8083 23216
rect 4521 23158 8083 23160
rect 4521 23155 4587 23158
rect 8017 23155 8083 23158
rect 0 22946 480 22976
rect 1577 22946 1643 22949
rect 0 22944 1643 22946
rect 0 22888 1582 22944
rect 1638 22888 1643 22944
rect 0 22886 1643 22888
rect 0 22856 480 22886
rect 1577 22883 1643 22886
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 3417 22674 3483 22677
rect 6177 22674 6243 22677
rect 7189 22674 7255 22677
rect 3417 22672 7255 22674
rect 3417 22616 3422 22672
rect 3478 22616 6182 22672
rect 6238 22616 7194 22672
rect 7250 22616 7255 22672
rect 3417 22614 7255 22616
rect 3417 22611 3483 22614
rect 6177 22611 6243 22614
rect 7189 22611 7255 22614
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 5349 22130 5415 22133
rect 10041 22130 10107 22133
rect 5349 22128 10107 22130
rect 5349 22072 5354 22128
rect 5410 22072 10046 22128
rect 10102 22072 10107 22128
rect 5349 22070 10107 22072
rect 5349 22067 5415 22070
rect 10041 22067 10107 22070
rect 14733 21994 14799 21997
rect 9446 21992 14799 21994
rect 9446 21936 14738 21992
rect 14794 21936 14799 21992
rect 9446 21934 14799 21936
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 6637 21722 6703 21725
rect 8569 21722 8635 21725
rect 6637 21720 8635 21722
rect 6637 21664 6642 21720
rect 6698 21664 8574 21720
rect 8630 21664 8635 21720
rect 6637 21662 8635 21664
rect 6637 21659 6703 21662
rect 8569 21659 8635 21662
rect 5441 21586 5507 21589
rect 7097 21586 7163 21589
rect 5441 21584 7163 21586
rect 5441 21528 5446 21584
rect 5502 21528 7102 21584
rect 7158 21528 7163 21584
rect 5441 21526 7163 21528
rect 5441 21523 5507 21526
rect 7097 21523 7163 21526
rect 5165 21450 5231 21453
rect 7465 21450 7531 21453
rect 8201 21452 8267 21453
rect 5165 21448 7531 21450
rect 5165 21392 5170 21448
rect 5226 21392 7470 21448
rect 7526 21392 7531 21448
rect 5165 21390 7531 21392
rect 5165 21387 5231 21390
rect 7465 21387 7531 21390
rect 8150 21388 8156 21452
rect 8220 21450 8267 21452
rect 8220 21448 8312 21450
rect 8262 21392 8312 21448
rect 8220 21390 8312 21392
rect 8220 21388 8267 21390
rect 8201 21387 8267 21388
rect 7741 21314 7807 21317
rect 9305 21314 9371 21317
rect 9446 21314 9506 21934
rect 14733 21931 14799 21934
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 7741 21312 9506 21314
rect 7741 21256 7746 21312
rect 7802 21256 9310 21312
rect 9366 21256 9506 21312
rect 7741 21254 9506 21256
rect 7741 21251 7807 21254
rect 9305 21251 9371 21254
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 9765 21178 9831 21181
rect 7974 21176 9831 21178
rect 7974 21120 9770 21176
rect 9826 21120 9831 21176
rect 7974 21118 9831 21120
rect 0 21042 480 21072
rect 1669 21042 1735 21045
rect 0 21040 1735 21042
rect 0 20984 1674 21040
rect 1730 20984 1735 21040
rect 0 20982 1735 20984
rect 0 20952 480 20982
rect 1669 20979 1735 20982
rect 4613 21042 4679 21045
rect 7974 21042 8034 21118
rect 9765 21115 9831 21118
rect 4613 21040 8034 21042
rect 4613 20984 4618 21040
rect 4674 20984 8034 21040
rect 4613 20982 8034 20984
rect 8109 21042 8175 21045
rect 12801 21042 12867 21045
rect 8109 21040 12867 21042
rect 8109 20984 8114 21040
rect 8170 20984 12806 21040
rect 12862 20984 12867 21040
rect 8109 20982 12867 20984
rect 4613 20979 4679 20982
rect 8109 20979 8175 20982
rect 12801 20979 12867 20982
rect 3141 20906 3207 20909
rect 3969 20906 4035 20909
rect 9857 20906 9923 20909
rect 3141 20904 9923 20906
rect 3141 20848 3146 20904
rect 3202 20848 3974 20904
rect 4030 20848 9862 20904
rect 9918 20848 9923 20904
rect 3141 20846 9923 20848
rect 3141 20843 3207 20846
rect 3969 20843 4035 20846
rect 9857 20843 9923 20846
rect 9765 20772 9831 20773
rect 9765 20770 9812 20772
rect 9720 20768 9812 20770
rect 9720 20712 9770 20768
rect 9720 20710 9812 20712
rect 9765 20708 9812 20710
rect 9876 20708 9882 20772
rect 9765 20707 9831 20708
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 9949 19954 10015 19957
rect 12433 19954 12499 19957
rect 9949 19952 12499 19954
rect 9949 19896 9954 19952
rect 10010 19896 12438 19952
rect 12494 19896 12499 19952
rect 9949 19894 12499 19896
rect 9949 19891 10015 19894
rect 12433 19891 12499 19894
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 4429 19410 4495 19413
rect 7649 19410 7715 19413
rect 4429 19408 7715 19410
rect 4429 19352 4434 19408
rect 4490 19352 7654 19408
rect 7710 19352 7715 19408
rect 4429 19350 7715 19352
rect 4429 19347 4495 19350
rect 7649 19347 7715 19350
rect 9438 19348 9444 19412
rect 9508 19410 9514 19412
rect 9581 19410 9647 19413
rect 9508 19408 9647 19410
rect 9508 19352 9586 19408
rect 9642 19352 9647 19408
rect 9508 19350 9647 19352
rect 9508 19348 9514 19350
rect 9581 19347 9647 19350
rect 7281 19274 7347 19277
rect 11789 19274 11855 19277
rect 12617 19274 12683 19277
rect 7281 19272 12683 19274
rect 7281 19216 7286 19272
rect 7342 19216 11794 19272
rect 11850 19216 12622 19272
rect 12678 19216 12683 19272
rect 7281 19214 12683 19216
rect 7281 19211 7347 19214
rect 11789 19211 11855 19214
rect 12617 19211 12683 19214
rect 7557 19138 7623 19141
rect 10869 19138 10935 19141
rect 7557 19136 10935 19138
rect 7557 19080 7562 19136
rect 7618 19080 10874 19136
rect 10930 19080 10935 19136
rect 7557 19078 10935 19080
rect 7557 19075 7623 19078
rect 10869 19075 10935 19078
rect 6277 19072 6597 19073
rect 0 19002 480 19032
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 1577 19002 1643 19005
rect 0 19000 1643 19002
rect 0 18944 1582 19000
rect 1638 18944 1643 19000
rect 0 18942 1643 18944
rect 0 18912 480 18942
rect 1577 18939 1643 18942
rect 1393 18866 1459 18869
rect 6729 18866 6795 18869
rect 1393 18864 6795 18866
rect 1393 18808 1398 18864
rect 1454 18808 6734 18864
rect 6790 18808 6795 18864
rect 1393 18806 6795 18808
rect 1393 18803 1459 18806
rect 6729 18803 6795 18806
rect 9438 18804 9444 18868
rect 9508 18866 9514 18868
rect 9581 18866 9647 18869
rect 11053 18866 11119 18869
rect 9508 18864 11119 18866
rect 9508 18808 9586 18864
rect 9642 18808 11058 18864
rect 11114 18808 11119 18864
rect 9508 18806 11119 18808
rect 9508 18804 9514 18806
rect 9581 18803 9647 18806
rect 11053 18803 11119 18806
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 8702 18260 8708 18324
rect 8772 18322 8778 18324
rect 9305 18322 9371 18325
rect 8772 18320 9371 18322
rect 8772 18264 9310 18320
rect 9366 18264 9371 18320
rect 8772 18262 9371 18264
rect 8772 18260 8778 18262
rect 9305 18259 9371 18262
rect 2221 18186 2287 18189
rect 10041 18186 10107 18189
rect 2221 18184 10107 18186
rect 2221 18128 2226 18184
rect 2282 18128 10046 18184
rect 10102 18128 10107 18184
rect 2221 18126 10107 18128
rect 2221 18123 2287 18126
rect 10041 18123 10107 18126
rect 9305 18050 9371 18053
rect 10777 18050 10843 18053
rect 9305 18048 10843 18050
rect 9305 17992 9310 18048
rect 9366 17992 10782 18048
rect 10838 17992 10843 18048
rect 9305 17990 10843 17992
rect 9305 17987 9371 17990
rect 10777 17987 10843 17990
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 9305 17914 9371 17917
rect 9581 17914 9647 17917
rect 11053 17914 11119 17917
rect 9305 17912 11119 17914
rect 9305 17856 9310 17912
rect 9366 17856 9586 17912
rect 9642 17856 11058 17912
rect 11114 17856 11119 17912
rect 9305 17854 11119 17856
rect 9305 17851 9371 17854
rect 9581 17851 9647 17854
rect 11053 17851 11119 17854
rect 5625 17642 5691 17645
rect 10593 17642 10659 17645
rect 5625 17640 10659 17642
rect 5625 17584 5630 17640
rect 5686 17584 10598 17640
rect 10654 17584 10659 17640
rect 5625 17582 10659 17584
rect 5625 17579 5691 17582
rect 10593 17579 10659 17582
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 5165 17234 5231 17237
rect 11329 17234 11395 17237
rect 12157 17234 12223 17237
rect 5165 17232 12223 17234
rect 5165 17176 5170 17232
rect 5226 17176 11334 17232
rect 11390 17176 12162 17232
rect 12218 17176 12223 17232
rect 5165 17174 12223 17176
rect 5165 17171 5231 17174
rect 11329 17171 11395 17174
rect 12157 17171 12223 17174
rect 0 16962 480 16992
rect 1577 16962 1643 16965
rect 0 16960 1643 16962
rect 0 16904 1582 16960
rect 1638 16904 1643 16960
rect 0 16902 1643 16904
rect 0 16872 480 16902
rect 1577 16899 1643 16902
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 3233 16826 3299 16829
rect 4153 16826 4219 16829
rect 3233 16824 4219 16826
rect 3233 16768 3238 16824
rect 3294 16768 4158 16824
rect 4214 16768 4219 16824
rect 3233 16766 4219 16768
rect 3233 16763 3299 16766
rect 4153 16763 4219 16766
rect 13537 16690 13603 16693
rect 15520 16690 16000 16720
rect 13537 16688 16000 16690
rect 13537 16632 13542 16688
rect 13598 16632 16000 16688
rect 13537 16630 16000 16632
rect 13537 16627 13603 16630
rect 15520 16600 16000 16630
rect 4613 16554 4679 16557
rect 10409 16554 10475 16557
rect 4613 16552 10475 16554
rect 4613 16496 4618 16552
rect 4674 16496 10414 16552
rect 10470 16496 10475 16552
rect 4613 16494 10475 16496
rect 4613 16491 4679 16494
rect 10409 16491 10475 16494
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 7649 16146 7715 16149
rect 9949 16146 10015 16149
rect 7649 16144 10015 16146
rect 7649 16088 7654 16144
rect 7710 16088 9954 16144
rect 10010 16088 10015 16144
rect 7649 16086 10015 16088
rect 7649 16083 7715 16086
rect 9949 16083 10015 16086
rect 6177 16010 6243 16013
rect 9857 16010 9923 16013
rect 6177 16008 9923 16010
rect 6177 15952 6182 16008
rect 6238 15952 9862 16008
rect 9918 15952 9923 16008
rect 6177 15950 9923 15952
rect 6177 15947 6243 15950
rect 9857 15947 9923 15950
rect 6821 15874 6887 15877
rect 8201 15874 8267 15877
rect 6821 15872 8267 15874
rect 6821 15816 6826 15872
rect 6882 15816 8206 15872
rect 8262 15816 8267 15872
rect 6821 15814 8267 15816
rect 6821 15811 6887 15814
rect 8201 15811 8267 15814
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 5901 15738 5967 15741
rect 5901 15736 6194 15738
rect 5901 15680 5906 15736
rect 5962 15680 6194 15736
rect 5901 15678 6194 15680
rect 5901 15675 5967 15678
rect 6134 15605 6194 15678
rect 2681 15602 2747 15605
rect 5901 15602 5967 15605
rect 2681 15600 5967 15602
rect 2681 15544 2686 15600
rect 2742 15544 5906 15600
rect 5962 15544 5967 15600
rect 2681 15542 5967 15544
rect 6134 15600 6243 15605
rect 6134 15544 6182 15600
rect 6238 15544 6243 15600
rect 6134 15542 6243 15544
rect 2681 15539 2747 15542
rect 5901 15539 5967 15542
rect 6177 15539 6243 15542
rect 8201 15602 8267 15605
rect 10133 15602 10199 15605
rect 10409 15602 10475 15605
rect 8201 15600 10475 15602
rect 8201 15544 8206 15600
rect 8262 15544 10138 15600
rect 10194 15544 10414 15600
rect 10470 15544 10475 15600
rect 8201 15542 10475 15544
rect 8201 15539 8267 15542
rect 10133 15539 10199 15542
rect 10409 15539 10475 15542
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 10777 15194 10843 15197
rect 11329 15194 11395 15197
rect 10777 15192 11395 15194
rect 10777 15136 10782 15192
rect 10838 15136 11334 15192
rect 11390 15136 11395 15192
rect 10777 15134 11395 15136
rect 10777 15131 10843 15134
rect 11329 15131 11395 15134
rect 7189 15058 7255 15061
rect 9857 15058 9923 15061
rect 7189 15056 9923 15058
rect 7189 15000 7194 15056
rect 7250 15000 9862 15056
rect 9918 15000 9923 15056
rect 7189 14998 9923 15000
rect 7189 14995 7255 14998
rect 9857 14995 9923 14998
rect 0 14922 480 14952
rect 1669 14922 1735 14925
rect 0 14920 1735 14922
rect 0 14864 1674 14920
rect 1730 14864 1735 14920
rect 0 14862 1735 14864
rect 0 14832 480 14862
rect 1669 14859 1735 14862
rect 2221 14922 2287 14925
rect 10041 14922 10107 14925
rect 2221 14920 10107 14922
rect 2221 14864 2226 14920
rect 2282 14864 10046 14920
rect 10102 14864 10107 14920
rect 2221 14862 10107 14864
rect 2221 14859 2287 14862
rect 10041 14859 10107 14862
rect 7189 14786 7255 14789
rect 9673 14786 9739 14789
rect 7189 14784 9739 14786
rect 7189 14728 7194 14784
rect 7250 14728 9678 14784
rect 9734 14728 9739 14784
rect 7189 14726 9739 14728
rect 7189 14723 7255 14726
rect 9673 14723 9739 14726
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 6177 14512 6243 14517
rect 6177 14456 6182 14512
rect 6238 14456 6243 14512
rect 6177 14451 6243 14456
rect 4429 14378 4495 14381
rect 6180 14378 6240 14451
rect 10133 14378 10199 14381
rect 4429 14376 10199 14378
rect 4429 14320 4434 14376
rect 4490 14320 10138 14376
rect 10194 14320 10199 14376
rect 4429 14318 10199 14320
rect 4429 14315 4495 14318
rect 10133 14315 10199 14318
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 4521 13970 4587 13973
rect 10225 13970 10291 13973
rect 4521 13968 10291 13970
rect 4521 13912 4526 13968
rect 4582 13912 10230 13968
rect 10286 13912 10291 13968
rect 4521 13910 10291 13912
rect 4521 13907 4587 13910
rect 10225 13907 10291 13910
rect 5809 13834 5875 13837
rect 7465 13834 7531 13837
rect 5809 13832 7531 13834
rect 5809 13776 5814 13832
rect 5870 13776 7470 13832
rect 7526 13776 7531 13832
rect 5809 13774 7531 13776
rect 5809 13771 5875 13774
rect 7465 13771 7531 13774
rect 8702 13772 8708 13836
rect 8772 13834 8778 13836
rect 9489 13834 9555 13837
rect 8772 13832 9555 13834
rect 8772 13776 9494 13832
rect 9550 13776 9555 13832
rect 8772 13774 9555 13776
rect 8772 13772 8778 13774
rect 9489 13771 9555 13774
rect 6729 13698 6795 13701
rect 8109 13698 8175 13701
rect 10317 13698 10383 13701
rect 6729 13696 10383 13698
rect 6729 13640 6734 13696
rect 6790 13640 8114 13696
rect 8170 13640 10322 13696
rect 10378 13640 10383 13696
rect 6729 13638 10383 13640
rect 6729 13635 6795 13638
rect 8109 13635 8175 13638
rect 10317 13635 10383 13638
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 4245 13426 4311 13429
rect 10317 13426 10383 13429
rect 4245 13424 10383 13426
rect 4245 13368 4250 13424
rect 4306 13368 10322 13424
rect 10378 13368 10383 13424
rect 4245 13366 10383 13368
rect 4245 13363 4311 13366
rect 10317 13363 10383 13366
rect 10869 13426 10935 13429
rect 12157 13426 12223 13429
rect 10869 13424 12223 13426
rect 10869 13368 10874 13424
rect 10930 13368 12162 13424
rect 12218 13368 12223 13424
rect 10869 13366 12223 13368
rect 10869 13363 10935 13366
rect 12157 13363 12223 13366
rect 12709 13290 12775 13293
rect 9584 13288 12775 13290
rect 9584 13232 12714 13288
rect 12770 13232 12775 13288
rect 9584 13230 12775 13232
rect 3610 13088 3930 13089
rect 0 13018 480 13048
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 1577 13018 1643 13021
rect 0 13016 1643 13018
rect 0 12960 1582 13016
rect 1638 12960 1643 13016
rect 0 12958 1643 12960
rect 0 12928 480 12958
rect 1577 12955 1643 12958
rect 8017 12882 8083 12885
rect 9584 12882 9644 13230
rect 12709 13227 12775 13230
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 8017 12880 9644 12882
rect 8017 12824 8022 12880
rect 8078 12824 9644 12880
rect 8017 12822 9644 12824
rect 8017 12819 8083 12822
rect 1669 12610 1735 12613
rect 5533 12610 5599 12613
rect 1669 12608 5599 12610
rect 1669 12552 1674 12608
rect 1730 12552 5538 12608
rect 5594 12552 5599 12608
rect 1669 12550 5599 12552
rect 1669 12547 1735 12550
rect 5533 12547 5599 12550
rect 6729 12610 6795 12613
rect 8845 12610 8911 12613
rect 6729 12608 8911 12610
rect 6729 12552 6734 12608
rect 6790 12552 8850 12608
rect 8906 12552 8911 12608
rect 6729 12550 8911 12552
rect 6729 12547 6795 12550
rect 8845 12547 8911 12550
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 4889 12474 4955 12477
rect 4846 12472 4955 12474
rect 4846 12416 4894 12472
rect 4950 12416 4955 12472
rect 4846 12411 4955 12416
rect 11053 12474 11119 12477
rect 11329 12474 11395 12477
rect 11053 12472 11395 12474
rect 11053 12416 11058 12472
rect 11114 12416 11334 12472
rect 11390 12416 11395 12472
rect 11053 12414 11395 12416
rect 11053 12411 11119 12414
rect 11329 12411 11395 12414
rect 4846 12341 4906 12411
rect 4846 12336 4955 12341
rect 4846 12280 4894 12336
rect 4950 12280 4955 12336
rect 4846 12278 4955 12280
rect 4889 12275 4955 12278
rect 8845 12338 8911 12341
rect 10777 12338 10843 12341
rect 11329 12338 11395 12341
rect 8845 12336 11395 12338
rect 8845 12280 8850 12336
rect 8906 12280 10782 12336
rect 10838 12280 11334 12336
rect 11390 12280 11395 12336
rect 8845 12278 11395 12280
rect 8845 12275 8911 12278
rect 10777 12275 10843 12278
rect 11329 12275 11395 12278
rect 5809 12202 5875 12205
rect 10685 12202 10751 12205
rect 5809 12200 10751 12202
rect 5809 12144 5814 12200
rect 5870 12144 10690 12200
rect 10746 12144 10751 12200
rect 5809 12142 10751 12144
rect 5809 12139 5875 12142
rect 10685 12139 10751 12142
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 8017 11794 8083 11797
rect 10041 11794 10107 11797
rect 8017 11792 10107 11794
rect 8017 11736 8022 11792
rect 8078 11736 10046 11792
rect 10102 11736 10107 11792
rect 8017 11734 10107 11736
rect 8017 11731 8083 11734
rect 10041 11731 10107 11734
rect 8477 11658 8543 11661
rect 11421 11658 11487 11661
rect 8477 11656 11487 11658
rect 8477 11600 8482 11656
rect 8538 11600 11426 11656
rect 11482 11600 11487 11656
rect 8477 11598 11487 11600
rect 8477 11595 8543 11598
rect 11421 11595 11487 11598
rect 2221 11522 2287 11525
rect 4797 11522 4863 11525
rect 2221 11520 4863 11522
rect 2221 11464 2226 11520
rect 2282 11464 4802 11520
rect 4858 11464 4863 11520
rect 2221 11462 4863 11464
rect 2221 11459 2287 11462
rect 4797 11459 4863 11462
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 5993 11114 6059 11117
rect 8201 11114 8267 11117
rect 5993 11112 8267 11114
rect 5993 11056 5998 11112
rect 6054 11056 8206 11112
rect 8262 11056 8267 11112
rect 5993 11054 8267 11056
rect 5993 11051 6059 11054
rect 8201 11051 8267 11054
rect 0 10978 480 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 480 10918
rect 1577 10915 1643 10918
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 9397 10842 9463 10845
rect 11881 10842 11947 10845
rect 9397 10840 11947 10842
rect 9397 10784 9402 10840
rect 9458 10784 11886 10840
rect 11942 10784 11947 10840
rect 9397 10782 11947 10784
rect 9397 10779 9463 10782
rect 11881 10779 11947 10782
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 8477 10298 8543 10301
rect 9397 10298 9463 10301
rect 8477 10296 9463 10298
rect 8477 10240 8482 10296
rect 8538 10240 9402 10296
rect 9458 10240 9463 10296
rect 8477 10238 9463 10240
rect 8477 10235 8543 10238
rect 9397 10235 9463 10238
rect 8937 10162 9003 10165
rect 9438 10162 9444 10164
rect 8937 10160 9444 10162
rect 8937 10104 8942 10160
rect 8998 10104 9444 10160
rect 8937 10102 9444 10104
rect 8937 10099 9003 10102
rect 9438 10100 9444 10102
rect 9508 10162 9514 10164
rect 15377 10162 15443 10165
rect 9508 10160 15443 10162
rect 9508 10104 15382 10160
rect 15438 10104 15443 10160
rect 9508 10102 15443 10104
rect 9508 10100 9514 10102
rect 15377 10099 15443 10102
rect 13905 10026 13971 10029
rect 15520 10026 16000 10056
rect 13905 10024 16000 10026
rect 13905 9968 13910 10024
rect 13966 9968 16000 10024
rect 13905 9966 16000 9968
rect 13905 9963 13971 9966
rect 15520 9936 16000 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 4705 9754 4771 9757
rect 6913 9754 6979 9757
rect 4705 9752 6979 9754
rect 4705 9696 4710 9752
rect 4766 9696 6918 9752
rect 6974 9696 6979 9752
rect 4705 9694 6979 9696
rect 4705 9691 4771 9694
rect 6913 9691 6979 9694
rect 2037 9618 2103 9621
rect 3877 9618 3943 9621
rect 2037 9616 3943 9618
rect 2037 9560 2042 9616
rect 2098 9560 3882 9616
rect 3938 9560 3943 9616
rect 2037 9558 3943 9560
rect 2037 9555 2103 9558
rect 3877 9555 3943 9558
rect 9305 9618 9371 9621
rect 10869 9618 10935 9621
rect 9305 9616 10935 9618
rect 9305 9560 9310 9616
rect 9366 9560 10874 9616
rect 10930 9560 10935 9616
rect 9305 9558 10935 9560
rect 9305 9555 9371 9558
rect 10869 9555 10935 9558
rect 5809 9482 5875 9485
rect 9121 9482 9187 9485
rect 5809 9480 9187 9482
rect 5809 9424 5814 9480
rect 5870 9424 9126 9480
rect 9182 9424 9187 9480
rect 5809 9422 9187 9424
rect 5809 9419 5875 9422
rect 9121 9419 9187 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 8109 9074 8175 9077
rect 9765 9074 9831 9077
rect 8109 9072 9831 9074
rect 8109 9016 8114 9072
rect 8170 9016 9770 9072
rect 9826 9016 9831 9072
rect 8109 9014 9831 9016
rect 8109 9011 8175 9014
rect 9765 9011 9831 9014
rect 0 8938 480 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 480 8878
rect 1577 8875 1643 8878
rect 5349 8938 5415 8941
rect 14181 8938 14247 8941
rect 5349 8936 14247 8938
rect 5349 8880 5354 8936
rect 5410 8880 14186 8936
rect 14242 8880 14247 8936
rect 5349 8878 14247 8880
rect 5349 8875 5415 8878
rect 14181 8875 14247 8878
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 7557 8666 7623 8669
rect 8569 8666 8635 8669
rect 7557 8664 8635 8666
rect 7557 8608 7562 8664
rect 7618 8608 8574 8664
rect 8630 8608 8635 8664
rect 7557 8606 8635 8608
rect 7557 8603 7623 8606
rect 8569 8603 8635 8606
rect 3785 8394 3851 8397
rect 3969 8394 4035 8397
rect 5809 8394 5875 8397
rect 3785 8392 5875 8394
rect 3785 8336 3790 8392
rect 3846 8336 3974 8392
rect 4030 8336 5814 8392
rect 5870 8336 5875 8392
rect 3785 8334 5875 8336
rect 3785 8331 3851 8334
rect 3969 8331 4035 8334
rect 5809 8331 5875 8334
rect 8201 8258 8267 8261
rect 10225 8258 10291 8261
rect 8201 8256 10291 8258
rect 8201 8200 8206 8256
rect 8262 8200 10230 8256
rect 10286 8200 10291 8256
rect 8201 8198 10291 8200
rect 8201 8195 8267 8198
rect 10225 8195 10291 8198
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 4981 7986 5047 7989
rect 8385 7986 8451 7989
rect 4981 7984 8451 7986
rect 4981 7928 4986 7984
rect 5042 7928 8390 7984
rect 8446 7928 8451 7984
rect 4981 7926 8451 7928
rect 4981 7923 5047 7926
rect 8385 7923 8451 7926
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 2497 7442 2563 7445
rect 4981 7442 5047 7445
rect 2497 7440 5047 7442
rect 2497 7384 2502 7440
rect 2558 7384 4986 7440
rect 5042 7384 5047 7440
rect 2497 7382 5047 7384
rect 2497 7379 2563 7382
rect 4981 7379 5047 7382
rect 8937 7442 9003 7445
rect 12801 7442 12867 7445
rect 8937 7440 12867 7442
rect 8937 7384 8942 7440
rect 8998 7384 12806 7440
rect 12862 7384 12867 7440
rect 8937 7382 12867 7384
rect 8937 7379 9003 7382
rect 12801 7379 12867 7382
rect 4061 7306 4127 7309
rect 9673 7306 9739 7309
rect 4061 7304 9739 7306
rect 4061 7248 4066 7304
rect 4122 7248 9678 7304
rect 9734 7248 9739 7304
rect 4061 7246 9739 7248
rect 4061 7243 4127 7246
rect 9673 7243 9739 7246
rect 8109 7170 8175 7173
rect 10133 7170 10199 7173
rect 8109 7168 10199 7170
rect 8109 7112 8114 7168
rect 8170 7112 10138 7168
rect 10194 7112 10199 7168
rect 8109 7110 10199 7112
rect 8109 7107 8175 7110
rect 10133 7107 10199 7110
rect 6277 7104 6597 7105
rect 0 7034 480 7064
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 2313 7034 2379 7037
rect 0 7032 2379 7034
rect 0 6976 2318 7032
rect 2374 6976 2379 7032
rect 0 6974 2379 6976
rect 0 6944 480 6974
rect 2313 6971 2379 6974
rect 6177 6898 6243 6901
rect 7925 6898 7991 6901
rect 6177 6896 7991 6898
rect 6177 6840 6182 6896
rect 6238 6840 7930 6896
rect 7986 6840 7991 6896
rect 6177 6838 7991 6840
rect 6177 6835 6243 6838
rect 7925 6835 7991 6838
rect 9213 6898 9279 6901
rect 9397 6898 9463 6901
rect 9213 6896 9463 6898
rect 9213 6840 9218 6896
rect 9274 6840 9402 6896
rect 9458 6840 9463 6896
rect 9213 6838 9463 6840
rect 9213 6835 9279 6838
rect 9397 6835 9463 6838
rect 5533 6626 5599 6629
rect 8569 6626 8635 6629
rect 5533 6624 8635 6626
rect 5533 6568 5538 6624
rect 5594 6568 8574 6624
rect 8630 6568 8635 6624
rect 5533 6566 8635 6568
rect 5533 6563 5599 6566
rect 8569 6563 8635 6566
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 6637 6490 6703 6493
rect 8201 6490 8267 6493
rect 6637 6488 8267 6490
rect 6637 6432 6642 6488
rect 6698 6432 8206 6488
rect 8262 6432 8267 6488
rect 6637 6430 8267 6432
rect 6637 6427 6703 6430
rect 8201 6427 8267 6430
rect 6637 6354 6703 6357
rect 12433 6354 12499 6357
rect 6637 6352 12499 6354
rect 6637 6296 6642 6352
rect 6698 6296 12438 6352
rect 12494 6296 12499 6352
rect 6637 6294 12499 6296
rect 6637 6291 6703 6294
rect 12433 6291 12499 6294
rect 4429 6218 4495 6221
rect 5073 6218 5139 6221
rect 8017 6218 8083 6221
rect 12249 6218 12315 6221
rect 4429 6216 7666 6218
rect 4429 6160 4434 6216
rect 4490 6160 5078 6216
rect 5134 6160 7666 6216
rect 4429 6158 7666 6160
rect 4429 6155 4495 6158
rect 5073 6155 5139 6158
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 1485 5810 1551 5813
rect 7465 5810 7531 5813
rect 1485 5808 7531 5810
rect 1485 5752 1490 5808
rect 1546 5752 7470 5808
rect 7526 5752 7531 5808
rect 1485 5750 7531 5752
rect 1485 5747 1551 5750
rect 7465 5747 7531 5750
rect 5257 5674 5323 5677
rect 6729 5674 6795 5677
rect 5257 5672 6795 5674
rect 5257 5616 5262 5672
rect 5318 5616 6734 5672
rect 6790 5616 6795 5672
rect 5257 5614 6795 5616
rect 7606 5674 7666 6158
rect 8017 6216 12315 6218
rect 8017 6160 8022 6216
rect 8078 6160 12254 6216
rect 12310 6160 12315 6216
rect 8017 6158 12315 6160
rect 8017 6155 8083 6158
rect 12249 6155 12315 6158
rect 9489 6084 9555 6085
rect 9438 6020 9444 6084
rect 9508 6082 9555 6084
rect 9508 6080 9600 6082
rect 9550 6024 9600 6080
rect 9508 6022 9600 6024
rect 9508 6020 9555 6022
rect 9489 6019 9555 6020
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 7741 5810 7807 5813
rect 11053 5810 11119 5813
rect 7741 5808 11119 5810
rect 7741 5752 7746 5808
rect 7802 5752 11058 5808
rect 11114 5752 11119 5808
rect 7741 5750 11119 5752
rect 7741 5747 7807 5750
rect 11053 5747 11119 5750
rect 12525 5674 12591 5677
rect 13445 5674 13511 5677
rect 7606 5672 13511 5674
rect 7606 5616 12530 5672
rect 12586 5616 13450 5672
rect 13506 5616 13511 5672
rect 7606 5614 13511 5616
rect 5257 5611 5323 5614
rect 6729 5611 6795 5614
rect 12525 5611 12591 5614
rect 13445 5611 13511 5614
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 3049 5266 3115 5269
rect 4521 5266 4587 5269
rect 9765 5266 9831 5269
rect 3049 5264 9831 5266
rect 3049 5208 3054 5264
rect 3110 5208 4526 5264
rect 4582 5208 9770 5264
rect 9826 5208 9831 5264
rect 3049 5206 9831 5208
rect 3049 5203 3115 5206
rect 4521 5203 4587 5206
rect 9765 5203 9831 5206
rect 5809 5130 5875 5133
rect 9305 5130 9371 5133
rect 11605 5130 11671 5133
rect 5809 5128 6010 5130
rect 5809 5072 5814 5128
rect 5870 5072 6010 5128
rect 5809 5070 6010 5072
rect 5809 5067 5875 5070
rect 0 4994 480 5024
rect 1577 4994 1643 4997
rect 0 4992 1643 4994
rect 0 4936 1582 4992
rect 1638 4936 1643 4992
rect 0 4934 1643 4936
rect 0 4904 480 4934
rect 1577 4931 1643 4934
rect 5950 4722 6010 5070
rect 9305 5128 11671 5130
rect 9305 5072 9310 5128
rect 9366 5072 11610 5128
rect 11666 5072 11671 5128
rect 9305 5070 11671 5072
rect 9305 5067 9371 5070
rect 11605 5067 11671 5070
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 10777 4858 10843 4861
rect 6686 4856 10843 4858
rect 6686 4800 10782 4856
rect 10838 4800 10843 4856
rect 6686 4798 10843 4800
rect 6686 4722 6746 4798
rect 10777 4795 10843 4798
rect 5950 4662 6746 4722
rect 7465 4722 7531 4725
rect 9857 4722 9923 4725
rect 7465 4720 9923 4722
rect 7465 4664 7470 4720
rect 7526 4664 9862 4720
rect 9918 4664 9923 4720
rect 7465 4662 9923 4664
rect 7465 4659 7531 4662
rect 9857 4659 9923 4662
rect 3877 4586 3943 4589
rect 5073 4586 5139 4589
rect 3877 4584 5139 4586
rect 3877 4528 3882 4584
rect 3938 4528 5078 4584
rect 5134 4528 5139 4584
rect 3877 4526 5139 4528
rect 3877 4523 3943 4526
rect 5073 4523 5139 4526
rect 6821 4586 6887 4589
rect 8477 4586 8543 4589
rect 6821 4584 8543 4586
rect 6821 4528 6826 4584
rect 6882 4528 8482 4584
rect 8538 4528 8543 4584
rect 6821 4526 8543 4528
rect 6821 4523 6887 4526
rect 8477 4523 8543 4526
rect 4153 4450 4219 4453
rect 7005 4450 7071 4453
rect 4153 4448 7071 4450
rect 4153 4392 4158 4448
rect 4214 4392 7010 4448
rect 7066 4392 7071 4448
rect 4153 4390 7071 4392
rect 4153 4387 4219 4390
rect 7005 4387 7071 4390
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 7005 4178 7071 4181
rect 11053 4178 11119 4181
rect 7005 4176 11119 4178
rect 7005 4120 7010 4176
rect 7066 4120 11058 4176
rect 11114 4120 11119 4176
rect 7005 4118 11119 4120
rect 7005 4115 7071 4118
rect 11053 4115 11119 4118
rect 4337 4042 4403 4045
rect 4797 4042 4863 4045
rect 4337 4040 4863 4042
rect 4337 3984 4342 4040
rect 4398 3984 4802 4040
rect 4858 3984 4863 4040
rect 4337 3982 4863 3984
rect 4337 3979 4403 3982
rect 4797 3979 4863 3982
rect 6177 4042 6243 4045
rect 8385 4042 8451 4045
rect 6177 4040 8451 4042
rect 6177 3984 6182 4040
rect 6238 3984 8390 4040
rect 8446 3984 8451 4040
rect 6177 3982 8451 3984
rect 6177 3979 6243 3982
rect 8385 3979 8451 3982
rect 8753 4042 8819 4045
rect 13353 4042 13419 4045
rect 8753 4040 13419 4042
rect 8753 3984 8758 4040
rect 8814 3984 13358 4040
rect 13414 3984 13419 4040
rect 8753 3982 13419 3984
rect 8753 3979 8819 3982
rect 13353 3979 13419 3982
rect 8017 3906 8083 3909
rect 10685 3906 10751 3909
rect 11329 3906 11395 3909
rect 8017 3904 11395 3906
rect 8017 3848 8022 3904
rect 8078 3848 10690 3904
rect 10746 3848 11334 3904
rect 11390 3848 11395 3904
rect 8017 3846 11395 3848
rect 8017 3843 8083 3846
rect 10685 3843 10751 3846
rect 11329 3843 11395 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 7189 3770 7255 3773
rect 8753 3770 8819 3773
rect 9673 3770 9739 3773
rect 7189 3768 9739 3770
rect 7189 3712 7194 3768
rect 7250 3712 8758 3768
rect 8814 3712 9678 3768
rect 9734 3712 9739 3768
rect 7189 3710 9739 3712
rect 7189 3707 7255 3710
rect 8753 3707 8819 3710
rect 9673 3707 9739 3710
rect 7833 3634 7899 3637
rect 10685 3634 10751 3637
rect 12617 3634 12683 3637
rect 7833 3632 10610 3634
rect 7833 3576 7838 3632
rect 7894 3576 10610 3632
rect 7833 3574 10610 3576
rect 7833 3571 7899 3574
rect 10550 3501 10610 3574
rect 10685 3632 12683 3634
rect 10685 3576 10690 3632
rect 10746 3576 12622 3632
rect 12678 3576 12683 3632
rect 10685 3574 12683 3576
rect 10685 3571 10751 3574
rect 12617 3571 12683 3574
rect 10225 3498 10291 3501
rect 8710 3496 10291 3498
rect 8710 3440 10230 3496
rect 10286 3440 10291 3496
rect 8710 3438 10291 3440
rect 10550 3496 10659 3501
rect 10550 3440 10598 3496
rect 10654 3440 10659 3496
rect 10550 3438 10659 3440
rect 6821 3362 6887 3365
rect 8710 3362 8770 3438
rect 10225 3435 10291 3438
rect 10593 3435 10659 3438
rect 12065 3498 12131 3501
rect 12065 3496 14842 3498
rect 12065 3440 12070 3496
rect 12126 3440 14842 3496
rect 12065 3438 14842 3440
rect 12065 3435 12131 3438
rect 6821 3360 8770 3362
rect 6821 3304 6826 3360
rect 6882 3304 8770 3360
rect 6821 3302 8770 3304
rect 14782 3362 14842 3438
rect 15520 3362 16000 3392
rect 14782 3302 16000 3362
rect 6821 3299 6887 3302
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 15520 3272 16000 3302
rect 14277 3231 14597 3232
rect 933 3090 999 3093
rect 6913 3090 6979 3093
rect 933 3088 6979 3090
rect 933 3032 938 3088
rect 994 3032 6918 3088
rect 6974 3032 6979 3088
rect 933 3030 6979 3032
rect 933 3027 999 3030
rect 6913 3027 6979 3030
rect 8477 3090 8543 3093
rect 14917 3090 14983 3093
rect 8477 3088 14983 3090
rect 8477 3032 8482 3088
rect 8538 3032 14922 3088
rect 14978 3032 14983 3088
rect 8477 3030 14983 3032
rect 8477 3027 8543 3030
rect 14917 3027 14983 3030
rect 0 2954 480 2984
rect 2221 2954 2287 2957
rect 13721 2954 13787 2957
rect 0 2952 2287 2954
rect 0 2896 2226 2952
rect 2282 2896 2287 2952
rect 0 2894 2287 2896
rect 0 2864 480 2894
rect 2221 2891 2287 2894
rect 6134 2952 13787 2954
rect 6134 2896 13726 2952
rect 13782 2896 13787 2952
rect 6134 2894 13787 2896
rect 2589 2818 2655 2821
rect 4245 2818 4311 2821
rect 2589 2816 4311 2818
rect 2589 2760 2594 2816
rect 2650 2760 4250 2816
rect 4306 2760 4311 2816
rect 2589 2758 4311 2760
rect 2589 2755 2655 2758
rect 4245 2755 4311 2758
rect 4613 2818 4679 2821
rect 4797 2818 4863 2821
rect 6134 2818 6194 2894
rect 13721 2891 13787 2894
rect 9489 2820 9555 2821
rect 9438 2818 9444 2820
rect 4613 2816 6194 2818
rect 4613 2760 4618 2816
rect 4674 2760 4802 2816
rect 4858 2760 6194 2816
rect 4613 2758 6194 2760
rect 9398 2758 9444 2818
rect 9508 2816 9555 2820
rect 9550 2760 9555 2816
rect 4613 2755 4679 2758
rect 4797 2755 4863 2758
rect 9438 2756 9444 2758
rect 9508 2756 9555 2760
rect 9489 2755 9555 2756
rect 12525 2818 12591 2821
rect 12893 2818 12959 2821
rect 12525 2816 12959 2818
rect 12525 2760 12530 2816
rect 12586 2760 12898 2816
rect 12954 2760 12959 2816
rect 12525 2758 12959 2760
rect 12525 2755 12591 2758
rect 12893 2755 12959 2758
rect 13077 2818 13143 2821
rect 14641 2818 14707 2821
rect 13077 2816 14707 2818
rect 13077 2760 13082 2816
rect 13138 2760 14646 2816
rect 14702 2760 14707 2816
rect 13077 2758 14707 2760
rect 13077 2755 13143 2758
rect 14641 2755 14707 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 2405 2682 2471 2685
rect 4705 2682 4771 2685
rect 2405 2680 4771 2682
rect 2405 2624 2410 2680
rect 2466 2624 4710 2680
rect 4766 2624 4771 2680
rect 2405 2622 4771 2624
rect 2405 2619 2471 2622
rect 4705 2619 4771 2622
rect 3877 2546 3943 2549
rect 7465 2546 7531 2549
rect 3877 2544 7531 2546
rect 3877 2488 3882 2544
rect 3938 2488 7470 2544
rect 7526 2488 7531 2544
rect 3877 2486 7531 2488
rect 3877 2483 3943 2486
rect 7465 2483 7531 2486
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 2129 1458 2195 1461
rect 7097 1458 7163 1461
rect 2129 1456 7163 1458
rect 2129 1400 2134 1456
rect 2190 1400 7102 1456
rect 7158 1400 7163 1456
rect 2129 1398 7163 1400
rect 2129 1395 2195 1398
rect 7097 1395 7163 1398
rect 0 1050 480 1080
rect 2497 1050 2563 1053
rect 0 1048 2563 1050
rect 0 992 2502 1048
rect 2558 992 2563 1048
rect 0 990 2563 992
rect 0 960 480 990
rect 2497 987 2563 990
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 8156 28732 8220 28796
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 9812 26964 9876 27028
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 9444 24380 9508 24444
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 8156 21448 8220 21452
rect 8156 21392 8206 21448
rect 8206 21392 8220 21448
rect 8156 21388 8220 21392
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 9812 20768 9876 20772
rect 9812 20712 9826 20768
rect 9826 20712 9876 20768
rect 9812 20708 9876 20712
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 9444 19348 9508 19412
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 9444 18804 9508 18868
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 8708 18260 8772 18324
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 8708 13772 8772 13836
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 9444 10100 9508 10164
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 9444 6080 9508 6084
rect 9444 6024 9494 6080
rect 9494 6024 9508 6080
rect 9444 6020 9508 6024
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 9444 2816 9508 2820
rect 9444 2760 9494 2816
rect 9494 2760 9508 2816
rect 9444 2756 9508 2760
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8155 28796 8221 28797
rect 8155 28732 8156 28796
rect 8220 28732 8221 28796
rect 8155 28731 8221 28732
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 8158 21453 8218 28731
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 9811 27028 9877 27029
rect 9811 26964 9812 27028
rect 9876 26964 9877 27028
rect 9811 26963 9877 26964
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 9443 24444 9509 24445
rect 9443 24380 9444 24444
rect 9508 24380 9509 24444
rect 9443 24379 9509 24380
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8155 21452 8221 21453
rect 8155 21388 8156 21452
rect 8220 21388 8221 21452
rect 8155 21387 8221 21388
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 9446 19413 9506 24379
rect 9814 20773 9874 26963
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 9811 20772 9877 20773
rect 9811 20708 9812 20772
rect 9876 20708 9877 20772
rect 9811 20707 9877 20708
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 9443 19412 9509 19413
rect 9443 19348 9444 19412
rect 9508 19348 9509 19412
rect 9443 19347 9509 19348
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 9443 18868 9509 18869
rect 9443 18804 9444 18868
rect 9508 18804 9509 18868
rect 9443 18803 9509 18804
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8707 18324 8773 18325
rect 8707 18260 8708 18324
rect 8772 18260 8773 18324
rect 8707 18259 8773 18260
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 8710 13837 8770 18259
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8707 13836 8773 13837
rect 8707 13772 8708 13836
rect 8772 13772 8773 13836
rect 8707 13771 8773 13772
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 9446 10165 9506 18803
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 9443 10164 9509 10165
rect 9443 10100 9444 10164
rect 9508 10100 9509 10164
rect 9443 10099 9509 10100
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 9443 6084 9509 6085
rect 9443 6020 9444 6084
rect 9508 6020 9509 6084
rect 9443 6019 9509 6020
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 9446 2821 9506 6019
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 9443 2820 9509 2821
rect 9443 2756 9444 2820
rect 9508 2756 9509 2820
rect 9443 2755 9509 2756
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_6
timestamp 1604681595
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _46_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _23_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_34 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4232 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36
timestamp 1604681595
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1604681595
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4784 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4876 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1604681595
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_50
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1604681595
transform 1 0 5980 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1604681595
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6256 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1604681595
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_66
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67
timestamp 1604681595
transform 1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7544 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_90
timestamp 1604681595
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98
timestamp 1604681595
transform 1 0 10120 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9936 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9752 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1604681595
transform 1 0 11500 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1604681595
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_142
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_136 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_36
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_40
timestamp 1604681595
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 6716 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_53
timestamp 1604681595
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_57
timestamp 1604681595
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65
timestamp 1604681595
transform 1 0 7084 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_71
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9844 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_104
timestamp 1604681595
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11408 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_108
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_128
timestamp 1604681595
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_132 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13248 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2944 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_13
timestamp 1604681595
transform 1 0 2300 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_16
timestamp 1604681595
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1604681595
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_40
timestamp 1604681595
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9936 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_88
timestamp 1604681595
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1604681595
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1604681595
transform 1 0 11500 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1604681595
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_105
timestamp 1604681595
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_136
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_144
timestamp 1604681595
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_10
timestamp 1604681595
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4600 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_54
timestamp 1604681595
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_58
timestamp 1604681595
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_78
timestamp 1604681595
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1604681595
transform 1 0 8648 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9936 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_98
timestamp 1604681595
transform 1 0 10120 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11776 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1604681595
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_136
timestamp 1604681595
transform 1 0 13616 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1604681595
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1604681595
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3404 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_21
timestamp 1604681595
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_41
timestamp 1604681595
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_45
timestamp 1604681595
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1604681595
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1604681595
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1604681595
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_106
timestamp 1604681595
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_126
timestamp 1604681595
transform 1 0 12696 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_138
timestamp 1604681595
transform 1 0 13800 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 2024 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_14
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_18
timestamp 1604681595
transform 1 0 2760 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_34
timestamp 1604681595
transform 1 0 4232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4508 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4692 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_41
timestamp 1604681595
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_45
timestamp 1604681595
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_48
timestamp 1604681595
transform 1 0 5520 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 5612 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1604681595
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_61
timestamp 1604681595
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 6348 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_67
timestamp 1604681595
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1604681595
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 6900 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1604681595
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_78
timestamp 1604681595
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_86
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_84
timestamp 1604681595
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_88
timestamp 1604681595
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9568 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1604681595
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1604681595
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_105
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_110
timestamp 1604681595
transform 1 0 11224 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1604681595
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 11132 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1604681595
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_120
timestamp 1604681595
transform 1 0 12144 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_132
timestamp 1604681595
transform 1 0 13248 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1604681595
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_143
timestamp 1604681595
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_12
timestamp 1604681595
transform 1 0 2208 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_19
timestamp 1604681595
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_40
timestamp 1604681595
transform 1 0 4784 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 5060 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 6164 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_47
timestamp 1604681595
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1604681595
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_59
timestamp 1604681595
transform 1 0 6532 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_71
timestamp 1604681595
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1604681595
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_101
timestamp 1604681595
transform 1 0 10396 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 11040 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp 1604681595
transform 1 0 10948 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_124
timestamp 1604681595
transform 1 0 12512 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_136
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1604681595
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_11
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_16
timestamp 1604681595
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_20
timestamp 1604681595
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_24
timestamp 1604681595
transform 1 0 3312 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_32
timestamp 1604681595
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_43
timestamp 1604681595
transform 1 0 5060 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_48
timestamp 1604681595
transform 1 0 5520 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 5612 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7820 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp 1604681595
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_82
timestamp 1604681595
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9384 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_99
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_103
timestamp 1604681595
transform 1 0 10580 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1604681595
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1604681595
transform 1 0 11500 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1604681595
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_143
timestamp 1604681595
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 4324 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_38
timestamp 1604681595
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 5336 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_42
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_62
timestamp 1604681595
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_70
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_104
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1604681595
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1604681595
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_143
timestamp 1604681595
transform 1 0 14260 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2668 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_9
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_13
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_16
timestamp 1604681595
transform 1 0 2576 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4232 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1604681595
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1604681595
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1604681595
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_78
timestamp 1604681595
transform 1 0 8280 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_83
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9108 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_103
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_115
timestamp 1604681595
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_9
timestamp 1604681595
transform 1 0 1932 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5612 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1604681595
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1604681595
transform 1 0 6440 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_64
timestamp 1604681595
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1604681595
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_102
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_114
timestamp 1604681595
transform 1 0 11592 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_126
timestamp 1604681595
transform 1 0 12696 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_9
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_14
timestamp 1604681595
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2760 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_38
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1604681595
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_46
timestamp 1604681595
transform 1 0 5336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_59
timestamp 1604681595
transform 1 0 6532 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_55
timestamp 1604681595
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_55
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 5888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_67
timestamp 1604681595
transform 1 0 7268 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7728 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7084 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_78
timestamp 1604681595
transform 1 0 8280 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_74
timestamp 1604681595
transform 1 0 7912 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_83
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_87
timestamp 1604681595
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1604681595
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604681595
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1604681595
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_102
timestamp 1604681595
transform 1 0 10488 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1604681595
transform 1 0 9936 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10304 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1604681595
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_107
timestamp 1604681595
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1604681595
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_122
timestamp 1604681595
transform 1 0 12328 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_116
timestamp 1604681595
transform 1 0 11776 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1604681595
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_143
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_20
timestamp 1604681595
transform 1 0 2944 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_28
timestamp 1604681595
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1604681595
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1604681595
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8556 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_73
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_77
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1604681595
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_94
timestamp 1604681595
transform 1 0 9752 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_101
timestamp 1604681595
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_144
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_9
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_13
timestamp 1604681595
transform 1 0 2300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4784 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_25
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6348 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_49
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_53
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_66
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_70
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604681595
transform 1 0 12328 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_114
timestamp 1604681595
transform 1 0 11592 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_125
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_137
timestamp 1604681595
transform 1 0 13708 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_9
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_13
timestamp 1604681595
transform 1 0 2300 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_25
timestamp 1604681595
transform 1 0 3404 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_33
timestamp 1604681595
transform 1 0 4140 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1604681595
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1604681595
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1604681595
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6900 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8464 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_72
timestamp 1604681595
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp 1604681595
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1604681595
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_143
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_17
timestamp 1604681595
transform 1 0 2668 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1604681595
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_48
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_54
timestamp 1604681595
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_67
timestamp 1604681595
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_71
timestamp 1604681595
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_96
timestamp 1604681595
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_100
timestamp 1604681595
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 11040 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_107
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_124
timestamp 1604681595
transform 1 0 12512 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_136
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1604681595
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_9
timestamp 1604681595
transform 1 0 1932 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_31
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_40
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_19_47
timestamp 1604681595
transform 1 0 5428 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1604681595
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp 1604681595
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_57
timestamp 1604681595
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 7084 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1604681595
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_82
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_81
timestamp 1604681595
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_102
timestamp 1604681595
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1604681595
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_106
timestamp 1604681595
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1604681595
transform 1 0 11132 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1604681595
transform 1 0 12236 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_133
timestamp 1604681595
transform 1 0 13340 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2300 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3864 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_22
timestamp 1604681595
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_26
timestamp 1604681595
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_46
timestamp 1604681595
transform 1 0 5336 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_55
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8464 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_66
timestamp 1604681595
transform 1 0 7176 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_76
timestamp 1604681595
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_89
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1604681595
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_143
timestamp 1604681595
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2300 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1604681595
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3128 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_21
timestamp 1604681595
transform 1 0 3036 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1604681595
transform 1 0 3312 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_28
timestamp 1604681595
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5612 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_45
timestamp 1604681595
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_58
timestamp 1604681595
transform 1 0 6440 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_64
timestamp 1604681595
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_72
timestamp 1604681595
transform 1 0 7728 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_75
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_79
timestamp 1604681595
transform 1 0 8372 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1604681595
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_86
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1604681595
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11500 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_106
timestamp 1604681595
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_110
timestamp 1604681595
transform 1 0 11224 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_9
timestamp 1604681595
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_13
timestamp 1604681595
transform 1 0 2300 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_19
timestamp 1604681595
transform 1 0 2852 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_31
timestamp 1604681595
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_35
timestamp 1604681595
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_75
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_79
timestamp 1604681595
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1604681595
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_95
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11868 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_111
timestamp 1604681595
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1604681595
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_119
timestamp 1604681595
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_131
timestamp 1604681595
transform 1 0 13156 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_142
timestamp 1604681595
transform 1 0 14168 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_21
timestamp 1604681595
transform 1 0 3036 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_24
timestamp 1604681595
transform 1 0 3312 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1604681595
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1604681595
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_58
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp 1604681595
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_67
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1604681595
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1604681595
transform 1 0 10396 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1604681595
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1604681595
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1604681595
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_143
timestamp 1604681595
transform 1 0 14260 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_30
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_38
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7084 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8648 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1604681595
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_91
timestamp 1604681595
transform 1 0 9476 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_97
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1604681595
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_143
timestamp 1604681595
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1604681595
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_16
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1604681595
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_16
timestamp 1604681595
transform 1 0 2576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_11
timestamp 1604681595
transform 1 0 2116 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2852 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_28
timestamp 1604681595
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_25
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_21
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_32
timestamp 1604681595
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4416 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_49
timestamp 1604681595
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_45
timestamp 1604681595
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_50
timestamp 1604681595
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_46
timestamp 1604681595
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_53
timestamp 1604681595
transform 1 0 5980 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_61
timestamp 1604681595
transform 1 0 6716 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5888 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7084 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_67
timestamp 1604681595
transform 1 0 7268 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_72
timestamp 1604681595
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1604681595
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_86
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_92
timestamp 1604681595
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_101
timestamp 1604681595
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_96
timestamp 1604681595
transform 1 0 9936 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1604681595
transform 1 0 11408 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_108
timestamp 1604681595
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11776 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_132
timestamp 1604681595
transform 1 0 13248 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_144
timestamp 1604681595
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_143
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_13
timestamp 1604681595
transform 1 0 2300 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 4324 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_38
timestamp 1604681595
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5336 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_42
timestamp 1604681595
transform 1 0 4968 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_62
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7544 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_67
timestamp 1604681595
transform 1 0 7268 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_79
timestamp 1604681595
transform 1 0 8372 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1604681595
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11960 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1604681595
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_113
timestamp 1604681595
transform 1 0 11500 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_120
timestamp 1604681595
transform 1 0 12144 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_132
timestamp 1604681595
transform 1 0 13248 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_144
timestamp 1604681595
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1604681595
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_35
timestamp 1604681595
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5060 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_52
timestamp 1604681595
transform 1 0 5888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1604681595
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_82
timestamp 1604681595
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1604681595
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1604681595
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_112
timestamp 1604681595
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_126
timestamp 1604681595
transform 1 0 12696 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_138
timestamp 1604681595
transform 1 0 13800 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_9
timestamp 1604681595
transform 1 0 1932 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1604681595
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4232 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_21
timestamp 1604681595
transform 1 0 3036 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6716 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_50
timestamp 1604681595
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1604681595
transform 1 0 6072 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_70
timestamp 1604681595
transform 1 0 7544 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11408 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1604681595
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1604681595
transform 1 0 11224 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_114
timestamp 1604681595
transform 1 0 11592 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_127
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_139
timestamp 1604681595
transform 1 0 13892 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2760 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_34
timestamp 1604681595
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1604681595
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4968 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7544 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1604681595
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_90
timestamp 1604681595
transform 1 0 9384 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_94
timestamp 1604681595
transform 1 0 9752 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_106
timestamp 1604681595
transform 1 0 10856 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_111
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_115
timestamp 1604681595
transform 1 0 11684 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_132
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1604681595
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1604681595
transform 1 0 2944 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_28
timestamp 1604681595
transform 1 0 3680 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_40
timestamp 1604681595
transform 1 0 4784 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_64
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_72
timestamp 1604681595
transform 1 0 7728 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_75
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_79
timestamp 1604681595
transform 1 0 8372 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1604681595
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_101
timestamp 1604681595
transform 1 0 10396 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1604681595
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4784 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 4324 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_37
timestamp 1604681595
transform 1 0 4508 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_50
timestamp 1604681595
transform 1 0 5704 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_42
timestamp 1604681595
transform 1 0 4968 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_52
timestamp 1604681595
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_47
timestamp 1604681595
transform 1 0 5428 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5888 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1604681595
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_56
timestamp 1604681595
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6440 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6072 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7820 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_78
timestamp 1604681595
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_82
timestamp 1604681595
transform 1 0 8648 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_63
timestamp 1604681595
transform 1 0 6900 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_69
timestamp 1604681595
transform 1 0 7452 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1604681595
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_86
timestamp 1604681595
transform 1 0 9016 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_90
timestamp 1604681595
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_97
timestamp 1604681595
transform 1 0 10028 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10212 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_115
timestamp 1604681595
transform 1 0 11684 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_34_125
timestamp 1604681595
transform 1 0 12604 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_132
timestamp 1604681595
transform 1 0 13248 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_144
timestamp 1604681595
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_137
timestamp 1604681595
transform 1 0 13708 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3496 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_23
timestamp 1604681595
transform 1 0 3220 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_28
timestamp 1604681595
transform 1 0 3680 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_36
timestamp 1604681595
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_49
timestamp 1604681595
transform 1 0 5612 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_54
timestamp 1604681595
transform 1 0 6072 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_58
timestamp 1604681595
transform 1 0 6440 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7268 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8648 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 7084 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8280 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_76
timestamp 1604681595
transform 1 0 8096 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_80
timestamp 1604681595
transform 1 0 8464 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8832 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_93
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_97
timestamp 1604681595
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_101
timestamp 1604681595
transform 1 0 10396 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 1604681595
transform 1 0 11500 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 1604681595
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_131
timestamp 1604681595
transform 1 0 13156 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_136
timestamp 1604681595
transform 1 0 13616 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_144
timestamp 1604681595
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2760 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_7
timestamp 1604681595
transform 1 0 1748 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_13
timestamp 1604681595
transform 1 0 2300 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_16
timestamp 1604681595
transform 1 0 2576 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_20
timestamp 1604681595
transform 1 0 2944 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4324 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3128 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1604681595
transform 1 0 3312 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_28
timestamp 1604681595
transform 1 0 3680 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5888 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 8096 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7912 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 7544 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_72
timestamp 1604681595
transform 1 0 7728 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_79
timestamp 1604681595
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_83
timestamp 1604681595
transform 1 0 8740 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1604681595
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_102
timestamp 1604681595
transform 1 0 10488 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_114
timestamp 1604681595
transform 1 0 11592 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 13432 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_126
timestamp 1604681595
transform 1 0 12696 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_138
timestamp 1604681595
transform 1 0 13800 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2760 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2208 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_9
timestamp 1604681595
transform 1 0 1932 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_14
timestamp 1604681595
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4324 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3772 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_31
timestamp 1604681595
transform 1 0 3956 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_44
timestamp 1604681595
transform 1 0 5152 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5336 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_48
timestamp 1604681595
transform 1 0 5520 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5704 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_56
timestamp 1604681595
transform 1 0 6256 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_52
timestamp 1604681595
transform 1 0 5888 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6072 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_60
timestamp 1604681595
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6440 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7360 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7176 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9568 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_84
timestamp 1604681595
transform 1 0 8832 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_88
timestamp 1604681595
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_101
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12604 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_105
timestamp 1604681595
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_109
timestamp 1604681595
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1604681595
transform 1 0 11500 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1604681595
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12972 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_127
timestamp 1604681595
transform 1 0 12788 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_131
timestamp 1604681595
transform 1 0 13156 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_143
timestamp 1604681595
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_11
timestamp 1604681595
transform 1 0 2116 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4140 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_23
timestamp 1604681595
transform 1 0 3220 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6440 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_38_49
timestamp 1604681595
transform 1 0 5612 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_57
timestamp 1604681595
transform 1 0 6348 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_67
timestamp 1604681595
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_71
timestamp 1604681595
transform 1 0 7636 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_84
timestamp 1604681595
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12328 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_109
timestamp 1604681595
transform 1 0 11132 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_113
timestamp 1604681595
transform 1 0 11500 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_121
timestamp 1604681595
transform 1 0 12236 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_138
timestamp 1604681595
transform 1 0 13800 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 3036 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 3036 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_37
timestamp 1604681595
transform 1 0 4508 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_41
timestamp 1604681595
transform 1 0 4876 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_23
timestamp 1604681595
transform 1 0 3220 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_40
timestamp 1604681595
transform 1 0 4784 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_45
timestamp 1604681595
transform 1 0 5244 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_48
timestamp 1604681595
transform 1 0 5520 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5060 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5060 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5704 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5336 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 5244 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_59
timestamp 1604681595
transform 1 0 6532 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_55
timestamp 1604681595
transform 1 0 6164 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_52
timestamp 1604681595
transform 1 0 5888 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6348 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6716 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_83
timestamp 1604681595
transform 1 0 8740 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_79
timestamp 1604681595
transform 1 0 8372 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_77
timestamp 1604681595
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_73
timestamp 1604681595
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8556 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6900 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_88
timestamp 1604681595
transform 1 0 9200 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_90
timestamp 1604681595
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_101
timestamp 1604681595
transform 1 0 10396 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_97
timestamp 1604681595
transform 1 0 10028 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_94
timestamp 1604681595
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10212 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10580 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_123
timestamp 1604681595
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10948 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 13156 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_132
timestamp 1604681595
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_136
timestamp 1604681595
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_140
timestamp 1604681595
transform 1 0 13984 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_127
timestamp 1604681595
transform 1 0 12788 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_134
timestamp 1604681595
transform 1 0 13432 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_19
timestamp 1604681595
transform 1 0 2852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4876 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4508 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3680 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_30
timestamp 1604681595
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_34
timestamp 1604681595
transform 1 0 4232 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5060 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_52
timestamp 1604681595
transform 1 0 5888 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7084 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_82
timestamp 1604681595
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_95
timestamp 1604681595
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_99
timestamp 1604681595
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_112
timestamp 1604681595
transform 1 0 11408 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_132
timestamp 1604681595
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_136
timestamp 1604681595
transform 1 0 13616 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_144
timestamp 1604681595
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_9
timestamp 1604681595
transform 1 0 1932 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_21
timestamp 1604681595
transform 1 0 3036 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1604681595
transform 1 0 3772 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5704 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_48
timestamp 1604681595
transform 1 0 5520 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_52
timestamp 1604681595
transform 1 0 5888 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_59
timestamp 1604681595
transform 1 0 6532 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7084 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_67
timestamp 1604681595
transform 1 0 7268 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_71
timestamp 1604681595
transform 1 0 7636 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_83
timestamp 1604681595
transform 1 0 8740 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10580 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10120 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_88
timestamp 1604681595
transform 1 0 9200 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_97
timestamp 1604681595
transform 1 0 10028 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_100
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12144 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11592 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_112
timestamp 1604681595
transform 1 0 11408 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_116
timestamp 1604681595
transform 1 0 11776 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13156 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_129
timestamp 1604681595
transform 1 0 12972 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_133
timestamp 1604681595
transform 1 0 13340 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_145
timestamp 1604681595
transform 1 0 14444 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604681595
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2484 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_9
timestamp 1604681595
transform 1 0 1932 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_13
timestamp 1604681595
transform 1 0 2300 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_17
timestamp 1604681595
transform 1 0 2668 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_29
timestamp 1604681595
transform 1 0 3772 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_34
timestamp 1604681595
transform 1 0 4232 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_38
timestamp 1604681595
transform 1 0 4600 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_42
timestamp 1604681595
transform 1 0 4968 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_53
timestamp 1604681595
transform 1 0 5980 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1604681595
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_62
timestamp 1604681595
transform 1 0 6808 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 7360 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1604681595
transform 1 0 7544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_82
timestamp 1604681595
transform 1 0 8648 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10120 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 9844 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9660 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9292 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8924 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_87
timestamp 1604681595
transform 1 0 9108 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_91
timestamp 1604681595
transform 1 0 9476 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11132 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 11500 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_107
timestamp 1604681595
transform 1 0 10948 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_111
timestamp 1604681595
transform 1 0 11316 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_115
timestamp 1604681595
transform 1 0 11684 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_121
timestamp 1604681595
transform 1 0 12236 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1604681595
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_135
timestamp 1604681595
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_143
timestamp 1604681595
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604681595
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604681595
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_9
timestamp 1604681595
transform 1 0 1932 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_21
timestamp 1604681595
transform 1 0 3036 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1604681595
transform 1 0 3772 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_41
timestamp 1604681595
transform 1 0 4876 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 5888 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 5152 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5520 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_46
timestamp 1604681595
transform 1 0 5336 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_50
timestamp 1604681595
transform 1 0 5704 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7544 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 7912 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_68
timestamp 1604681595
transform 1 0 7360 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_72
timestamp 1604681595
transform 1 0 7728 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_76
timestamp 1604681595
transform 1 0 8096 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_88
timestamp 1604681595
transform 1 0 9200 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_102
timestamp 1604681595
transform 1 0 10488 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_106
timestamp 1604681595
transform 1 0 10856 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_110
timestamp 1604681595
transform 1 0 11224 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_122
timestamp 1604681595
transform 1 0 12328 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_134
timestamp 1604681595
transform 1 0 13432 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604681595
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604681595
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1604681595
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_15
timestamp 1604681595
transform 1 0 2484 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4232 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4048 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3680 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3312 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_23
timestamp 1604681595
transform 1 0 3220 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_26
timestamp 1604681595
transform 1 0 3496 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_30
timestamp 1604681595
transform 1 0 3864 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 5888 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6256 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_50
timestamp 1604681595
transform 1 0 5704 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1604681595
transform 1 0 6072 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_62
timestamp 1604681595
transform 1 0 6808 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7452 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7268 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_66
timestamp 1604681595
transform 1 0 7176 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9936 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9568 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9200 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_85
timestamp 1604681595
transform 1 0 8924 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_90
timestamp 1604681595
transform 1 0 9384 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_94
timestamp 1604681595
transform 1 0 9752 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_98
timestamp 1604681595
transform 1 0 10120 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11500 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11868 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_110
timestamp 1604681595
transform 1 0 11224 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_115
timestamp 1604681595
transform 1 0 11684 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_119
timestamp 1604681595
transform 1 0 12052 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1604681595
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_135
timestamp 1604681595
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_143
timestamp 1604681595
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604681595
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 1380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604681595
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604681595
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 1932 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1604681595
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1604681595
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_7
timestamp 1604681595
transform 1 0 1748 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_11
timestamp 1604681595
transform 1 0 2116 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_19
timestamp 1604681595
transform 1 0 2852 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_23
timestamp 1604681595
transform 1 0 3220 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1604681595
transform 1 0 3772 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3036 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3588 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_40
timestamp 1604681595
transform 1 0 4784 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_36
timestamp 1604681595
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_40
timestamp 1604681595
transform 1 0 4784 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_36
timestamp 1604681595
transform 1 0 4416 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_32
timestamp 1604681595
transform 1 0 4048 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4968 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_62
timestamp 1604681595
transform 1 0 6808 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1604681595
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_53
timestamp 1604681595
transform 1 0 5980 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_60
timestamp 1604681595
transform 1 0 6624 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6164 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5152 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_46_66
timestamp 1604681595
transform 1 0 7176 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6992 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6992 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_81
timestamp 1604681595
transform 1 0 8556 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_77
timestamp 1604681595
transform 1 0 8188 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_73
timestamp 1604681595
transform 1 0 7820 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8372 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8004 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 8740 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 1604681595
transform 1 0 9660 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_88
timestamp 1604681595
transform 1 0 9200 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_84
timestamp 1604681595
transform 1 0 8832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_102
timestamp 1604681595
transform 1 0 10488 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10672 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9936 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9016 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_47_114
timestamp 1604681595
transform 1 0 11592 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1604681595
transform 1 0 11224 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_106
timestamp 1604681595
transform 1 0 10856 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_109
timestamp 1604681595
transform 1 0 11132 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_105
timestamp 1604681595
transform 1 0 10764 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10948 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11408 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1604681595
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11500 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_46_129
timestamp 1604681595
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1604681595
transform 1 0 14076 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_145
timestamp 1604681595
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1604681595
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_143
timestamp 1604681595
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604681595
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604681595
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604681595
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_3
timestamp 1604681595
transform 1 0 1380 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_11
timestamp 1604681595
transform 1 0 2116 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_16
timestamp 1604681595
transform 1 0 2576 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_24
timestamp 1604681595
transform 1 0 3312 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1604681595
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_41
timestamp 1604681595
transform 1 0 4876 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 5704 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5060 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5428 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6256 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_45
timestamp 1604681595
transform 1 0 5244 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_49
timestamp 1604681595
transform 1 0 5612 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_53
timestamp 1604681595
transform 1 0 5980 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_58
timestamp 1604681595
transform 1 0 6440 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_62
timestamp 1604681595
transform 1 0 6808 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7084 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6900 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8096 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 8464 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_74
timestamp 1604681595
transform 1 0 7912 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_78
timestamp 1604681595
transform 1 0 8280 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_82
timestamp 1604681595
transform 1 0 8648 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10304 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9108 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_86
timestamp 1604681595
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_89
timestamp 1604681595
transform 1 0 9292 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1604681595
transform 1 0 9660 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_97
timestamp 1604681595
transform 1 0 10028 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1604681595
transform 1 0 11132 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1604681595
transform 1 0 12236 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_133
timestamp 1604681595
transform 1 0 13340 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1604681595
transform 1 0 14444 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604681595
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604681595
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 1932 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_7
timestamp 1604681595
transform 1 0 1748 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_11
timestamp 1604681595
transform 1 0 2116 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_16
timestamp 1604681595
transform 1 0 2576 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_20
timestamp 1604681595
transform 1 0 2944 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3404 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3220 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4692 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_34
timestamp 1604681595
transform 1 0 4232 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_38
timestamp 1604681595
transform 1 0 4600 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_41
timestamp 1604681595
transform 1 0 4876 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6256 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1604681595
transform 1 0 5980 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_58
timestamp 1604681595
transform 1 0 6440 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_62
timestamp 1604681595
transform 1 0 6808 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 7268 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 8280 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6992 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_66
timestamp 1604681595
transform 1 0 7176 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_70
timestamp 1604681595
transform 1 0 7544 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_74
timestamp 1604681595
transform 1 0 7912 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_77
timestamp 1604681595
transform 1 0 8188 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_81
timestamp 1604681595
transform 1 0 8556 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 10120 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 10488 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_96
timestamp 1604681595
transform 1 0 9936 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_100
timestamp 1604681595
transform 1 0 10304 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_104
timestamp 1604681595
transform 1 0 10672 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10856 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11224 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_108
timestamp 1604681595
transform 1 0 11040 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_112
timestamp 1604681595
transform 1 0 11408 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_120
timestamp 1604681595
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1604681595
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1604681595
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_143
timestamp 1604681595
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604681595
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604681595
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1604681595
transform 1 0 1380 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_11
timestamp 1604681595
transform 1 0 2116 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4692 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4232 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_23
timestamp 1604681595
transform 1 0 3220 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_27
timestamp 1604681595
transform 1 0 3588 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_32
timestamp 1604681595
transform 1 0 4048 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_36
timestamp 1604681595
transform 1 0 4416 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6256 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 5704 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6072 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_48
timestamp 1604681595
transform 1 0 5520 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_52
timestamp 1604681595
transform 1 0 5888 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7360 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7728 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_65
timestamp 1604681595
transform 1 0 7084 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_70
timestamp 1604681595
transform 1 0 7544 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_74
timestamp 1604681595
transform 1 0 7912 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 10396 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9108 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_84
timestamp 1604681595
transform 1 0 8832 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_89
timestamp 1604681595
transform 1 0 9292 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_93
timestamp 1604681595
transform 1 0 9660 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_104
timestamp 1604681595
transform 1 0 10672 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10856 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_122
timestamp 1604681595
transform 1 0 12328 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_134
timestamp 1604681595
transform 1 0 13432 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604681595
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2852 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604681595
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2668 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_9
timestamp 1604681595
transform 1 0 1932 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_13
timestamp 1604681595
transform 1 0 2300 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4876 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4508 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_35
timestamp 1604681595
transform 1 0 4324 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_39
timestamp 1604681595
transform 1 0 4692 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5060 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_52
timestamp 1604681595
transform 1 0 5888 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1604681595
transform 1 0 6348 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_62
timestamp 1604681595
transform 1 0 6808 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7360 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8740 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6992 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8372 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_66
timestamp 1604681595
transform 1 0 7176 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_77
timestamp 1604681595
transform 1 0 8188 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_81
timestamp 1604681595
transform 1 0 8556 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8924 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10488 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10304 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9936 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_94
timestamp 1604681595
transform 1 0 9752 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_98
timestamp 1604681595
transform 1 0 10120 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11500 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 11868 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_111
timestamp 1604681595
transform 1 0 11316 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_115
timestamp 1604681595
transform 1 0 11684 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_119
timestamp 1604681595
transform 1 0 12052 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1604681595
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1604681595
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_143
timestamp 1604681595
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604681595
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604681595
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604681595
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 2852 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1604681595
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1604681595
transform 1 0 2484 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1604681595
transform 1 0 1380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_7
timestamp 1604681595
transform 1 0 1748 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_19
timestamp 1604681595
transform 1 0 2852 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 3680 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 3496 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_21
timestamp 1604681595
transform 1 0 3036 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_41
timestamp 1604681595
transform 1 0 4876 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_25
timestamp 1604681595
transform 1 0 3404 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_48
timestamp 1604681595
transform 1 0 5520 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_44
timestamp 1604681595
transform 1 0 5152 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_45
timestamp 1604681595
transform 1 0 5244 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5704 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5336 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5060 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 5612 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_58
timestamp 1604681595
transform 1 0 6440 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_52
timestamp 1604681595
transform 1 0 5888 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_52
timestamp 1604681595
transform 1 0 5888 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6624 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_53_62
timestamp 1604681595
transform 1 0 6808 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_67
timestamp 1604681595
transform 1 0 7268 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_69
timestamp 1604681595
transform 1 0 7452 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7084 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7452 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7636 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_80
timestamp 1604681595
transform 1 0 8464 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_77
timestamp 1604681595
transform 1 0 8188 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_73
timestamp 1604681595
transform 1 0 7820 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_84
timestamp 1604681595
transform 1 0 8832 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_93
timestamp 1604681595
transform 1 0 9660 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1604681595
transform 1 0 9476 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_87
timestamp 1604681595
transform 1 0 9108 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9568 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8924 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_94
timestamp 1604681595
transform 1 0 9752 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_100
timestamp 1604681595
transform 1 0 10304 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_97
timestamp 1604681595
transform 1 0 10028 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9936 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10396 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_53_111
timestamp 1604681595
transform 1 0 11316 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_107
timestamp 1604681595
transform 1 0 10948 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11500 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11132 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_119
timestamp 1604681595
transform 1 0 12052 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_115
timestamp 1604681595
transform 1 0 11684 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11868 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_123
timestamp 1604681595
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_117
timestamp 1604681595
transform 1 0 11868 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_129
timestamp 1604681595
transform 1 0 12972 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1604681595
transform 1 0 14076 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_145
timestamp 1604681595
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_135
timestamp 1604681595
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_143
timestamp 1604681595
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604681595
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604681595
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604681595
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_9
timestamp 1604681595
transform 1 0 1932 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4876 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4692 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 3680 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1604681595
transform 1 0 3036 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1604681595
transform 1 0 3588 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_30
timestamp 1604681595
transform 1 0 3864 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_32
timestamp 1604681595
transform 1 0 4048 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_38
timestamp 1604681595
transform 1 0 4600 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_57
timestamp 1604681595
transform 1 0 6348 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_61
timestamp 1604681595
transform 1 0 6716 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7360 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7176 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_64
timestamp 1604681595
transform 1 0 6992 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 9660 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10120 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_84
timestamp 1604681595
transform 1 0 8832 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_96
timestamp 1604681595
transform 1 0 9936 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_100
timestamp 1604681595
transform 1 0 10304 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_104
timestamp 1604681595
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11040 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12052 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10856 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_117
timestamp 1604681595
transform 1 0 11868 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1604681595
transform 1 0 12236 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_133
timestamp 1604681595
transform 1 0 13340 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_145
timestamp 1604681595
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604681595
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604681595
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1604681595
transform 1 0 1380 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_7
timestamp 1604681595
transform 1 0 1748 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_19
timestamp 1604681595
transform 1 0 2852 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4232 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_31
timestamp 1604681595
transform 1 0 3956 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_36
timestamp 1604681595
transform 1 0 4416 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_40
timestamp 1604681595
transform 1 0 4784 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_53
timestamp 1604681595
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1604681595
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8648 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8280 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 7820 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_71
timestamp 1604681595
transform 1 0 7636 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_75
timestamp 1604681595
transform 1 0 8004 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_80
timestamp 1604681595
transform 1 0 8464 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8832 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10488 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10304 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_93
timestamp 1604681595
transform 1 0 9660 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_98
timestamp 1604681595
transform 1 0 10120 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 12420 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 11500 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11868 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_111
timestamp 1604681595
transform 1 0 11316 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_115
timestamp 1604681595
transform 1 0 11684 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_119
timestamp 1604681595
transform 1 0 12052 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_126
timestamp 1604681595
transform 1 0 12696 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_138
timestamp 1604681595
transform 1 0 13800 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604681595
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604681595
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 2484 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_9
timestamp 1604681595
transform 1 0 1932 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_17
timestamp 1604681595
transform 1 0 2668 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4876 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1604681595
transform 1 0 3772 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_32
timestamp 1604681595
transform 1 0 4048 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_40
timestamp 1604681595
transform 1 0 4784 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6624 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5060 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_56_52
timestamp 1604681595
transform 1 0 5888 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_76
timestamp 1604681595
transform 1 0 8096 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8832 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_86
timestamp 1604681595
transform 1 0 9016 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_93
timestamp 1604681595
transform 1 0 9660 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11500 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12512 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_105
timestamp 1604681595
transform 1 0 10764 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_122
timestamp 1604681595
transform 1 0 12328 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_126
timestamp 1604681595
transform 1 0 12696 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_138
timestamp 1604681595
transform 1 0 13800 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604681595
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 2484 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 1380 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604681595
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 1932 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 2300 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_7
timestamp 1604681595
transform 1 0 1748 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_11
timestamp 1604681595
transform 1 0 2116 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_19
timestamp 1604681595
transform 1 0 2852 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 3036 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 4140 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_23
timestamp 1604681595
transform 1 0 3220 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_31
timestamp 1604681595
transform 1 0 3956 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_35
timestamp 1604681595
transform 1 0 4324 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 5796 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_45
timestamp 1604681595
transform 1 0 5244 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_53
timestamp 1604681595
transform 1 0 5980 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_62
timestamp 1604681595
transform 1 0 6808 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 7176 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 7728 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 8096 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8556 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_70
timestamp 1604681595
transform 1 0 7544 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_74
timestamp 1604681595
transform 1 0 7912 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_78
timestamp 1604681595
transform 1 0 8280 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_83
timestamp 1604681595
transform 1 0 8740 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9476 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10488 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_87
timestamp 1604681595
transform 1 0 9108 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_100
timestamp 1604681595
transform 1 0 10304 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_104
timestamp 1604681595
transform 1 0 10672 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11776 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11408 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1604681595
transform 1 0 11224 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_114
timestamp 1604681595
transform 1 0 11592 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_118
timestamp 1604681595
transform 1 0 11960 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_132
timestamp 1604681595
transform 1 0 13248 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_136
timestamp 1604681595
transform 1 0 13616 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_144
timestamp 1604681595
transform 1 0 14352 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604681595
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 2484 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 1380 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604681595
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_7
timestamp 1604681595
transform 1 0 1748 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_19
timestamp 1604681595
transform 1 0 2852 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 4140 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_32
timestamp 1604681595
transform 1 0 4048 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_37
timestamp 1604681595
transform 1 0 4508 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 5796 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_49
timestamp 1604681595
transform 1 0 5612 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_55
timestamp 1604681595
transform 1 0 6164 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 7544 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_67
timestamp 1604681595
transform 1 0 7268 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_74
timestamp 1604681595
transform 1 0 7912 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9752 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_86
timestamp 1604681595
transform 1 0 9016 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_93
timestamp 1604681595
transform 1 0 9660 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11960 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11408 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_110
timestamp 1604681595
transform 1 0 11224 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_114
timestamp 1604681595
transform 1 0 11592 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_127
timestamp 1604681595
transform 1 0 12788 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_139
timestamp 1604681595
transform 1 0 13892 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_145
timestamp 1604681595
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604681595
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_7
timestamp 1604681595
transform 1 0 1748 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604681595
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604681595
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 1380 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_15
timestamp 1604681595
transform 1 0 2484 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_19
timestamp 1604681595
transform 1 0 2852 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_11
timestamp 1604681595
transform 1 0 2116 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 2300 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 2484 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 2852 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1604681595
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_23
timestamp 1604681595
transform 1 0 3220 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_23
timestamp 1604681595
transform 1 0 3220 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 3404 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 3036 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 3588 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_36
timestamp 1604681595
transform 1 0 4416 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_35
timestamp 1604681595
transform 1 0 4324 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_31
timestamp 1604681595
transform 1 0 3956 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 4140 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 4048 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_48
timestamp 1604681595
transform 1 0 5520 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_46
timestamp 1604681595
transform 1 0 5336 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_43
timestamp 1604681595
transform 1 0 5060 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 5152 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 5152 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 5520 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_56
timestamp 1604681595
transform 1 0 6256 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_56
timestamp 1604681595
transform 1 0 6256 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_52
timestamp 1604681595
transform 1 0 5888 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 6440 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 6072 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 6348 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_61
timestamp 1604681595
transform 1 0 6716 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_62
timestamp 1604681595
transform 1 0 6808 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_60
timestamp 1604681595
transform 1 0 6624 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_67
timestamp 1604681595
transform 1 0 7268 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_71
timestamp 1604681595
transform 1 0 7636 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_67
timestamp 1604681595
transform 1 0 7268 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 7084 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 7452 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 7084 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 7452 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_73
timestamp 1604681595
transform 1 0 7820 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 8004 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_77
timestamp 1604681595
transform 1 0 8188 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 7820 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10028 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9844 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10028 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_89
timestamp 1604681595
transform 1 0 9292 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_89
timestamp 1604681595
transform 1 0 9292 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_93
timestamp 1604681595
transform 1 0 9660 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_99
timestamp 1604681595
transform 1 0 10212 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11040 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11684 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1604681595
transform 1 0 11500 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_117
timestamp 1604681595
transform 1 0 11868 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_121
timestamp 1604681595
transform 1 0 12236 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_123
timestamp 1604681595
transform 1 0 12420 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_107
timestamp 1604681595
transform 1 0 10948 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_124
timestamp 1604681595
transform 1 0 12512 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 13432 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 13984 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_131
timestamp 1604681595
transform 1 0 13156 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_138
timestamp 1604681595
transform 1 0 13800 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_142
timestamp 1604681595
transform 1 0 14168 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_136
timestamp 1604681595
transform 1 0 13616 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_144
timestamp 1604681595
transform 1 0 14352 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604681595
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604681595
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604681595
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604681595
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1604681595
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1604681595
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_39
timestamp 1604681595
transform 1 0 4692 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 5152 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 5704 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_43
timestamp 1604681595
transform 1 0 5060 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_48
timestamp 1604681595
transform 1 0 5520 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_52
timestamp 1604681595
transform 1 0 5888 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_60
timestamp 1604681595
transform 1 0 6624 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_62
timestamp 1604681595
transform 1 0 6808 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 7084 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 7636 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_69
timestamp 1604681595
transform 1 0 7452 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_73
timestamp 1604681595
transform 1 0 7820 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_85
timestamp 1604681595
transform 1 0 8924 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_97
timestamp 1604681595
transform 1 0 10028 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_109
timestamp 1604681595
transform 1 0 11132 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_121
timestamp 1604681595
transform 1 0 12236 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1604681595
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1604681595
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_143
timestamp 1604681595
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604681595
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604681595
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604681595
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604681595
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604681595
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1604681595
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1604681595
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_56
timestamp 1604681595
transform 1 0 6256 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 7084 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_64
timestamp 1604681595
transform 1 0 6992 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_69
timestamp 1604681595
transform 1 0 7452 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_81
timestamp 1604681595
transform 1 0 8556 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_89
timestamp 1604681595
transform 1 0 9292 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604681595
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1604681595
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1604681595
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1604681595
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1604681595
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1604681595
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604681595
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604681595
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604681595
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604681595
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604681595
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1604681595
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1604681595
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1604681595
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1604681595
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1604681595
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1604681595
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1604681595
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1604681595
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604681595
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1604681595
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_143
timestamp 1604681595
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604681595
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604681595
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604681595
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604681595
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604681595
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604681595
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604681595
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604681595
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604681595
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604681595
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604681595
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604681595
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604681595
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604681595
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604681595
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_137
timestamp 1604681595
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1604681595
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604681595
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 2864 480 2984 6 ccff_head
port 0 nsew default input
rlabel metal3 s 15520 9936 16000 10056 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8206 39520 8262 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12162 39520 12218 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 12990 39520 13046 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 13358 39520 13414 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14922 39520 14978 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15750 39520 15806 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 8942 39520 8998 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9402 39520 9458 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 9770 39520 9826 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10598 39520 10654 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 10966 39520 11022 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 11794 39520 11850 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 39520 258 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4158 39520 4214 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5354 39520 5410 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6182 39520 6238 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 6918 39520 6974 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 7746 39520 7802 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 938 39520 994 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 39520 1454 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1766 39520 1822 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2594 39520 2650 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 2962 39520 3018 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3790 39520 3846 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 15520 23264 16000 23384 6 gfpga_pad_EMBEDDED_IO_SOC_DIR
port 82 nsew default tristate
rlabel metal3 s 15520 29928 16000 30048 6 gfpga_pad_EMBEDDED_IO_SOC_IN
port 83 nsew default input
rlabel metal3 s 15520 36592 16000 36712 6 gfpga_pad_EMBEDDED_IO_SOC_OUT
port 84 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 left_grid_pin_16_
port 85 nsew default tristate
rlabel metal3 s 0 6944 480 7064 6 left_grid_pin_17_
port 86 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 left_grid_pin_18_
port 87 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 left_grid_pin_19_
port 88 nsew default tristate
rlabel metal3 s 0 12928 480 13048 6 left_grid_pin_20_
port 89 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 left_grid_pin_21_
port 90 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 left_grid_pin_22_
port 91 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 left_grid_pin_23_
port 92 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 left_grid_pin_24_
port 93 nsew default tristate
rlabel metal3 s 0 22856 480 22976 6 left_grid_pin_25_
port 94 nsew default tristate
rlabel metal3 s 0 24896 480 25016 6 left_grid_pin_26_
port 95 nsew default tristate
rlabel metal3 s 0 26936 480 27056 6 left_grid_pin_27_
port 96 nsew default tristate
rlabel metal3 s 0 28840 480 28960 6 left_grid_pin_28_
port 97 nsew default tristate
rlabel metal3 s 0 30880 480 31000 6 left_grid_pin_29_
port 98 nsew default tristate
rlabel metal3 s 0 32920 480 33040 6 left_grid_pin_30_
port 99 nsew default tristate
rlabel metal3 s 0 34824 480 34944 6 left_grid_pin_31_
port 100 nsew default tristate
rlabel metal3 s 0 36864 480 36984 6 left_width_0_height_0__pin_0_
port 101 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_width_0_height_0__pin_1_lower
port 102 nsew default tristate
rlabel metal3 s 0 38904 480 39024 6 left_width_0_height_0__pin_1_upper
port 103 nsew default tristate
rlabel metal3 s 15520 3272 16000 3392 6 prog_clk
port 104 nsew default input
rlabel metal3 s 15520 16600 16000 16720 6 right_grid_pin_0_
port 105 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 VPWR
port 106 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 VGND
port 107 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
