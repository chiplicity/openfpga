VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__2_
  CLASS BLOCK ;
  FOREIGN cbx_1__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 85.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 81.000 5.890 85.000 ;
    END
  END IO_ISOL_N
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 81.000 16.930 85.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 81.000 27.970 85.000 ;
    END
  END SC_OUT_TOP
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END bottom_grid_pin_11_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END bottom_grid_pin_13_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END bottom_grid_pin_15_
  PIN bottom_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END bottom_grid_pin_1_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END bottom_grid_pin_3_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END bottom_grid_pin_5_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END bottom_grid_pin_7_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END bottom_grid_pin_8_
  PIN bottom_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END bottom_grid_pin_9_
  PIN bottom_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END bottom_width_0_height_0__pin_0_
  PIN bottom_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END bottom_width_0_height_0__pin_1_lower
  PIN bottom_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END bottom_width_0_height_0__pin_1_upper
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 81.000 39.010 85.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 81.000 50.050 85.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 42.880 100.000 43.480 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 63.960 100.000 64.560 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 66.000 100.000 66.600 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 68.720 100.000 69.320 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 70.760 100.000 71.360 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 72.800 100.000 73.400 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 74.840 100.000 75.440 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 76.880 100.000 77.480 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 78.920 100.000 79.520 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 80.960 100.000 81.560 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 83.000 100.000 83.600 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 44.920 100.000 45.520 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 46.960 100.000 47.560 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 49.000 100.000 49.600 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 51.720 100.000 52.320 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 53.760 100.000 54.360 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.800 100.000 56.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 57.840 100.000 58.440 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 59.880 100.000 60.480 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 61.920 100.000 62.520 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 0.720 100.000 1.320 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 21.800 100.000 22.400 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 23.840 100.000 24.440 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 25.880 100.000 26.480 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 27.920 100.000 28.520 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 29.960 100.000 30.560 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 32.000 100.000 32.600 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 34.720 100.000 35.320 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 36.760 100.000 37.360 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 38.800 100.000 39.400 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 40.840 100.000 41.440 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 2.760 100.000 3.360 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 4.800 100.000 5.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 6.840 100.000 7.440 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 8.880 100.000 9.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 10.920 100.000 11.520 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 12.960 100.000 13.560 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 15.000 100.000 15.600 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 17.720 100.000 18.320 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 19.760 100.000 20.360 ;
    END
  END chanx_right_out[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.850 81.000 72.130 85.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 81.000 83.170 85.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 81.000 94.210 85.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END prog_clk_0_S_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END prog_clk_0_W_out
  PIN top_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 81.000 61.090 85.000 ;
    END
  END top_grid_pin_0_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.545 10.640 21.145 73.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.375 10.640 35.975 73.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 73.525 ;
      LAYER met1 ;
        RECT 1.910 6.840 94.300 76.800 ;
      LAYER met2 ;
        RECT 1.940 80.720 5.330 83.485 ;
        RECT 6.170 80.720 16.370 83.485 ;
        RECT 17.210 80.720 27.410 83.485 ;
        RECT 28.250 80.720 38.450 83.485 ;
        RECT 39.290 80.720 49.490 83.485 ;
        RECT 50.330 80.720 60.530 83.485 ;
        RECT 61.370 80.720 71.570 83.485 ;
        RECT 72.410 80.720 82.610 83.485 ;
        RECT 83.450 80.720 93.650 83.485 ;
        RECT 94.490 80.720 97.430 83.485 ;
        RECT 1.940 4.280 97.430 80.720 ;
        RECT 2.490 0.835 5.790 4.280 ;
        RECT 6.630 0.835 10.390 4.280 ;
        RECT 11.230 0.835 14.990 4.280 ;
        RECT 15.830 0.835 19.590 4.280 ;
        RECT 20.430 0.835 24.190 4.280 ;
        RECT 25.030 0.835 28.790 4.280 ;
        RECT 29.630 0.835 33.390 4.280 ;
        RECT 34.230 0.835 37.530 4.280 ;
        RECT 38.370 0.835 42.130 4.280 ;
        RECT 42.970 0.835 46.730 4.280 ;
        RECT 47.570 0.835 51.330 4.280 ;
        RECT 52.170 0.835 55.930 4.280 ;
        RECT 56.770 0.835 60.530 4.280 ;
        RECT 61.370 0.835 65.130 4.280 ;
        RECT 65.970 0.835 69.270 4.280 ;
        RECT 70.110 0.835 73.870 4.280 ;
        RECT 74.710 0.835 78.470 4.280 ;
        RECT 79.310 0.835 83.070 4.280 ;
        RECT 83.910 0.835 87.670 4.280 ;
        RECT 88.510 0.835 92.270 4.280 ;
        RECT 93.110 0.835 96.870 4.280 ;
      LAYER met3 ;
        RECT 4.400 82.600 95.600 83.465 ;
        RECT 4.000 81.960 97.455 82.600 ;
        RECT 4.400 80.560 95.600 81.960 ;
        RECT 4.000 79.920 97.455 80.560 ;
        RECT 4.400 78.520 95.600 79.920 ;
        RECT 4.000 77.880 97.455 78.520 ;
        RECT 4.400 76.480 95.600 77.880 ;
        RECT 4.000 75.840 97.455 76.480 ;
        RECT 4.400 74.440 95.600 75.840 ;
        RECT 4.000 73.800 97.455 74.440 ;
        RECT 4.400 72.400 95.600 73.800 ;
        RECT 4.000 71.760 97.455 72.400 ;
        RECT 4.400 70.360 95.600 71.760 ;
        RECT 4.000 69.720 97.455 70.360 ;
        RECT 4.400 68.320 95.600 69.720 ;
        RECT 4.000 67.680 97.455 68.320 ;
        RECT 4.400 67.000 97.455 67.680 ;
        RECT 4.400 66.280 95.600 67.000 ;
        RECT 4.000 65.640 95.600 66.280 ;
        RECT 4.400 65.600 95.600 65.640 ;
        RECT 4.400 64.960 97.455 65.600 ;
        RECT 4.400 64.240 95.600 64.960 ;
        RECT 4.000 63.600 95.600 64.240 ;
        RECT 4.400 63.560 95.600 63.600 ;
        RECT 4.400 62.920 97.455 63.560 ;
        RECT 4.400 62.200 95.600 62.920 ;
        RECT 4.000 61.560 95.600 62.200 ;
        RECT 4.400 61.520 95.600 61.560 ;
        RECT 4.400 60.880 97.455 61.520 ;
        RECT 4.400 60.160 95.600 60.880 ;
        RECT 4.000 59.520 95.600 60.160 ;
        RECT 4.400 59.480 95.600 59.520 ;
        RECT 4.400 58.840 97.455 59.480 ;
        RECT 4.400 58.120 95.600 58.840 ;
        RECT 4.000 57.480 95.600 58.120 ;
        RECT 4.400 57.440 95.600 57.480 ;
        RECT 4.400 56.800 97.455 57.440 ;
        RECT 4.400 56.080 95.600 56.800 ;
        RECT 4.000 55.440 95.600 56.080 ;
        RECT 4.400 55.400 95.600 55.440 ;
        RECT 4.400 54.760 97.455 55.400 ;
        RECT 4.400 54.040 95.600 54.760 ;
        RECT 4.000 53.400 95.600 54.040 ;
        RECT 4.400 53.360 95.600 53.400 ;
        RECT 4.400 52.720 97.455 53.360 ;
        RECT 4.400 52.000 95.600 52.720 ;
        RECT 4.000 51.360 95.600 52.000 ;
        RECT 4.400 51.320 95.600 51.360 ;
        RECT 4.400 50.000 97.455 51.320 ;
        RECT 4.400 49.960 95.600 50.000 ;
        RECT 4.000 49.320 95.600 49.960 ;
        RECT 4.400 48.600 95.600 49.320 ;
        RECT 4.400 47.960 97.455 48.600 ;
        RECT 4.400 47.920 95.600 47.960 ;
        RECT 4.000 47.280 95.600 47.920 ;
        RECT 4.400 46.560 95.600 47.280 ;
        RECT 4.400 45.920 97.455 46.560 ;
        RECT 4.400 45.880 95.600 45.920 ;
        RECT 4.000 45.240 95.600 45.880 ;
        RECT 4.400 44.520 95.600 45.240 ;
        RECT 4.400 43.880 97.455 44.520 ;
        RECT 4.400 43.840 95.600 43.880 ;
        RECT 4.000 42.520 95.600 43.840 ;
        RECT 4.400 42.480 95.600 42.520 ;
        RECT 4.400 41.840 97.455 42.480 ;
        RECT 4.400 41.120 95.600 41.840 ;
        RECT 4.000 40.480 95.600 41.120 ;
        RECT 4.400 40.440 95.600 40.480 ;
        RECT 4.400 39.800 97.455 40.440 ;
        RECT 4.400 39.080 95.600 39.800 ;
        RECT 4.000 38.440 95.600 39.080 ;
        RECT 4.400 38.400 95.600 38.440 ;
        RECT 4.400 37.760 97.455 38.400 ;
        RECT 4.400 37.040 95.600 37.760 ;
        RECT 4.000 36.400 95.600 37.040 ;
        RECT 4.400 36.360 95.600 36.400 ;
        RECT 4.400 35.720 97.455 36.360 ;
        RECT 4.400 35.000 95.600 35.720 ;
        RECT 4.000 34.360 95.600 35.000 ;
        RECT 4.400 34.320 95.600 34.360 ;
        RECT 4.400 33.000 97.455 34.320 ;
        RECT 4.400 32.960 95.600 33.000 ;
        RECT 4.000 32.320 95.600 32.960 ;
        RECT 4.400 31.600 95.600 32.320 ;
        RECT 4.400 30.960 97.455 31.600 ;
        RECT 4.400 30.920 95.600 30.960 ;
        RECT 4.000 30.280 95.600 30.920 ;
        RECT 4.400 29.560 95.600 30.280 ;
        RECT 4.400 28.920 97.455 29.560 ;
        RECT 4.400 28.880 95.600 28.920 ;
        RECT 4.000 28.240 95.600 28.880 ;
        RECT 4.400 27.520 95.600 28.240 ;
        RECT 4.400 26.880 97.455 27.520 ;
        RECT 4.400 26.840 95.600 26.880 ;
        RECT 4.000 26.200 95.600 26.840 ;
        RECT 4.400 25.480 95.600 26.200 ;
        RECT 4.400 24.840 97.455 25.480 ;
        RECT 4.400 24.800 95.600 24.840 ;
        RECT 4.000 24.160 95.600 24.800 ;
        RECT 4.400 23.440 95.600 24.160 ;
        RECT 4.400 22.800 97.455 23.440 ;
        RECT 4.400 22.760 95.600 22.800 ;
        RECT 4.000 22.120 95.600 22.760 ;
        RECT 4.400 21.400 95.600 22.120 ;
        RECT 4.400 20.760 97.455 21.400 ;
        RECT 4.400 20.720 95.600 20.760 ;
        RECT 4.000 20.080 95.600 20.720 ;
        RECT 4.400 19.360 95.600 20.080 ;
        RECT 4.400 18.720 97.455 19.360 ;
        RECT 4.400 18.680 95.600 18.720 ;
        RECT 4.000 18.040 95.600 18.680 ;
        RECT 4.400 17.320 95.600 18.040 ;
        RECT 4.400 16.640 97.455 17.320 ;
        RECT 4.000 16.000 97.455 16.640 ;
        RECT 4.400 14.600 95.600 16.000 ;
        RECT 4.000 13.960 97.455 14.600 ;
        RECT 4.400 12.560 95.600 13.960 ;
        RECT 4.000 11.920 97.455 12.560 ;
        RECT 4.400 10.520 95.600 11.920 ;
        RECT 4.000 9.880 97.455 10.520 ;
        RECT 4.400 8.480 95.600 9.880 ;
        RECT 4.000 7.840 97.455 8.480 ;
        RECT 4.400 6.440 95.600 7.840 ;
        RECT 4.000 5.800 97.455 6.440 ;
        RECT 4.400 4.400 95.600 5.800 ;
        RECT 4.000 3.760 97.455 4.400 ;
        RECT 4.400 2.360 95.600 3.760 ;
        RECT 4.000 1.720 97.455 2.360 ;
        RECT 4.400 0.855 95.600 1.720 ;
      LAYER met4 ;
        RECT 21.545 10.640 33.975 73.680 ;
        RECT 36.375 10.640 81.585 73.680 ;
  END
END cbx_1__2_
END LIBRARY

