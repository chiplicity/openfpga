VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__3_
  CLASS BLOCK ;
  FOREIGN sb_1__3_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 137.600 4.050 140.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 137.600 11.870 140.000 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 137.600 20.150 140.000 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 137.600 28.430 140.000 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.400 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 2.400 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 137.600 36.710 140.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 2.760 140.000 3.360 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 8.200 140.000 8.800 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 14.320 140.000 14.920 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 19.760 140.000 20.360 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 25.880 140.000 26.480 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 31.320 140.000 31.920 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.710 137.600 44.990 140.000 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 2.400 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 2.400 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 37.440 140.000 38.040 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 2.400 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 2.400 34.640 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 43.560 140.000 44.160 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 2.400 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 49.000 140.000 49.600 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 137.600 53.270 140.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 137.600 61.550 140.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.400 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 55.120 140.000 55.720 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 137.600 77.650 140.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 2.400 60.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 60.560 140.000 61.160 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 66.680 140.000 67.280 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.400 66.600 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 72.800 140.000 73.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 137.600 85.930 140.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 137.600 94.210 140.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.400 92.440 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 78.240 140.000 78.840 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 84.360 140.000 84.960 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 2.400 98.560 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 2.400 104.680 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 137.600 102.490 140.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.800 140.000 90.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 2.400 111.480 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 137.600 110.770 140.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.920 140.000 96.520 ;
    END
  END chany_bottom_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 2.400 ;
    END
  END left_top_grid_pin_11_
  PIN left_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 125.160 140.000 125.760 ;
    END
  END left_top_grid_pin_13_
  PIN left_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 2.400 ;
    END
  END left_top_grid_pin_15_
  PIN left_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 107.480 140.000 108.080 ;
    END
  END left_top_grid_pin_1_
  PIN left_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 113.600 140.000 114.200 ;
    END
  END left_top_grid_pin_3_
  PIN left_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 119.040 140.000 119.640 ;
    END
  END left_top_grid_pin_5_
  PIN left_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 137.600 119.050 140.000 ;
    END
  END left_top_grid_pin_7_
  PIN left_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 2.400 ;
    END
  END left_top_grid_pin_9_
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 137.600 127.330 140.000 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.720 140.000 137.320 ;
    END
  END right_top_grid_pin_11_
  PIN right_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 2.400 ;
    END
  END right_top_grid_pin_13_
  PIN right_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 2.400 136.640 ;
    END
  END right_top_grid_pin_15_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 2.400 117.600 ;
    END
  END right_top_grid_pin_1_
  PIN right_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 130.600 140.000 131.200 ;
    END
  END right_top_grid_pin_3_
  PIN right_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 2.400 123.720 ;
    END
  END right_top_grid_pin_5_
  PIN right_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.330 137.600 135.610 140.000 ;
    END
  END right_top_grid_pin_7_
  PIN right_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 2.400 130.520 ;
    END
  END right_top_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.070 0.380 138.390 137.660 ;
      LAYER met2 ;
        RECT 0.090 137.320 3.490 137.770 ;
        RECT 4.330 137.320 11.310 137.770 ;
        RECT 12.150 137.320 19.590 137.770 ;
        RECT 20.430 137.320 27.870 137.770 ;
        RECT 28.710 137.320 36.150 137.770 ;
        RECT 36.990 137.320 44.430 137.770 ;
        RECT 45.270 137.320 52.710 137.770 ;
        RECT 53.550 137.320 60.990 137.770 ;
        RECT 61.830 137.320 69.270 137.770 ;
        RECT 70.110 137.320 77.090 137.770 ;
        RECT 77.930 137.320 85.370 137.770 ;
        RECT 86.210 137.320 93.650 137.770 ;
        RECT 94.490 137.320 101.930 137.770 ;
        RECT 102.770 137.320 110.210 137.770 ;
        RECT 111.050 137.320 118.490 137.770 ;
        RECT 119.330 137.320 126.770 137.770 ;
        RECT 127.610 137.320 135.050 137.770 ;
        RECT 135.890 137.320 138.370 137.770 ;
        RECT 0.090 2.680 138.370 137.320 ;
        RECT 0.090 0.270 3.030 2.680 ;
        RECT 3.870 0.270 9.930 2.680 ;
        RECT 10.770 0.270 16.830 2.680 ;
        RECT 17.670 0.270 23.730 2.680 ;
        RECT 24.570 0.270 30.630 2.680 ;
        RECT 31.470 0.270 37.990 2.680 ;
        RECT 38.830 0.270 44.890 2.680 ;
        RECT 45.730 0.270 51.790 2.680 ;
        RECT 52.630 0.270 58.690 2.680 ;
        RECT 59.530 0.270 65.590 2.680 ;
        RECT 66.430 0.270 72.950 2.680 ;
        RECT 73.790 0.270 79.850 2.680 ;
        RECT 80.690 0.270 86.750 2.680 ;
        RECT 87.590 0.270 93.650 2.680 ;
        RECT 94.490 0.270 100.550 2.680 ;
        RECT 101.390 0.270 107.910 2.680 ;
        RECT 108.750 0.270 114.810 2.680 ;
        RECT 115.650 0.270 121.710 2.680 ;
        RECT 122.550 0.270 128.610 2.680 ;
        RECT 129.450 0.270 135.510 2.680 ;
        RECT 136.350 0.270 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 136.320 137.200 136.720 ;
        RECT 2.800 135.640 138.650 136.320 ;
        RECT 0.270 131.600 138.650 135.640 ;
        RECT 0.270 130.920 137.200 131.600 ;
        RECT 2.800 130.200 137.200 130.920 ;
        RECT 2.800 129.520 138.650 130.200 ;
        RECT 0.270 126.160 138.650 129.520 ;
        RECT 0.270 124.760 137.200 126.160 ;
        RECT 0.270 124.120 138.650 124.760 ;
        RECT 2.800 122.720 138.650 124.120 ;
        RECT 0.270 120.040 138.650 122.720 ;
        RECT 0.270 118.640 137.200 120.040 ;
        RECT 0.270 118.000 138.650 118.640 ;
        RECT 2.800 116.600 138.650 118.000 ;
        RECT 0.270 114.600 138.650 116.600 ;
        RECT 0.270 113.200 137.200 114.600 ;
        RECT 0.270 111.880 138.650 113.200 ;
        RECT 2.800 110.480 138.650 111.880 ;
        RECT 0.270 108.480 138.650 110.480 ;
        RECT 0.270 107.080 137.200 108.480 ;
        RECT 0.270 105.080 138.650 107.080 ;
        RECT 2.800 103.680 138.650 105.080 ;
        RECT 0.270 102.360 138.650 103.680 ;
        RECT 0.270 100.960 137.200 102.360 ;
        RECT 0.270 98.960 138.650 100.960 ;
        RECT 2.800 97.560 138.650 98.960 ;
        RECT 0.270 96.920 138.650 97.560 ;
        RECT 0.270 95.520 137.200 96.920 ;
        RECT 0.270 92.840 138.650 95.520 ;
        RECT 2.800 91.440 138.650 92.840 ;
        RECT 0.270 90.800 138.650 91.440 ;
        RECT 0.270 89.400 137.200 90.800 ;
        RECT 0.270 86.040 138.650 89.400 ;
        RECT 2.800 85.360 138.650 86.040 ;
        RECT 2.800 84.640 137.200 85.360 ;
        RECT 0.270 83.960 137.200 84.640 ;
        RECT 0.270 79.920 138.650 83.960 ;
        RECT 2.800 79.240 138.650 79.920 ;
        RECT 2.800 78.520 137.200 79.240 ;
        RECT 0.270 77.840 137.200 78.520 ;
        RECT 0.270 73.800 138.650 77.840 ;
        RECT 2.800 72.400 137.200 73.800 ;
        RECT 0.270 67.680 138.650 72.400 ;
        RECT 0.270 67.000 137.200 67.680 ;
        RECT 2.800 66.280 137.200 67.000 ;
        RECT 2.800 65.600 138.650 66.280 ;
        RECT 0.270 61.560 138.650 65.600 ;
        RECT 0.270 60.880 137.200 61.560 ;
        RECT 2.800 60.160 137.200 60.880 ;
        RECT 2.800 59.480 138.650 60.160 ;
        RECT 0.270 56.120 138.650 59.480 ;
        RECT 0.270 54.720 137.200 56.120 ;
        RECT 0.270 54.080 138.650 54.720 ;
        RECT 2.800 52.680 138.650 54.080 ;
        RECT 0.270 50.000 138.650 52.680 ;
        RECT 0.270 48.600 137.200 50.000 ;
        RECT 0.270 47.960 138.650 48.600 ;
        RECT 2.800 46.560 138.650 47.960 ;
        RECT 0.270 44.560 138.650 46.560 ;
        RECT 0.270 43.160 137.200 44.560 ;
        RECT 0.270 41.840 138.650 43.160 ;
        RECT 2.800 40.440 138.650 41.840 ;
        RECT 0.270 38.440 138.650 40.440 ;
        RECT 0.270 37.040 137.200 38.440 ;
        RECT 0.270 35.040 138.650 37.040 ;
        RECT 2.800 33.640 138.650 35.040 ;
        RECT 0.270 32.320 138.650 33.640 ;
        RECT 0.270 30.920 137.200 32.320 ;
        RECT 0.270 28.920 138.650 30.920 ;
        RECT 2.800 27.520 138.650 28.920 ;
        RECT 0.270 26.880 138.650 27.520 ;
        RECT 0.270 25.480 137.200 26.880 ;
        RECT 0.270 22.800 138.650 25.480 ;
        RECT 2.800 21.400 138.650 22.800 ;
        RECT 0.270 20.760 138.650 21.400 ;
        RECT 0.270 19.360 137.200 20.760 ;
        RECT 0.270 16.000 138.650 19.360 ;
        RECT 2.800 15.320 138.650 16.000 ;
        RECT 2.800 14.600 137.200 15.320 ;
        RECT 0.270 13.920 137.200 14.600 ;
        RECT 0.270 9.880 138.650 13.920 ;
        RECT 2.800 9.200 138.650 9.880 ;
        RECT 2.800 8.480 137.200 9.200 ;
        RECT 0.270 7.800 137.200 8.480 ;
        RECT 0.270 3.760 138.650 7.800 ;
        RECT 2.800 3.360 137.200 3.760 ;
      LAYER met4 ;
        RECT 0.295 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 138.625 128.080 ;
  END
END sb_1__3_
END LIBRARY

