magic
tech EFS8A
magscale 1 2
timestamp 1604337187
<< locali >>
rect 7665 25687 7699 25993
rect 12081 25755 12115 26605
rect 12173 25823 12207 26401
rect 12449 26367 12483 26741
rect 12449 25823 12483 26197
rect 19901 26027 19935 26197
rect 19993 25959 20027 26197
rect 17785 25823 17819 25925
rect 7665 24667 7699 24837
rect 12081 23511 12115 23681
rect 22569 23511 22603 23817
rect 11621 22423 11655 22729
rect 17233 22423 17267 22593
rect 20269 22423 20303 22525
rect 19901 21879 19935 21981
rect 10057 21335 10091 21437
rect 11621 21403 11655 21641
rect 17601 21403 17635 21641
rect 2881 20247 2915 20553
rect 19901 19703 19935 20009
rect 4537 19159 4571 19261
rect 6101 18615 6135 18921
rect 11989 18071 12023 18241
rect 22201 18071 22235 18377
rect 8309 17595 8343 17765
rect 12081 16983 12115 17153
rect 15209 14807 15243 15113
rect 6009 12699 6043 12937
rect 19717 12767 19751 12937
rect 5549 12087 5583 12189
rect 9321 12087 9355 12393
rect 6377 11543 6411 11849
rect 10333 11543 10367 11781
rect 22661 9911 22695 10217
rect 6377 9367 6411 9469
rect 22109 9367 22143 9469
rect 24501 9367 24535 9673
rect 21833 8823 21867 9129
rect 11161 8279 11195 8449
rect 20821 8347 20855 8517
rect 20269 3927 20303 4097
rect 3249 3519 3283 3621
rect 10793 3451 10827 3553
rect 12081 2839 12115 2941
<< viali >>
rect 12449 26741 12483 26775
rect 12081 26605 12115 26639
rect 7665 25993 7699 26027
rect 12173 26401 12207 26435
rect 12449 26333 12483 26367
rect 12173 25789 12207 25823
rect 12449 26197 12483 26231
rect 19901 26197 19935 26231
rect 19901 25993 19935 26027
rect 19993 26197 20027 26231
rect 12449 25789 12483 25823
rect 17785 25925 17819 25959
rect 19993 25925 20027 25959
rect 17785 25789 17819 25823
rect 12081 25721 12115 25755
rect 7665 25653 7699 25687
rect 7665 25449 7699 25483
rect 8769 25449 8803 25483
rect 10057 25449 10091 25483
rect 11529 25449 11563 25483
rect 14473 25449 14507 25483
rect 14933 25449 14967 25483
rect 19717 25449 19751 25483
rect 21925 25449 21959 25483
rect 12449 25381 12483 25415
rect 13185 25381 13219 25415
rect 15853 25381 15887 25415
rect 16037 25381 16071 25415
rect 7481 25313 7515 25347
rect 8585 25313 8619 25347
rect 9873 25313 9907 25347
rect 11345 25313 11379 25347
rect 13001 25313 13035 25347
rect 14289 25313 14323 25347
rect 17141 25313 17175 25347
rect 18429 25313 18463 25347
rect 19533 25313 19567 25347
rect 21741 25313 21775 25347
rect 22845 25313 22879 25347
rect 24593 25313 24627 25347
rect 9597 25245 9631 25279
rect 10517 25245 10551 25279
rect 10885 25245 10919 25279
rect 11621 25245 11655 25279
rect 13277 25245 13311 25279
rect 15301 25245 15335 25279
rect 16129 25245 16163 25279
rect 13737 25177 13771 25211
rect 15577 25177 15611 25211
rect 17325 25177 17359 25211
rect 18613 25177 18647 25211
rect 23029 25177 23063 25211
rect 6653 25109 6687 25143
rect 7389 25109 7423 25143
rect 8033 25109 8067 25143
rect 8401 25109 8435 25143
rect 9229 25109 9263 25143
rect 11069 25109 11103 25143
rect 11989 25109 12023 25143
rect 12725 25109 12759 25143
rect 14013 25109 14047 25143
rect 17877 25109 17911 25143
rect 20085 25109 20119 25143
rect 20545 25109 20579 25143
rect 21465 25109 21499 25143
rect 22293 25109 22327 25143
rect 23673 25109 23707 25143
rect 24777 25109 24811 25143
rect 11437 24905 11471 24939
rect 17509 24905 17543 24939
rect 7389 24837 7423 24871
rect 7665 24837 7699 24871
rect 11069 24837 11103 24871
rect 12265 24837 12299 24871
rect 6653 24701 6687 24735
rect 6837 24701 6871 24735
rect 7757 24769 7791 24803
rect 8401 24769 8435 24803
rect 13001 24769 13035 24803
rect 15209 24769 15243 24803
rect 20453 24769 20487 24803
rect 22201 24769 22235 24803
rect 22661 24769 22695 24803
rect 9413 24701 9447 24735
rect 11253 24701 11287 24735
rect 14013 24701 14047 24735
rect 15761 24701 15795 24735
rect 16405 24701 16439 24735
rect 18889 24701 18923 24735
rect 19441 24701 19475 24735
rect 25237 24701 25271 24735
rect 25789 24701 25823 24735
rect 6285 24633 6319 24667
rect 7665 24633 7699 24667
rect 8493 24633 8527 24667
rect 8585 24633 8619 24667
rect 9873 24633 9907 24667
rect 10149 24633 10183 24667
rect 13001 24633 13035 24667
rect 13093 24633 13127 24667
rect 13829 24633 13863 24667
rect 14289 24633 14323 24667
rect 15945 24633 15979 24667
rect 16037 24633 16071 24667
rect 16773 24633 16807 24667
rect 16957 24633 16991 24667
rect 20637 24633 20671 24667
rect 21189 24633 21223 24667
rect 21723 24633 21757 24667
rect 22293 24633 22327 24667
rect 24041 24633 24075 24667
rect 24317 24633 24351 24667
rect 4813 24565 4847 24599
rect 5273 24565 5307 24599
rect 5549 24565 5583 24599
rect 7021 24565 7055 24599
rect 8015 24565 8049 24599
rect 9045 24565 9079 24599
rect 9587 24565 9621 24599
rect 10057 24565 10091 24599
rect 10609 24565 10643 24599
rect 11805 24565 11839 24599
rect 12531 24565 12565 24599
rect 13461 24565 13495 24599
rect 14749 24565 14783 24599
rect 15475 24565 15509 24599
rect 17785 24565 17819 24599
rect 18521 24565 18555 24599
rect 19073 24565 19107 24599
rect 19809 24565 19843 24599
rect 20075 24565 20109 24599
rect 20545 24565 20579 24599
rect 21465 24565 21499 24599
rect 22201 24565 22235 24599
rect 23029 24565 23063 24599
rect 23489 24565 23523 24599
rect 23755 24565 23789 24599
rect 24225 24565 24259 24599
rect 24685 24565 24719 24599
rect 25421 24565 25455 24599
rect 1593 24361 1627 24395
rect 6009 24361 6043 24395
rect 6469 24361 6503 24395
rect 7113 24361 7147 24395
rect 10517 24361 10551 24395
rect 14933 24361 14967 24395
rect 15485 24361 15519 24395
rect 15853 24361 15887 24395
rect 18797 24361 18831 24395
rect 19901 24361 19935 24395
rect 20269 24361 20303 24395
rect 22937 24361 22971 24395
rect 8585 24293 8619 24327
rect 13737 24293 13771 24327
rect 16773 24293 16807 24327
rect 17233 24293 17267 24327
rect 18337 24293 18371 24327
rect 22017 24293 22051 24327
rect 23673 24293 23707 24327
rect 1409 24225 1443 24259
rect 5825 24225 5859 24259
rect 6929 24225 6963 24259
rect 7941 24225 7975 24259
rect 8401 24225 8435 24259
rect 10876 24225 10910 24259
rect 13553 24225 13587 24259
rect 14565 24225 14599 24259
rect 16865 24225 16899 24259
rect 19717 24225 19751 24259
rect 23765 24225 23799 24259
rect 24501 24225 24535 24259
rect 24685 24225 24719 24259
rect 4537 24157 4571 24191
rect 5273 24157 5307 24191
rect 8677 24157 8711 24191
rect 10609 24157 10643 24191
rect 13829 24157 13863 24191
rect 16681 24157 16715 24191
rect 18245 24157 18279 24191
rect 18429 24157 18463 24191
rect 21925 24157 21959 24191
rect 22109 24157 22143 24191
rect 23581 24157 23615 24191
rect 4905 24089 4939 24123
rect 8125 24089 8159 24123
rect 12725 24089 12759 24123
rect 13277 24089 13311 24123
rect 14289 24089 14323 24123
rect 21373 24089 21407 24123
rect 5733 24021 5767 24055
rect 6837 24021 6871 24055
rect 7573 24021 7607 24055
rect 9137 24021 9171 24055
rect 9505 24021 9539 24055
rect 9873 24021 9907 24055
rect 11989 24021 12023 24055
rect 13093 24021 13127 24055
rect 16313 24021 16347 24055
rect 17601 24021 17635 24055
rect 17877 24021 17911 24055
rect 19165 24021 19199 24055
rect 19533 24021 19567 24055
rect 20729 24021 20763 24055
rect 21557 24021 21591 24055
rect 22569 24021 22603 24055
rect 23213 24021 23247 24055
rect 24133 24021 24167 24055
rect 24869 24021 24903 24055
rect 1593 23817 1627 23851
rect 5825 23817 5859 23851
rect 7573 23817 7607 23851
rect 12541 23817 12575 23851
rect 15577 23817 15611 23851
rect 18153 23817 18187 23851
rect 19165 23817 19199 23851
rect 19625 23817 19659 23851
rect 21189 23817 21223 23851
rect 22569 23817 22603 23851
rect 22845 23817 22879 23851
rect 25697 23817 25731 23851
rect 11437 23749 11471 23783
rect 19809 23749 19843 23783
rect 21373 23749 21407 23783
rect 7389 23681 7423 23715
rect 8033 23681 8067 23715
rect 12081 23681 12115 23715
rect 13093 23681 13127 23715
rect 17509 23681 17543 23715
rect 18705 23681 18739 23715
rect 21925 23681 21959 23715
rect 1409 23613 1443 23647
rect 5089 23613 5123 23647
rect 5641 23613 5675 23647
rect 9045 23613 9079 23647
rect 9301 23613 9335 23647
rect 11069 23613 11103 23647
rect 3617 23545 3651 23579
rect 4353 23545 4387 23579
rect 5549 23545 5583 23579
rect 6653 23545 6687 23579
rect 8125 23545 8159 23579
rect 11897 23545 11931 23579
rect 12817 23613 12851 23647
rect 13461 23613 13495 23647
rect 14197 23613 14231 23647
rect 16681 23613 16715 23647
rect 20085 23613 20119 23647
rect 21649 23613 21683 23647
rect 13001 23545 13035 23579
rect 14464 23545 14498 23579
rect 16957 23545 16991 23579
rect 18429 23545 18463 23579
rect 18613 23545 18647 23579
rect 20361 23545 20395 23579
rect 21833 23545 21867 23579
rect 24041 23749 24075 23783
rect 24593 23681 24627 23715
rect 25513 23613 25547 23647
rect 26065 23613 26099 23647
rect 23121 23545 23155 23579
rect 24317 23545 24351 23579
rect 2053 23477 2087 23511
rect 2421 23477 2455 23511
rect 3249 23477 3283 23511
rect 3893 23477 3927 23511
rect 4721 23477 4755 23511
rect 6193 23477 6227 23511
rect 8033 23477 8067 23511
rect 8493 23477 8527 23511
rect 8861 23477 8895 23511
rect 10425 23477 10459 23511
rect 12081 23477 12115 23511
rect 12173 23477 12207 23511
rect 14013 23477 14047 23511
rect 16221 23477 16255 23511
rect 17877 23477 17911 23511
rect 20269 23477 20303 23511
rect 20821 23477 20855 23511
rect 22385 23477 22419 23511
rect 22569 23477 22603 23511
rect 24501 23477 24535 23511
rect 24961 23477 24995 23511
rect 1593 23273 1627 23307
rect 5549 23273 5583 23307
rect 11069 23273 11103 23307
rect 12817 23273 12851 23307
rect 13277 23273 13311 23307
rect 16405 23273 16439 23307
rect 18153 23273 18187 23307
rect 20177 23273 20211 23307
rect 21465 23273 21499 23307
rect 21925 23273 21959 23307
rect 22835 23273 22869 23307
rect 24869 23273 24903 23307
rect 25329 23273 25363 23307
rect 7021 23205 7055 23239
rect 8401 23205 8435 23239
rect 8585 23205 8619 23239
rect 8677 23205 8711 23239
rect 15669 23205 15703 23239
rect 15853 23205 15887 23239
rect 17417 23205 17451 23239
rect 18797 23205 18831 23239
rect 18981 23205 19015 23239
rect 23305 23205 23339 23239
rect 24685 23205 24719 23239
rect 1409 23137 1443 23171
rect 2513 23137 2547 23171
rect 5365 23137 5399 23171
rect 7113 23137 7147 23171
rect 9956 23137 9990 23171
rect 12633 23137 12667 23171
rect 13921 23137 13955 23171
rect 17509 23137 17543 23171
rect 23397 23137 23431 23171
rect 4537 23069 4571 23103
rect 7021 23069 7055 23103
rect 9137 23069 9171 23103
rect 9689 23069 9723 23103
rect 12909 23069 12943 23103
rect 14105 23069 14139 23103
rect 15945 23069 15979 23103
rect 17417 23069 17451 23103
rect 19073 23069 19107 23103
rect 21373 23069 21407 23103
rect 21557 23069 21591 23103
rect 23305 23069 23339 23103
rect 24961 23069 24995 23103
rect 3433 23001 3467 23035
rect 6377 23001 6411 23035
rect 7849 23001 7883 23035
rect 8125 23001 8159 23035
rect 12357 23001 12391 23035
rect 15117 23001 15151 23035
rect 15393 23001 15427 23035
rect 16957 23001 16991 23035
rect 21005 23001 21039 23035
rect 25697 23001 25731 23035
rect 1961 22933 1995 22967
rect 2329 22933 2363 22967
rect 2697 22933 2731 22967
rect 3065 22933 3099 22967
rect 3801 22933 3835 22967
rect 4813 22933 4847 22967
rect 5273 22933 5307 22967
rect 6009 22933 6043 22967
rect 6561 22933 6595 22967
rect 7573 22933 7607 22967
rect 9505 22933 9539 22967
rect 11621 22933 11655 22967
rect 11989 22933 12023 22967
rect 13737 22933 13771 22967
rect 14657 22933 14691 22967
rect 16681 22933 16715 22967
rect 18521 22933 18555 22967
rect 19717 22933 19751 22967
rect 20545 22933 20579 22967
rect 22569 22933 22603 22967
rect 23949 22933 23983 22967
rect 24409 22933 24443 22967
rect 2697 22729 2731 22763
rect 7389 22729 7423 22763
rect 7757 22729 7791 22763
rect 9321 22729 9355 22763
rect 10885 22729 10919 22763
rect 11621 22729 11655 22763
rect 14749 22729 14783 22763
rect 15669 22729 15703 22763
rect 16497 22729 16531 22763
rect 17417 22729 17451 22763
rect 20085 22729 20119 22763
rect 23397 22729 23431 22763
rect 1593 22661 1627 22695
rect 5273 22661 5307 22695
rect 8769 22661 8803 22695
rect 2421 22593 2455 22627
rect 4721 22593 4755 22627
rect 5733 22593 5767 22627
rect 8125 22593 8159 22627
rect 9781 22593 9815 22627
rect 11253 22593 11287 22627
rect 11437 22593 11471 22627
rect 1409 22525 1443 22559
rect 2513 22525 2547 22559
rect 3617 22525 3651 22559
rect 5825 22525 5859 22559
rect 8309 22525 8343 22559
rect 9045 22525 9079 22559
rect 9873 22525 9907 22559
rect 10609 22525 10643 22559
rect 3433 22457 3467 22491
rect 4353 22457 4387 22491
rect 9781 22457 9815 22491
rect 10333 22457 10367 22491
rect 16313 22661 16347 22695
rect 20637 22661 20671 22695
rect 23765 22661 23799 22695
rect 17049 22593 17083 22627
rect 17233 22593 17267 22627
rect 20453 22593 20487 22627
rect 21097 22593 21131 22627
rect 22385 22593 22419 22627
rect 25421 22593 25455 22627
rect 12173 22525 12207 22559
rect 13369 22525 13403 22559
rect 12725 22457 12759 22491
rect 13636 22457 13670 22491
rect 16773 22457 16807 22491
rect 16957 22457 16991 22491
rect 17785 22525 17819 22559
rect 18061 22525 18095 22559
rect 20269 22525 20303 22559
rect 21189 22525 21223 22559
rect 22109 22525 22143 22559
rect 24685 22525 24719 22559
rect 25237 22525 25271 22559
rect 25973 22525 26007 22559
rect 18306 22457 18340 22491
rect 21557 22457 21591 22491
rect 24041 22457 24075 22491
rect 24317 22457 24351 22491
rect 1961 22389 1995 22423
rect 3065 22389 3099 22423
rect 3801 22389 3835 22423
rect 5089 22389 5123 22423
rect 5733 22389 5767 22423
rect 6561 22389 6595 22423
rect 7113 22389 7147 22423
rect 8217 22389 8251 22423
rect 11345 22389 11379 22423
rect 11621 22389 11655 22423
rect 11897 22389 11931 22423
rect 13185 22389 13219 22423
rect 15301 22389 15335 22423
rect 17233 22389 17267 22423
rect 19441 22389 19475 22423
rect 20269 22389 20303 22423
rect 21097 22389 21131 22423
rect 22017 22389 22051 22423
rect 23121 22389 23155 22423
rect 24225 22389 24259 22423
rect 25053 22389 25087 22423
rect 1961 22185 1995 22219
rect 5457 22185 5491 22219
rect 6551 22185 6585 22219
rect 16497 22185 16531 22219
rect 17969 22185 18003 22219
rect 21465 22185 21499 22219
rect 24593 22185 24627 22219
rect 7021 22117 7055 22151
rect 8585 22117 8619 22151
rect 10241 22117 10275 22151
rect 11253 22117 11287 22151
rect 12173 22117 12207 22151
rect 13691 22117 13725 22151
rect 18889 22117 18923 22151
rect 19625 22117 19659 22151
rect 20987 22117 21021 22151
rect 21281 22117 21315 22151
rect 22385 22117 22419 22151
rect 23029 22117 23063 22151
rect 1409 22049 1443 22083
rect 2513 22049 2547 22083
rect 6377 22049 6411 22083
rect 7113 22049 7147 22083
rect 7757 22049 7791 22083
rect 8401 22049 8435 22083
rect 10333 22049 10367 22083
rect 11989 22049 12023 22083
rect 15301 22049 15335 22083
rect 15577 22049 15611 22083
rect 16856 22049 16890 22083
rect 18613 22049 18647 22083
rect 20637 22049 20671 22083
rect 24409 22049 24443 22083
rect 25053 22049 25087 22083
rect 5365 21981 5399 22015
rect 5549 21981 5583 22015
rect 7021 21981 7055 22015
rect 8677 21981 8711 22015
rect 9137 21981 9171 22015
rect 10241 21981 10275 22015
rect 12265 21981 12299 22015
rect 13093 21981 13127 22015
rect 13737 21981 13771 22015
rect 13829 21981 13863 22015
rect 15117 21981 15151 22015
rect 16589 21981 16623 22015
rect 19533 21981 19567 22015
rect 19717 21981 19751 22015
rect 19901 21981 19935 22015
rect 21557 21981 21591 22015
rect 23029 21981 23063 22015
rect 23121 21981 23155 22015
rect 24685 21981 24719 22015
rect 25421 21981 25455 22015
rect 2697 21913 2731 21947
rect 4997 21913 5031 21947
rect 9781 21913 9815 21947
rect 13277 21913 13311 21947
rect 14749 21913 14783 21947
rect 19165 21913 19199 21947
rect 22569 21913 22603 21947
rect 24133 21913 24167 21947
rect 1593 21845 1627 21879
rect 2421 21845 2455 21879
rect 3065 21845 3099 21879
rect 3617 21845 3651 21879
rect 4261 21845 4295 21879
rect 4629 21845 4663 21879
rect 6009 21845 6043 21879
rect 8125 21845 8159 21879
rect 9413 21845 9447 21879
rect 10793 21845 10827 21879
rect 11713 21845 11747 21879
rect 12725 21845 12759 21879
rect 14289 21845 14323 21879
rect 16037 21845 16071 21879
rect 19901 21845 19935 21879
rect 20177 21845 20211 21879
rect 21925 21845 21959 21879
rect 23673 21845 23707 21879
rect 25789 21845 25823 21879
rect 2973 21641 3007 21675
rect 5273 21641 5307 21675
rect 10885 21641 10919 21675
rect 11621 21641 11655 21675
rect 13829 21641 13863 21675
rect 15209 21641 15243 21675
rect 15485 21641 15519 21675
rect 16497 21641 16531 21675
rect 17601 21641 17635 21675
rect 18245 21641 18279 21675
rect 22569 21641 22603 21675
rect 23765 21641 23799 21675
rect 26341 21641 26375 21675
rect 3709 21573 3743 21607
rect 4997 21573 5031 21607
rect 2053 21505 2087 21539
rect 11345 21505 11379 21539
rect 1777 21437 1811 21471
rect 3525 21437 3559 21471
rect 6929 21437 6963 21471
rect 8217 21437 8251 21471
rect 8473 21437 8507 21471
rect 10057 21437 10091 21471
rect 3985 21369 4019 21403
rect 4261 21369 4295 21403
rect 5549 21369 5583 21403
rect 5825 21369 5859 21403
rect 6469 21369 6503 21403
rect 7205 21369 7239 21403
rect 7757 21369 7791 21403
rect 14473 21505 14507 21539
rect 16865 21505 16899 21539
rect 12173 21437 12207 21471
rect 12449 21437 12483 21471
rect 12716 21437 12750 21471
rect 14841 21437 14875 21471
rect 15301 21437 15335 21471
rect 16313 21437 16347 21471
rect 17049 21437 17083 21471
rect 21373 21573 21407 21607
rect 21833 21505 21867 21539
rect 23397 21505 23431 21539
rect 24225 21505 24259 21539
rect 17877 21437 17911 21471
rect 18797 21437 18831 21471
rect 19053 21437 19087 21471
rect 21925 21437 21959 21471
rect 24685 21437 24719 21471
rect 25237 21437 25271 21471
rect 10517 21369 10551 21403
rect 11345 21369 11379 21403
rect 11437 21369 11471 21403
rect 11621 21369 11655 21403
rect 17417 21369 17451 21403
rect 17601 21369 17635 21403
rect 18705 21369 18739 21403
rect 24317 21369 24351 21403
rect 25513 21369 25547 21403
rect 1685 21301 1719 21335
rect 2605 21301 2639 21335
rect 4169 21301 4203 21335
rect 5733 21301 5767 21335
rect 8033 21301 8067 21335
rect 9597 21301 9631 21335
rect 10057 21301 10091 21335
rect 10149 21301 10183 21335
rect 11897 21301 11931 21335
rect 15945 21301 15979 21335
rect 16957 21301 16991 21335
rect 20177 21301 20211 21335
rect 21005 21301 21039 21335
rect 21833 21301 21867 21335
rect 23121 21301 23155 21335
rect 24225 21301 24259 21335
rect 25145 21301 25179 21335
rect 25973 21301 26007 21335
rect 2973 21097 3007 21131
rect 5641 21097 5675 21131
rect 6561 21097 6595 21131
rect 8033 21097 8067 21131
rect 8953 21097 8987 21131
rect 9505 21097 9539 21131
rect 11069 21097 11103 21131
rect 12081 21097 12115 21131
rect 13921 21097 13955 21131
rect 14289 21097 14323 21131
rect 15025 21097 15059 21131
rect 15853 21097 15887 21131
rect 16497 21097 16531 21131
rect 19533 21097 19567 21131
rect 21465 21097 21499 21131
rect 25421 21097 25455 21131
rect 26157 21097 26191 21131
rect 2789 21029 2823 21063
rect 3065 21029 3099 21063
rect 8585 21029 8619 21063
rect 9934 21029 9968 21063
rect 13093 21029 13127 21063
rect 15669 21029 15703 21063
rect 17233 21029 17267 21063
rect 17371 21029 17405 21063
rect 17509 21029 17543 21063
rect 18981 21029 19015 21063
rect 20085 21029 20119 21063
rect 21557 21029 21591 21063
rect 23029 21029 23063 21063
rect 24593 21029 24627 21063
rect 25053 21029 25087 21063
rect 3709 20961 3743 20995
rect 6193 20961 6227 20995
rect 6920 20961 6954 20995
rect 12909 20961 12943 20995
rect 14105 20961 14139 20995
rect 18797 20961 18831 20995
rect 22845 20961 22879 20995
rect 4077 20893 4111 20927
rect 5549 20893 5583 20927
rect 5733 20893 5767 20927
rect 6653 20893 6687 20927
rect 9689 20893 9723 20927
rect 11713 20893 11747 20927
rect 13185 20893 13219 20927
rect 15945 20893 15979 20927
rect 19073 20893 19107 20927
rect 21373 20893 21407 20927
rect 23121 20893 23155 20927
rect 24593 20893 24627 20927
rect 24685 20893 24719 20927
rect 25789 20893 25823 20927
rect 5181 20825 5215 20859
rect 12449 20825 12483 20859
rect 15393 20825 15427 20859
rect 16957 20825 16991 20859
rect 18153 20825 18187 20859
rect 21005 20825 21039 20859
rect 22569 20825 22603 20859
rect 24133 20825 24167 20859
rect 1777 20757 1811 20791
rect 2053 20757 2087 20791
rect 2513 20757 2547 20791
rect 4537 20757 4571 20791
rect 4997 20757 5031 20791
rect 12633 20757 12667 20791
rect 13645 20757 13679 20791
rect 18521 20757 18555 20791
rect 20361 20757 20395 20791
rect 22017 20757 22051 20791
rect 22385 20757 22419 20791
rect 23673 20757 23707 20791
rect 2881 20553 2915 20587
rect 3433 20553 3467 20587
rect 3709 20553 3743 20587
rect 4721 20553 4755 20587
rect 7573 20553 7607 20587
rect 9321 20553 9355 20587
rect 10885 20553 10919 20587
rect 12265 20553 12299 20587
rect 14841 20553 14875 20587
rect 15945 20553 15979 20587
rect 16773 20553 16807 20587
rect 17049 20553 17083 20587
rect 17877 20553 17911 20587
rect 18521 20553 18555 20587
rect 20453 20553 20487 20587
rect 22017 20553 22051 20587
rect 23765 20553 23799 20587
rect 2145 20485 2179 20519
rect 2697 20417 2731 20451
rect 1961 20281 1995 20315
rect 2421 20281 2455 20315
rect 5273 20485 5307 20519
rect 10333 20485 10367 20519
rect 15025 20485 15059 20519
rect 17417 20485 17451 20519
rect 18889 20485 18923 20519
rect 21741 20485 21775 20519
rect 4261 20417 4295 20451
rect 5825 20417 5859 20451
rect 8125 20417 8159 20451
rect 8309 20417 8343 20451
rect 9781 20417 9815 20451
rect 11345 20417 11379 20451
rect 15393 20417 15427 20451
rect 19257 20417 19291 20451
rect 20269 20417 20303 20451
rect 20913 20417 20947 20451
rect 22569 20417 22603 20451
rect 3985 20349 4019 20383
rect 5549 20349 5583 20383
rect 7739 20349 7773 20383
rect 9137 20349 9171 20383
rect 9873 20349 9907 20383
rect 10701 20349 10735 20383
rect 11437 20349 11471 20383
rect 11805 20349 11839 20383
rect 12449 20349 12483 20383
rect 12705 20349 12739 20383
rect 16871 20349 16905 20383
rect 21005 20349 21039 20383
rect 25237 20349 25271 20383
rect 25973 20349 26007 20383
rect 6561 20281 6595 20315
rect 9781 20281 9815 20315
rect 11345 20281 11379 20315
rect 15485 20281 15519 20315
rect 15577 20281 15611 20315
rect 19441 20281 19475 20315
rect 22293 20281 22327 20315
rect 22477 20281 22511 20315
rect 23121 20281 23155 20315
rect 24041 20281 24075 20315
rect 24317 20281 24351 20315
rect 25513 20281 25547 20315
rect 2605 20213 2639 20247
rect 2881 20213 2915 20247
rect 3157 20213 3191 20247
rect 4169 20213 4203 20247
rect 4997 20213 5031 20247
rect 5733 20213 5767 20247
rect 6285 20213 6319 20247
rect 7205 20213 7239 20247
rect 8217 20213 8251 20247
rect 8677 20213 8711 20247
rect 13829 20213 13863 20247
rect 14381 20213 14415 20247
rect 16405 20213 16439 20247
rect 19349 20213 19383 20247
rect 19809 20213 19843 20247
rect 20913 20213 20947 20247
rect 21373 20213 21407 20247
rect 23489 20213 23523 20247
rect 24225 20213 24259 20247
rect 24685 20213 24719 20247
rect 25053 20213 25087 20247
rect 26341 20213 26375 20247
rect 1777 20009 1811 20043
rect 2145 20009 2179 20043
rect 2973 20009 3007 20043
rect 4905 20009 4939 20043
rect 7297 20009 7331 20043
rect 7941 20009 7975 20043
rect 8309 20009 8343 20043
rect 9505 20009 9539 20043
rect 13645 20009 13679 20043
rect 14197 20009 14231 20043
rect 14657 20009 14691 20043
rect 15025 20009 15059 20043
rect 15761 20009 15795 20043
rect 17693 20009 17727 20043
rect 18889 20009 18923 20043
rect 19533 20009 19567 20043
rect 19901 20009 19935 20043
rect 25421 20009 25455 20043
rect 4721 19941 4755 19975
rect 5825 19941 5859 19975
rect 10241 19941 10275 19975
rect 12081 19941 12115 19975
rect 15301 19941 15335 19975
rect 16558 19941 16592 19975
rect 19625 19941 19659 19975
rect 2789 19873 2823 19907
rect 3709 19873 3743 19907
rect 5457 19873 5491 19907
rect 5917 19873 5951 19907
rect 6184 19873 6218 19907
rect 9137 19873 9171 19907
rect 10057 19873 10091 19907
rect 11437 19873 11471 19907
rect 12173 19873 12207 19907
rect 13001 19873 13035 19907
rect 13737 19873 13771 19907
rect 3065 19805 3099 19839
rect 4997 19805 5031 19839
rect 8585 19805 8619 19839
rect 10333 19805 10367 19839
rect 11989 19805 12023 19839
rect 13645 19805 13679 19839
rect 16313 19805 16347 19839
rect 19533 19805 19567 19839
rect 2513 19737 2547 19771
rect 4445 19737 4479 19771
rect 12633 19737 12667 19771
rect 19073 19737 19107 19771
rect 20085 19941 20119 19975
rect 23397 19941 23431 19975
rect 24409 19941 24443 19975
rect 20453 19873 20487 19907
rect 21373 19873 21407 19907
rect 21640 19873 21674 19907
rect 25881 19873 25915 19907
rect 23673 19805 23707 19839
rect 24409 19805 24443 19839
rect 24501 19805 24535 19839
rect 25237 19737 25271 19771
rect 9781 19669 9815 19703
rect 10793 19669 10827 19703
rect 11621 19669 11655 19703
rect 13185 19669 13219 19703
rect 16129 19669 16163 19703
rect 18337 19669 18371 19703
rect 19901 19669 19935 19703
rect 21097 19669 21131 19703
rect 22753 19669 22787 19703
rect 23949 19669 23983 19703
rect 24961 19669 24995 19703
rect 3709 19465 3743 19499
rect 5273 19465 5307 19499
rect 7021 19465 7055 19499
rect 10609 19465 10643 19499
rect 13461 19465 13495 19499
rect 16221 19465 16255 19499
rect 19625 19465 19659 19499
rect 20637 19465 20671 19499
rect 22109 19465 22143 19499
rect 23765 19465 23799 19499
rect 23121 19397 23155 19431
rect 4261 19329 4295 19363
rect 5825 19329 5859 19363
rect 6285 19329 6319 19363
rect 16589 19329 16623 19363
rect 20729 19329 20763 19363
rect 2421 19261 2455 19295
rect 3433 19261 3467 19295
rect 3985 19261 4019 19295
rect 4537 19261 4571 19295
rect 5549 19261 5583 19295
rect 6837 19261 6871 19295
rect 7849 19261 7883 19295
rect 8033 19261 8067 19295
rect 10333 19261 10367 19295
rect 11161 19261 11195 19295
rect 12541 19261 12575 19295
rect 13645 19261 13679 19295
rect 13912 19261 13946 19295
rect 15577 19261 15611 19295
rect 16773 19261 16807 19295
rect 17233 19261 17267 19295
rect 17877 19261 17911 19295
rect 18245 19261 18279 19295
rect 20996 19261 21030 19295
rect 25053 19261 25087 19295
rect 25237 19261 25271 19295
rect 25789 19261 25823 19295
rect 1961 19193 1995 19227
rect 2605 19193 2639 19227
rect 2697 19193 2731 19227
rect 4721 19193 4755 19227
rect 6653 19193 6687 19227
rect 8300 19193 8334 19227
rect 10885 19193 10919 19227
rect 18512 19193 18546 19227
rect 22753 19193 22787 19227
rect 24041 19193 24075 19227
rect 24225 19193 24259 19227
rect 24317 19193 24351 19227
rect 24685 19193 24719 19227
rect 2135 19125 2169 19159
rect 3065 19125 3099 19159
rect 4169 19125 4203 19159
rect 4537 19125 4571 19159
rect 4997 19125 5031 19159
rect 5733 19125 5767 19159
rect 7481 19125 7515 19159
rect 9413 19125 9447 19159
rect 10057 19125 10091 19159
rect 11069 19125 11103 19159
rect 11529 19125 11563 19159
rect 11897 19125 11931 19159
rect 12725 19125 12759 19159
rect 13185 19125 13219 19159
rect 15025 19125 15059 19159
rect 16037 19125 16071 19159
rect 16681 19125 16715 19159
rect 20177 19125 20211 19159
rect 23489 19125 23523 19159
rect 25421 19125 25455 19159
rect 26249 19125 26283 19159
rect 2495 18921 2529 18955
rect 2973 18921 3007 18955
rect 4721 18921 4755 18955
rect 6009 18921 6043 18955
rect 6101 18921 6135 18955
rect 9137 18921 9171 18955
rect 11805 18921 11839 18955
rect 13921 18921 13955 18955
rect 16405 18921 16439 18955
rect 18153 18921 18187 18955
rect 19901 18921 19935 18955
rect 20729 18921 20763 18955
rect 22017 18921 22051 18955
rect 25421 18921 25455 18955
rect 1961 18853 1995 18887
rect 3709 18853 3743 18887
rect 5273 18853 5307 18887
rect 5457 18853 5491 18887
rect 1409 18717 1443 18751
rect 2881 18717 2915 18751
rect 3065 18717 3099 18751
rect 5549 18717 5583 18751
rect 2329 18649 2363 18683
rect 4997 18649 5031 18683
rect 7021 18853 7055 18887
rect 8585 18853 8619 18887
rect 9505 18853 9539 18887
rect 13461 18853 13495 18887
rect 15853 18853 15887 18887
rect 17417 18853 17451 18887
rect 18981 18853 19015 18887
rect 19073 18853 19107 18887
rect 20177 18853 20211 18887
rect 21465 18853 21499 18887
rect 23029 18853 23063 18887
rect 24593 18853 24627 18887
rect 25053 18853 25087 18887
rect 10692 18785 10726 18819
rect 13553 18785 13587 18819
rect 15117 18785 15151 18819
rect 15669 18785 15703 18819
rect 15945 18785 15979 18819
rect 16681 18785 16715 18819
rect 17509 18785 17543 18819
rect 18797 18785 18831 18819
rect 21557 18785 21591 18819
rect 23121 18785 23155 18819
rect 7021 18717 7055 18751
rect 7113 18717 7147 18751
rect 8493 18717 8527 18751
rect 8677 18717 8711 18751
rect 10425 18717 10459 18751
rect 13369 18717 13403 18751
rect 14657 18717 14691 18751
rect 17325 18717 17359 18751
rect 21465 18717 21499 18751
rect 22937 18717 22971 18751
rect 24593 18717 24627 18751
rect 24685 18717 24719 18751
rect 6377 18649 6411 18683
rect 8125 18649 8159 18683
rect 15393 18649 15427 18683
rect 16957 18649 16991 18683
rect 18521 18649 18555 18683
rect 21005 18649 21039 18683
rect 22569 18649 22603 18683
rect 4353 18581 4387 18615
rect 6101 18581 6135 18615
rect 6561 18581 6595 18615
rect 7481 18581 7515 18615
rect 7849 18581 7883 18615
rect 9965 18581 9999 18615
rect 10241 18581 10275 18615
rect 12449 18581 12483 18615
rect 12725 18581 12759 18615
rect 13001 18581 13035 18615
rect 14289 18581 14323 18615
rect 19533 18581 19567 18615
rect 22385 18581 22419 18615
rect 23673 18581 23707 18615
rect 24133 18581 24167 18615
rect 2237 18377 2271 18411
rect 3801 18377 3835 18411
rect 4169 18377 4203 18411
rect 6285 18377 6319 18411
rect 8125 18377 8159 18411
rect 8585 18377 8619 18411
rect 9781 18377 9815 18411
rect 12541 18377 12575 18411
rect 13461 18377 13495 18411
rect 14197 18377 14231 18411
rect 15669 18377 15703 18411
rect 17049 18377 17083 18411
rect 19073 18377 19107 18411
rect 19441 18377 19475 18411
rect 21373 18377 21407 18411
rect 21925 18377 21959 18411
rect 22201 18377 22235 18411
rect 22661 18377 22695 18411
rect 23489 18377 23523 18411
rect 25053 18377 25087 18411
rect 25421 18377 25455 18411
rect 25789 18377 25823 18411
rect 2789 18309 2823 18343
rect 6929 18309 6963 18343
rect 18153 18309 18187 18343
rect 2605 18241 2639 18275
rect 3249 18241 3283 18275
rect 4261 18241 4295 18275
rect 7481 18241 7515 18275
rect 9873 18241 9907 18275
rect 11989 18241 12023 18275
rect 13001 18241 13035 18275
rect 14289 18241 14323 18275
rect 17785 18241 17819 18275
rect 18613 18241 18647 18275
rect 1409 18173 1443 18207
rect 6653 18173 6687 18207
rect 8401 18173 8435 18207
rect 1685 18105 1719 18139
rect 3341 18105 3375 18139
rect 4528 18105 4562 18139
rect 7205 18105 7239 18139
rect 7389 18105 7423 18139
rect 10140 18105 10174 18139
rect 13093 18173 13127 18207
rect 16865 18173 16899 18207
rect 18705 18173 18739 18207
rect 19993 18173 20027 18207
rect 20249 18173 20283 18207
rect 14556 18105 14590 18139
rect 23765 18309 23799 18343
rect 26249 18309 26283 18343
rect 24317 18241 24351 18275
rect 22477 18173 22511 18207
rect 24041 18173 24075 18207
rect 25237 18173 25271 18207
rect 23029 18105 23063 18139
rect 24225 18105 24259 18139
rect 3249 18037 3283 18071
rect 5641 18037 5675 18071
rect 9045 18037 9079 18071
rect 9413 18037 9447 18071
rect 11253 18037 11287 18071
rect 11805 18037 11839 18071
rect 11989 18037 12023 18071
rect 12265 18037 12299 18071
rect 13001 18037 13035 18071
rect 16221 18037 16255 18071
rect 16773 18037 16807 18071
rect 17417 18037 17451 18071
rect 18613 18037 18647 18071
rect 19901 18037 19935 18071
rect 22201 18037 22235 18071
rect 22293 18037 22327 18071
rect 24685 18037 24719 18071
rect 1961 17833 1995 17867
rect 3525 17833 3559 17867
rect 3801 17833 3835 17867
rect 6929 17833 6963 17867
rect 7297 17833 7331 17867
rect 8493 17833 8527 17867
rect 12541 17833 12575 17867
rect 13461 17833 13495 17867
rect 15117 17833 15151 17867
rect 15761 17833 15795 17867
rect 18061 17833 18095 17867
rect 18613 17833 18647 17867
rect 20729 17833 20763 17867
rect 21925 17833 21959 17867
rect 22293 17833 22327 17867
rect 23673 17833 23707 17867
rect 24593 17833 24627 17867
rect 25053 17833 25087 17867
rect 2329 17765 2363 17799
rect 2973 17765 3007 17799
rect 8033 17765 8067 17799
rect 8309 17765 8343 17799
rect 9505 17765 9539 17799
rect 10333 17765 10367 17799
rect 11897 17765 11931 17799
rect 13277 17765 13311 17799
rect 16948 17765 16982 17799
rect 19809 17765 19843 17799
rect 21281 17765 21315 17799
rect 21465 17765 21499 17799
rect 22845 17765 22879 17799
rect 23029 17765 23063 17799
rect 25421 17765 25455 17799
rect 4905 17697 4939 17731
rect 5264 17697 5298 17731
rect 1409 17629 1443 17663
rect 2973 17629 3007 17663
rect 3065 17629 3099 17663
rect 4997 17629 5031 17663
rect 7941 17629 7975 17663
rect 8125 17629 8159 17663
rect 10149 17697 10183 17731
rect 11989 17697 12023 17731
rect 15577 17697 15611 17731
rect 16681 17697 16715 17731
rect 19901 17697 19935 17731
rect 24409 17697 24443 17731
rect 25789 17697 25823 17731
rect 10425 17629 10459 17663
rect 11897 17629 11931 17663
rect 13553 17629 13587 17663
rect 19717 17629 19751 17663
rect 21557 17629 21591 17663
rect 23121 17629 23155 17663
rect 24685 17629 24719 17663
rect 8309 17561 8343 17595
rect 9873 17561 9907 17595
rect 11437 17561 11471 17595
rect 14381 17561 14415 17595
rect 16221 17561 16255 17595
rect 19073 17561 19107 17595
rect 20361 17561 20395 17595
rect 24133 17561 24167 17595
rect 2513 17493 2547 17527
rect 4353 17493 4387 17527
rect 6377 17493 6411 17527
rect 7573 17493 7607 17527
rect 8953 17493 8987 17527
rect 10793 17493 10827 17527
rect 11161 17493 11195 17527
rect 13001 17493 13035 17527
rect 13921 17493 13955 17527
rect 14657 17493 14691 17527
rect 16589 17493 16623 17527
rect 19349 17493 19383 17527
rect 21005 17493 21039 17527
rect 22569 17493 22603 17527
rect 4353 17289 4387 17323
rect 5273 17289 5307 17323
rect 6929 17289 6963 17323
rect 12541 17289 12575 17323
rect 13553 17289 13587 17323
rect 14105 17289 14139 17323
rect 16221 17289 16255 17323
rect 17049 17289 17083 17323
rect 19993 17289 20027 17323
rect 23029 17289 23063 17323
rect 23765 17289 23799 17323
rect 25421 17289 25455 17323
rect 2789 17221 2823 17255
rect 4169 17221 4203 17255
rect 8585 17221 8619 17255
rect 10149 17221 10183 17255
rect 12173 17221 12207 17255
rect 15577 17221 15611 17255
rect 16773 17221 16807 17255
rect 17509 17221 17543 17255
rect 19073 17221 19107 17255
rect 20637 17221 20671 17255
rect 24685 17221 24719 17255
rect 4813 17153 4847 17187
rect 6285 17153 6319 17187
rect 7481 17153 7515 17187
rect 8769 17153 8803 17187
rect 11345 17153 11379 17187
rect 12081 17153 12115 17187
rect 13001 17153 13035 17187
rect 14197 17153 14231 17187
rect 18797 17153 18831 17187
rect 19533 17153 19567 17187
rect 19625 17153 19659 17187
rect 21097 17153 21131 17187
rect 22477 17153 22511 17187
rect 24133 17153 24167 17187
rect 1409 17085 1443 17119
rect 1685 17085 1719 17119
rect 2513 17085 2547 17119
rect 4905 17085 4939 17119
rect 3065 17017 3099 17051
rect 3249 17017 3283 17051
rect 3341 17017 3375 17051
rect 4813 17017 4847 17051
rect 7205 17017 7239 17051
rect 7389 17017 7423 17051
rect 7941 17017 7975 17051
rect 8309 17017 8343 17051
rect 9036 17017 9070 17051
rect 16865 17085 16899 17119
rect 21189 17085 21223 17119
rect 22293 17085 22327 17119
rect 25237 17085 25271 17119
rect 25789 17085 25823 17119
rect 13001 17017 13035 17051
rect 13093 17017 13127 17051
rect 14442 17017 14476 17051
rect 24317 17017 24351 17051
rect 25053 17017 25087 17051
rect 3709 16949 3743 16983
rect 5641 16949 5675 16983
rect 6653 16949 6687 16983
rect 10885 16949 10919 16983
rect 11161 16949 11195 16983
rect 11805 16949 11839 16983
rect 12081 16949 12115 16983
rect 17877 16949 17911 16983
rect 18521 16949 18555 16983
rect 19533 16949 19567 16983
rect 20361 16949 20395 16983
rect 21097 16949 21131 16983
rect 21557 16949 21591 16983
rect 22109 16949 22143 16983
rect 23489 16949 23523 16983
rect 24225 16949 24259 16983
rect 2329 16745 2363 16779
rect 3433 16745 3467 16779
rect 3893 16745 3927 16779
rect 5457 16745 5491 16779
rect 6929 16745 6963 16779
rect 8493 16745 8527 16779
rect 9873 16745 9907 16779
rect 10701 16745 10735 16779
rect 12449 16745 12483 16779
rect 13635 16745 13669 16779
rect 15025 16745 15059 16779
rect 15853 16745 15887 16779
rect 18889 16745 18923 16779
rect 19441 16745 19475 16779
rect 20545 16745 20579 16779
rect 22845 16745 22879 16779
rect 23949 16745 23983 16779
rect 24869 16745 24903 16779
rect 25145 16745 25179 16779
rect 2973 16677 3007 16711
rect 7358 16677 7392 16711
rect 11314 16677 11348 16711
rect 13461 16677 13495 16711
rect 14105 16677 14139 16711
rect 15669 16677 15703 16711
rect 17776 16677 17810 16711
rect 20269 16677 20303 16711
rect 1409 16609 1443 16643
rect 2789 16609 2823 16643
rect 3065 16609 3099 16643
rect 4344 16609 4378 16643
rect 6561 16609 6595 16643
rect 7113 16609 7147 16643
rect 9045 16609 9079 16643
rect 9505 16609 9539 16643
rect 9689 16609 9723 16643
rect 13001 16609 13035 16643
rect 14197 16609 14231 16643
rect 16313 16609 16347 16643
rect 16681 16609 16715 16643
rect 17509 16609 17543 16643
rect 21180 16609 21214 16643
rect 23765 16609 23799 16643
rect 24961 16609 24995 16643
rect 4077 16541 4111 16575
rect 11069 16541 11103 16575
rect 14013 16541 14047 16575
rect 15945 16541 15979 16575
rect 20913 16541 20947 16575
rect 24041 16541 24075 16575
rect 15393 16473 15427 16507
rect 17049 16473 17083 16507
rect 19901 16473 19935 16507
rect 24409 16473 24443 16507
rect 1961 16405 1995 16439
rect 2513 16405 2547 16439
rect 6009 16405 6043 16439
rect 10333 16405 10367 16439
rect 14657 16405 14691 16439
rect 22293 16405 22327 16439
rect 23213 16405 23247 16439
rect 23489 16405 23523 16439
rect 1593 16201 1627 16235
rect 2513 16201 2547 16235
rect 4537 16201 4571 16235
rect 5181 16201 5215 16235
rect 6561 16201 6595 16235
rect 9137 16201 9171 16235
rect 12173 16201 12207 16235
rect 13553 16201 13587 16235
rect 13921 16201 13955 16235
rect 16037 16201 16071 16235
rect 17233 16201 17267 16235
rect 17509 16201 17543 16235
rect 22293 16201 22327 16235
rect 23029 16201 23063 16235
rect 23489 16201 23523 16235
rect 24961 16201 24995 16235
rect 25421 16201 25455 16235
rect 2145 16133 2179 16167
rect 10333 16133 10367 16167
rect 12541 16133 12575 16167
rect 23765 16133 23799 16167
rect 5733 16065 5767 16099
rect 6101 16065 6135 16099
rect 10885 16065 10919 16099
rect 13093 16065 13127 16099
rect 24133 16065 24167 16099
rect 24317 16065 24351 16099
rect 1409 15997 1443 16031
rect 2605 15997 2639 16031
rect 5457 15997 5491 16031
rect 7757 15997 7791 16031
rect 10149 15997 10183 16031
rect 10609 15997 10643 16031
rect 14565 15997 14599 16031
rect 14657 15997 14691 16031
rect 18337 15997 18371 16031
rect 18429 15997 18463 16031
rect 20913 15997 20947 16031
rect 21180 15997 21214 16031
rect 25237 15997 25271 16031
rect 25789 15997 25823 16031
rect 2850 15929 2884 15963
rect 5641 15929 5675 15963
rect 8002 15929 8036 15963
rect 12817 15929 12851 15963
rect 14924 15929 14958 15963
rect 18674 15929 18708 15963
rect 20453 15929 20487 15963
rect 20821 15929 20855 15963
rect 3985 15861 4019 15895
rect 4997 15861 5031 15895
rect 7205 15861 7239 15895
rect 7573 15861 7607 15895
rect 9689 15861 9723 15895
rect 10793 15861 10827 15895
rect 11345 15861 11379 15895
rect 11805 15861 11839 15895
rect 13001 15861 13035 15895
rect 16589 15861 16623 15895
rect 19809 15861 19843 15895
rect 24225 15861 24259 15895
rect 1961 15657 1995 15691
rect 3893 15657 3927 15691
rect 4261 15657 4295 15691
rect 5181 15657 5215 15691
rect 5641 15657 5675 15691
rect 6745 15657 6779 15691
rect 7297 15657 7331 15691
rect 8309 15657 8343 15691
rect 9873 15657 9907 15691
rect 10333 15657 10367 15691
rect 10977 15657 11011 15691
rect 13093 15657 13127 15691
rect 13461 15657 13495 15691
rect 14105 15657 14139 15691
rect 15025 15657 15059 15691
rect 17141 15657 17175 15691
rect 17877 15657 17911 15691
rect 18429 15657 18463 15691
rect 21465 15657 21499 15691
rect 23029 15657 23063 15691
rect 23673 15657 23707 15691
rect 24041 15657 24075 15691
rect 2973 15589 3007 15623
rect 3525 15589 3559 15623
rect 5273 15589 5307 15623
rect 6561 15589 6595 15623
rect 14197 15589 14231 15623
rect 15669 15589 15703 15623
rect 15853 15589 15887 15623
rect 16773 15589 16807 15623
rect 17693 15589 17727 15623
rect 19441 15589 19475 15623
rect 24685 15589 24719 15623
rect 25145 15589 25179 15623
rect 1409 15521 1443 15555
rect 3065 15521 3099 15555
rect 8125 15521 8159 15555
rect 9137 15521 9171 15555
rect 9689 15521 9723 15555
rect 11325 15521 11359 15555
rect 14749 15521 14783 15555
rect 15945 15521 15979 15555
rect 21905 15521 21939 15555
rect 24777 15521 24811 15555
rect 2881 15453 2915 15487
rect 5181 15453 5215 15487
rect 6837 15453 6871 15487
rect 8401 15453 8435 15487
rect 8769 15453 8803 15487
rect 11069 15453 11103 15487
rect 14105 15453 14139 15487
rect 17969 15453 18003 15487
rect 19349 15453 19383 15487
rect 19533 15453 19567 15487
rect 19901 15453 19935 15487
rect 21649 15453 21683 15487
rect 24685 15453 24719 15487
rect 2513 15385 2547 15419
rect 4721 15385 4755 15419
rect 6285 15385 6319 15419
rect 13645 15385 13679 15419
rect 15393 15385 15427 15419
rect 20269 15385 20303 15419
rect 20729 15385 20763 15419
rect 24225 15385 24259 15419
rect 6101 15317 6135 15351
rect 7665 15317 7699 15351
rect 7849 15317 7883 15351
rect 12449 15317 12483 15351
rect 16405 15317 16439 15351
rect 17417 15317 17451 15351
rect 18981 15317 19015 15351
rect 21189 15317 21223 15351
rect 1777 15113 1811 15147
rect 3341 15113 3375 15147
rect 4353 15113 4387 15147
rect 4905 15113 4939 15147
rect 6285 15113 6319 15147
rect 6561 15113 6595 15147
rect 7021 15113 7055 15147
rect 7481 15113 7515 15147
rect 10517 15113 10551 15147
rect 13645 15113 13679 15147
rect 14105 15113 14139 15147
rect 15209 15113 15243 15147
rect 17509 15113 17543 15147
rect 17785 15113 17819 15147
rect 18981 15113 19015 15147
rect 21005 15113 21039 15147
rect 21649 15113 21683 15147
rect 23029 15113 23063 15147
rect 23397 15113 23431 15147
rect 23765 15113 23799 15147
rect 24777 15113 24811 15147
rect 2053 15045 2087 15079
rect 4721 15045 4755 15079
rect 12541 15045 12575 15079
rect 2605 14977 2639 15011
rect 5457 14977 5491 15011
rect 9965 14977 9999 15011
rect 11069 14977 11103 15011
rect 11897 14977 11931 15011
rect 12909 14977 12943 15011
rect 2329 14909 2363 14943
rect 3525 14909 3559 14943
rect 5181 14909 5215 14943
rect 6837 14909 6871 14943
rect 7941 14909 7975 14943
rect 13093 14909 13127 14943
rect 2513 14841 2547 14875
rect 3801 14841 3835 14875
rect 5917 14841 5951 14875
rect 8208 14841 8242 14875
rect 10333 14841 10367 14875
rect 10793 14841 10827 14875
rect 10977 14841 11011 14875
rect 12265 14841 12299 14875
rect 13001 14841 13035 14875
rect 14381 14841 14415 14875
rect 14657 14841 14691 14875
rect 15025 14841 15059 14875
rect 18521 15045 18555 15079
rect 16957 14977 16991 15011
rect 18061 14977 18095 15011
rect 22109 14977 22143 15011
rect 24317 14977 24351 15011
rect 15945 14909 15979 14943
rect 19073 14909 19107 14943
rect 22201 14909 22235 14943
rect 22569 14909 22603 14943
rect 25053 14909 25087 14943
rect 25237 14909 25271 14943
rect 25973 14909 26007 14943
rect 16479 14841 16513 14875
rect 16957 14841 16991 14875
rect 17049 14841 17083 14875
rect 19340 14841 19374 14875
rect 22109 14841 22143 14875
rect 24041 14841 24075 14875
rect 25513 14841 25547 14875
rect 3065 14773 3099 14807
rect 5365 14773 5399 14807
rect 7849 14773 7883 14807
rect 9321 14773 9355 14807
rect 11529 14773 11563 14807
rect 14565 14773 14599 14807
rect 15209 14773 15243 14807
rect 15393 14773 15427 14807
rect 16313 14773 16347 14807
rect 20453 14773 20487 14807
rect 21465 14773 21499 14807
rect 24225 14773 24259 14807
rect 2881 14569 2915 14603
rect 6653 14569 6687 14603
rect 6929 14569 6963 14603
rect 8861 14569 8895 14603
rect 10241 14569 10275 14603
rect 11161 14569 11195 14603
rect 11805 14569 11839 14603
rect 16681 14569 16715 14603
rect 18337 14569 18371 14603
rect 19441 14569 19475 14603
rect 19901 14569 19935 14603
rect 20269 14569 20303 14603
rect 20729 14569 20763 14603
rect 22753 14569 22787 14603
rect 24685 14569 24719 14603
rect 5733 14501 5767 14535
rect 8401 14501 8435 14535
rect 9229 14501 9263 14535
rect 15546 14501 15580 14535
rect 21465 14501 21499 14535
rect 21557 14501 21591 14535
rect 21925 14501 21959 14535
rect 1501 14433 1535 14467
rect 1768 14433 1802 14467
rect 4077 14433 4111 14467
rect 5549 14433 5583 14467
rect 6745 14433 6779 14467
rect 7389 14433 7423 14467
rect 12153 14433 12187 14467
rect 15301 14433 15335 14467
rect 19717 14433 19751 14467
rect 23561 14433 23595 14467
rect 5089 14365 5123 14399
rect 5825 14365 5859 14399
rect 8401 14365 8435 14399
rect 8493 14365 8527 14399
rect 10149 14365 10183 14399
rect 10333 14365 10367 14399
rect 11897 14365 11931 14399
rect 18245 14365 18279 14399
rect 18429 14365 18463 14399
rect 21465 14365 21499 14399
rect 23305 14365 23339 14399
rect 3893 14297 3927 14331
rect 5273 14297 5307 14331
rect 6285 14297 6319 14331
rect 7941 14297 7975 14331
rect 14473 14297 14507 14331
rect 17417 14297 17451 14331
rect 21005 14297 21039 14331
rect 3433 14229 3467 14263
rect 4261 14229 4295 14263
rect 4721 14229 4755 14263
rect 7757 14229 7791 14263
rect 9781 14229 9815 14263
rect 10793 14229 10827 14263
rect 13277 14229 13311 14263
rect 14013 14229 14047 14263
rect 14749 14229 14783 14263
rect 17877 14229 17911 14263
rect 19073 14229 19107 14263
rect 22293 14229 22327 14263
rect 23029 14229 23063 14263
rect 25237 14229 25271 14263
rect 3065 14025 3099 14059
rect 3709 14025 3743 14059
rect 6653 14025 6687 14059
rect 7113 14025 7147 14059
rect 9965 14025 9999 14059
rect 10517 14025 10551 14059
rect 14473 14025 14507 14059
rect 16497 14025 16531 14059
rect 18521 14025 18555 14059
rect 20637 14025 20671 14059
rect 21189 14025 21223 14059
rect 23029 14025 23063 14059
rect 23765 14025 23799 14059
rect 25421 14025 25455 14059
rect 8125 13957 8159 13991
rect 17417 13957 17451 13991
rect 22109 13957 22143 13991
rect 1685 13889 1719 13923
rect 4077 13889 4111 13923
rect 4169 13889 4203 13923
rect 7665 13889 7699 13923
rect 16313 13889 16347 13923
rect 16957 13889 16991 13923
rect 17049 13889 17083 13923
rect 17877 13889 17911 13923
rect 21005 13889 21039 13923
rect 21557 13889 21591 13923
rect 21741 13889 21775 13923
rect 24133 13889 24167 13923
rect 8401 13821 8435 13855
rect 8585 13821 8619 13855
rect 8852 13821 8886 13855
rect 13093 13821 13127 13855
rect 15945 13821 15979 13855
rect 18613 13821 18647 13855
rect 22661 13821 22695 13855
rect 24317 13821 24351 13855
rect 25053 13821 25087 13855
rect 25237 13821 25271 13855
rect 25789 13821 25823 13855
rect 1952 13753 1986 13787
rect 4414 13753 4448 13787
rect 7389 13753 7423 13787
rect 7573 13753 7607 13787
rect 11345 13753 11379 13787
rect 13338 13753 13372 13787
rect 16957 13753 16991 13787
rect 18880 13753 18914 13787
rect 5549 13685 5583 13719
rect 6101 13685 6135 13719
rect 11161 13685 11195 13719
rect 11989 13685 12023 13719
rect 13001 13685 13035 13719
rect 15393 13685 15427 13719
rect 19993 13685 20027 13719
rect 21649 13685 21683 13719
rect 23489 13685 23523 13719
rect 24225 13685 24259 13719
rect 24685 13685 24719 13719
rect 1869 13481 1903 13515
rect 2237 13481 2271 13515
rect 2973 13481 3007 13515
rect 5273 13481 5307 13515
rect 8585 13481 8619 13515
rect 9873 13481 9907 13515
rect 13185 13481 13219 13515
rect 14197 13481 14231 13515
rect 16497 13481 16531 13515
rect 16773 13481 16807 13515
rect 19441 13481 19475 13515
rect 21465 13481 21499 13515
rect 22293 13481 22327 13515
rect 24041 13481 24075 13515
rect 25329 13481 25363 13515
rect 3065 13413 3099 13447
rect 5917 13413 5951 13447
rect 8677 13413 8711 13447
rect 11713 13413 11747 13447
rect 15945 13413 15979 13447
rect 17224 13413 17258 13447
rect 18981 13413 19015 13447
rect 21281 13413 21315 13447
rect 22928 13413 22962 13447
rect 4077 13345 4111 13379
rect 5733 13345 5767 13379
rect 6929 13345 6963 13379
rect 9689 13345 9723 13379
rect 11529 13345 11563 13379
rect 14657 13345 14691 13379
rect 15117 13345 15151 13379
rect 15761 13345 15795 13379
rect 16957 13345 16991 13379
rect 22017 13345 22051 13379
rect 22668 13345 22702 13379
rect 25145 13345 25179 13379
rect 1409 13277 1443 13311
rect 2973 13277 3007 13311
rect 3525 13277 3559 13311
rect 4353 13277 4387 13311
rect 6009 13277 6043 13311
rect 8585 13277 8619 13311
rect 11805 13277 11839 13311
rect 12541 13277 12575 13311
rect 14197 13277 14231 13311
rect 14289 13277 14323 13311
rect 16037 13277 16071 13311
rect 21557 13277 21591 13311
rect 24961 13277 24995 13311
rect 2513 13209 2547 13243
rect 4905 13209 4939 13243
rect 5457 13209 5491 13243
rect 6745 13209 6779 13243
rect 7113 13209 7147 13243
rect 8125 13209 8159 13243
rect 9505 13209 9539 13243
rect 11253 13209 11287 13243
rect 13737 13209 13771 13243
rect 15485 13209 15519 13243
rect 21005 13209 21039 13243
rect 3893 13141 3927 13175
rect 6377 13141 6411 13175
rect 7573 13141 7607 13175
rect 7849 13141 7883 13175
rect 9045 13141 9079 13175
rect 10517 13141 10551 13175
rect 10885 13141 10919 13175
rect 13553 13141 13587 13175
rect 18337 13141 18371 13175
rect 19349 13141 19383 13175
rect 20085 13141 20119 13175
rect 20729 13141 20763 13175
rect 24593 13141 24627 13175
rect 1777 12937 1811 12971
rect 5273 12937 5307 12971
rect 6009 12937 6043 12971
rect 6285 12937 6319 12971
rect 7205 12937 7239 12971
rect 8125 12937 8159 12971
rect 8585 12937 8619 12971
rect 9689 12937 9723 12971
rect 10333 12937 10367 12971
rect 12173 12937 12207 12971
rect 13461 12937 13495 12971
rect 14105 12937 14139 12971
rect 15485 12937 15519 12971
rect 16497 12937 16531 12971
rect 17509 12937 17543 12971
rect 19441 12937 19475 12971
rect 19717 12937 19751 12971
rect 19809 12937 19843 12971
rect 21649 12937 21683 12971
rect 23765 12937 23799 12971
rect 24685 12937 24719 12971
rect 25421 12937 25455 12971
rect 3341 12869 3375 12903
rect 5089 12869 5123 12903
rect 3893 12801 3927 12835
rect 4353 12801 4387 12835
rect 5825 12801 5859 12835
rect 2053 12733 2087 12767
rect 4721 12733 4755 12767
rect 8769 12869 8803 12903
rect 10885 12869 10919 12903
rect 13921 12869 13955 12903
rect 16313 12869 16347 12903
rect 18521 12869 18555 12903
rect 7757 12801 7791 12835
rect 11253 12801 11287 12835
rect 11805 12801 11839 12835
rect 12909 12801 12943 12835
rect 14473 12801 14507 12835
rect 15117 12801 15151 12835
rect 15945 12801 15979 12835
rect 17049 12801 17083 12835
rect 19073 12801 19107 12835
rect 20085 12869 20119 12903
rect 21097 12869 21131 12903
rect 25789 12869 25823 12903
rect 20637 12801 20671 12835
rect 22201 12801 22235 12835
rect 24317 12801 24351 12835
rect 7481 12733 7515 12767
rect 9045 12733 9079 12767
rect 9321 12733 9355 12767
rect 10609 12733 10643 12767
rect 11437 12733 11471 12767
rect 14657 12733 14691 12767
rect 16773 12733 16807 12767
rect 17877 12733 17911 12767
rect 19717 12733 19751 12767
rect 20361 12733 20395 12767
rect 25237 12733 25271 12767
rect 26157 12733 26191 12767
rect 2329 12665 2363 12699
rect 3157 12665 3191 12699
rect 3617 12665 3651 12699
rect 5549 12665 5583 12699
rect 5733 12665 5767 12699
rect 6009 12665 6043 12699
rect 6653 12665 6687 12699
rect 7665 12665 7699 12699
rect 11345 12665 11379 12699
rect 12523 12665 12557 12699
rect 13001 12665 13035 12699
rect 13093 12665 13127 12699
rect 14565 12665 14599 12699
rect 18337 12665 18371 12699
rect 18797 12665 18831 12699
rect 21925 12665 21959 12699
rect 24041 12665 24075 12699
rect 2237 12597 2271 12631
rect 2789 12597 2823 12631
rect 3801 12597 3835 12631
rect 9229 12597 9263 12631
rect 16957 12597 16991 12631
rect 18981 12597 19015 12631
rect 20545 12597 20579 12631
rect 21373 12597 21407 12631
rect 22109 12597 22143 12631
rect 22661 12597 22695 12631
rect 23121 12597 23155 12631
rect 23489 12597 23523 12631
rect 24225 12597 24259 12631
rect 25053 12597 25087 12631
rect 1409 12393 1443 12427
rect 1961 12393 1995 12427
rect 2329 12393 2363 12427
rect 3525 12393 3559 12427
rect 5273 12393 5307 12427
rect 5733 12393 5767 12427
rect 7205 12393 7239 12427
rect 8677 12393 8711 12427
rect 9045 12393 9079 12427
rect 9321 12393 9355 12427
rect 15669 12393 15703 12427
rect 17233 12393 17267 12427
rect 18521 12393 18555 12427
rect 21005 12393 21039 12427
rect 23397 12393 23431 12427
rect 23949 12393 23983 12427
rect 2789 12325 2823 12359
rect 2973 12325 3007 12359
rect 4629 12325 4663 12359
rect 4813 12325 4847 12359
rect 4905 12325 4939 12359
rect 6377 12325 6411 12359
rect 8217 12325 8251 12359
rect 6193 12257 6227 12291
rect 8033 12257 8067 12291
rect 3065 12189 3099 12223
rect 5549 12189 5583 12223
rect 6469 12189 6503 12223
rect 8309 12189 8343 12223
rect 2513 12121 2547 12155
rect 4353 12121 4387 12155
rect 9689 12325 9723 12359
rect 12725 12325 12759 12359
rect 13737 12325 13771 12359
rect 16098 12325 16132 12359
rect 19165 12325 19199 12359
rect 20269 12325 20303 12359
rect 20729 12325 20763 12359
rect 25053 12325 25087 12359
rect 10609 12257 10643 12291
rect 10968 12257 11002 12291
rect 13093 12257 13127 12291
rect 19257 12257 19291 12291
rect 22017 12257 22051 12291
rect 22284 12257 22318 12291
rect 10701 12189 10735 12223
rect 13737 12189 13771 12223
rect 13829 12189 13863 12223
rect 14933 12189 14967 12223
rect 15853 12189 15887 12223
rect 19165 12189 19199 12223
rect 24317 12189 24351 12223
rect 24961 12189 24995 12223
rect 25145 12189 25179 12223
rect 9413 12121 9447 12155
rect 14565 12121 14599 12155
rect 25513 12121 25547 12155
rect 3801 12053 3835 12087
rect 5549 12053 5583 12087
rect 5917 12053 5951 12087
rect 7573 12053 7607 12087
rect 7757 12053 7791 12087
rect 9321 12053 9355 12087
rect 10241 12053 10275 12087
rect 12081 12053 12115 12087
rect 13277 12053 13311 12087
rect 14289 12053 14323 12087
rect 17785 12053 17819 12087
rect 18705 12053 18739 12087
rect 19993 12053 20027 12087
rect 21557 12053 21591 12087
rect 24593 12053 24627 12087
rect 2789 11849 2823 11883
rect 5641 11849 5675 11883
rect 6377 11849 6411 11883
rect 8493 11849 8527 11883
rect 10517 11849 10551 11883
rect 15209 11849 15243 11883
rect 19441 11849 19475 11883
rect 21557 11849 21591 11883
rect 22569 11849 22603 11883
rect 25053 11849 25087 11883
rect 4169 11781 4203 11815
rect 6193 11781 6227 11815
rect 3249 11713 3283 11747
rect 4261 11713 4295 11747
rect 1409 11645 1443 11679
rect 2513 11645 2547 11679
rect 3341 11645 3375 11679
rect 1685 11577 1719 11611
rect 3249 11577 3283 11611
rect 3801 11577 3835 11611
rect 4506 11577 4540 11611
rect 6929 11781 6963 11815
rect 10333 11781 10367 11815
rect 10701 11781 10735 11815
rect 16405 11781 16439 11815
rect 18429 11781 18463 11815
rect 19993 11781 20027 11815
rect 8953 11713 8987 11747
rect 10149 11713 10183 11747
rect 7481 11645 7515 11679
rect 7849 11645 7883 11679
rect 8217 11645 8251 11679
rect 9045 11645 9079 11679
rect 9413 11645 9447 11679
rect 7205 11577 7239 11611
rect 8953 11577 8987 11611
rect 11253 11713 11287 11747
rect 15853 11713 15887 11747
rect 16773 11713 16807 11747
rect 18889 11713 18923 11747
rect 22109 11713 22143 11747
rect 23489 11713 23523 11747
rect 23673 11713 23707 11747
rect 10977 11645 11011 11679
rect 12725 11645 12759 11679
rect 13737 11645 13771 11679
rect 13829 11645 13863 11679
rect 17877 11645 17911 11679
rect 18981 11645 19015 11679
rect 20545 11645 20579 11679
rect 21005 11645 21039 11679
rect 25605 11645 25639 11679
rect 11161 11577 11195 11611
rect 11713 11577 11747 11611
rect 13369 11577 13403 11611
rect 14096 11577 14130 11611
rect 16957 11577 16991 11611
rect 17325 11577 17359 11611
rect 18889 11577 18923 11611
rect 20269 11577 20303 11611
rect 20453 11577 20487 11611
rect 21833 11577 21867 11611
rect 22017 11577 22051 11611
rect 23121 11577 23155 11611
rect 23940 11577 23974 11611
rect 6377 11509 6411 11543
rect 6653 11509 6687 11543
rect 7389 11509 7423 11543
rect 10333 11509 10367 11543
rect 12173 11509 12207 11543
rect 12909 11509 12943 11543
rect 16221 11509 16255 11543
rect 16865 11509 16899 11543
rect 19717 11509 19751 11543
rect 21281 11509 21315 11543
rect 25973 11509 26007 11543
rect 1409 11305 1443 11339
rect 1961 11305 1995 11339
rect 2329 11305 2363 11339
rect 3433 11305 3467 11339
rect 3801 11305 3835 11339
rect 6009 11305 6043 11339
rect 7757 11305 7791 11339
rect 15853 11305 15887 11339
rect 18429 11305 18463 11339
rect 20177 11305 20211 11339
rect 20729 11305 20763 11339
rect 21465 11305 21499 11339
rect 22293 11305 22327 11339
rect 24593 11305 24627 11339
rect 2973 11237 3007 11271
rect 3065 11237 3099 11271
rect 7113 11237 7147 11271
rect 10302 11237 10336 11271
rect 12808 11237 12842 11271
rect 16488 11237 16522 11271
rect 18705 11237 18739 11271
rect 19717 11237 19751 11271
rect 21925 11237 21959 11271
rect 22845 11237 22879 11271
rect 23029 11237 23063 11271
rect 24685 11237 24719 11271
rect 4077 11169 4111 11203
rect 4344 11169 4378 11203
rect 6929 11169 6963 11203
rect 8125 11169 8159 11203
rect 10057 11169 10091 11203
rect 12541 11169 12575 11203
rect 15025 11169 15059 11203
rect 16221 11169 16255 11203
rect 19809 11169 19843 11203
rect 21557 11169 21591 11203
rect 24409 11169 24443 11203
rect 25789 11169 25823 11203
rect 2973 11101 3007 11135
rect 7205 11101 7239 11135
rect 8309 11101 8343 11135
rect 9229 11101 9263 11135
rect 12449 11101 12483 11135
rect 15485 11101 15519 11135
rect 19717 11101 19751 11135
rect 21465 11101 21499 11135
rect 23121 11101 23155 11135
rect 25053 11101 25087 11135
rect 2513 11033 2547 11067
rect 5457 11033 5491 11067
rect 6653 11033 6687 11067
rect 8861 11033 8895 11067
rect 11437 11033 11471 11067
rect 17601 11033 17635 11067
rect 19257 11033 19291 11067
rect 21005 11033 21039 11067
rect 22569 11033 22603 11067
rect 24133 11033 24167 11067
rect 6469 10965 6503 10999
rect 9873 10965 9907 10999
rect 12081 10965 12115 10999
rect 13921 10965 13955 10999
rect 14657 10965 14691 10999
rect 23673 10965 23707 10999
rect 25421 10965 25455 10999
rect 1869 10761 1903 10795
rect 3249 10761 3283 10795
rect 5641 10761 5675 10795
rect 9137 10761 9171 10795
rect 10057 10761 10091 10795
rect 11621 10761 11655 10795
rect 12265 10761 12299 10795
rect 14565 10761 14599 10795
rect 15853 10761 15887 10795
rect 16497 10761 16531 10795
rect 17417 10761 17451 10795
rect 18429 10761 18463 10795
rect 18613 10761 18647 10795
rect 21465 10761 21499 10795
rect 21741 10761 21775 10795
rect 22753 10761 22787 10795
rect 23489 10761 23523 10795
rect 24685 10761 24719 10795
rect 10333 10693 10367 10727
rect 11345 10693 11379 10727
rect 12725 10693 12759 10727
rect 14749 10693 14783 10727
rect 19533 10693 19567 10727
rect 20177 10693 20211 10727
rect 21189 10693 21223 10727
rect 23765 10693 23799 10727
rect 2421 10625 2455 10659
rect 3341 10625 3375 10659
rect 10701 10625 10735 10659
rect 13737 10625 13771 10659
rect 14197 10625 14231 10659
rect 17049 10625 17083 10659
rect 19073 10625 19107 10659
rect 22201 10625 22235 10659
rect 23029 10625 23063 10659
rect 25053 10625 25087 10659
rect 25513 10625 25547 10659
rect 1685 10557 1719 10591
rect 7757 10557 7791 10591
rect 8013 10557 8047 10591
rect 13461 10557 13495 10591
rect 15301 10557 15335 10591
rect 24317 10557 24351 10591
rect 25237 10557 25271 10591
rect 25973 10557 26007 10591
rect 2145 10489 2179 10523
rect 2329 10489 2363 10523
rect 2881 10489 2915 10523
rect 3586 10489 3620 10523
rect 6561 10489 6595 10523
rect 10885 10489 10919 10523
rect 13167 10489 13201 10523
rect 13645 10489 13679 10523
rect 15025 10489 15059 10523
rect 16221 10489 16255 10523
rect 16773 10489 16807 10523
rect 17877 10489 17911 10523
rect 19165 10489 19199 10523
rect 20453 10489 20487 10523
rect 20729 10489 20763 10523
rect 22293 10489 22327 10523
rect 24041 10489 24075 10523
rect 4721 10421 4755 10455
rect 5273 10421 5307 10455
rect 6009 10421 6043 10455
rect 7021 10421 7055 10455
rect 7573 10421 7607 10455
rect 9781 10421 9815 10455
rect 10793 10421 10827 10455
rect 15209 10421 15243 10455
rect 16957 10421 16991 10455
rect 19073 10421 19107 10455
rect 19993 10421 20027 10455
rect 20637 10421 20671 10455
rect 22201 10421 22235 10455
rect 24225 10421 24259 10455
rect 1961 10217 1995 10251
rect 2329 10217 2363 10251
rect 3617 10217 3651 10251
rect 4353 10217 4387 10251
rect 5273 10217 5307 10251
rect 7665 10217 7699 10251
rect 8861 10217 8895 10251
rect 12633 10217 12667 10251
rect 16405 10217 16439 10251
rect 16865 10217 16899 10251
rect 18337 10217 18371 10251
rect 19533 10217 19567 10251
rect 20637 10217 20671 10251
rect 22293 10217 22327 10251
rect 22661 10217 22695 10251
rect 22937 10217 22971 10251
rect 25329 10217 25363 10251
rect 25697 10217 25731 10251
rect 2973 10149 3007 10183
rect 3065 10149 3099 10183
rect 5089 10149 5123 10183
rect 6193 10149 6227 10183
rect 6530 10149 6564 10183
rect 10241 10149 10275 10183
rect 10333 10149 10367 10183
rect 12725 10149 12759 10183
rect 14197 10149 14231 10183
rect 15945 10149 15979 10183
rect 17509 10149 17543 10183
rect 17969 10149 18003 10183
rect 19073 10149 19107 10183
rect 20085 10149 20119 10183
rect 21158 10149 21192 10183
rect 5365 10081 5399 10115
rect 6285 10081 6319 10115
rect 9137 10081 9171 10115
rect 13185 10081 13219 10115
rect 13553 10081 13587 10115
rect 16037 10081 16071 10115
rect 1409 10013 1443 10047
rect 2973 10013 3007 10047
rect 5733 10013 5767 10047
rect 10241 10013 10275 10047
rect 11529 10013 11563 10047
rect 12633 10013 12667 10047
rect 14197 10013 14231 10047
rect 14289 10013 14323 10047
rect 15945 10013 15979 10047
rect 17417 10013 17451 10047
rect 17601 10013 17635 10047
rect 19073 10013 19107 10047
rect 19165 10013 19199 10047
rect 20913 10013 20947 10047
rect 2513 9945 2547 9979
rect 4813 9945 4847 9979
rect 9781 9945 9815 9979
rect 12173 9945 12207 9979
rect 13737 9945 13771 9979
rect 15025 9945 15059 9979
rect 15485 9945 15519 9979
rect 18613 9945 18647 9979
rect 23664 10081 23698 10115
rect 23397 10013 23431 10047
rect 24777 9945 24811 9979
rect 8493 9877 8527 9911
rect 10793 9877 10827 9911
rect 11253 9877 11287 9911
rect 11897 9877 11931 9911
rect 14657 9877 14691 9911
rect 17049 9877 17083 9911
rect 22661 9877 22695 9911
rect 23213 9877 23247 9911
rect 26065 9877 26099 9911
rect 4629 9673 4663 9707
rect 6929 9673 6963 9707
rect 7849 9673 7883 9707
rect 16865 9673 16899 9707
rect 17509 9673 17543 9707
rect 18337 9673 18371 9707
rect 20913 9673 20947 9707
rect 24501 9673 24535 9707
rect 2145 9605 2179 9639
rect 3709 9605 3743 9639
rect 5273 9605 5307 9639
rect 8493 9605 8527 9639
rect 10885 9605 10919 9639
rect 12081 9605 12115 9639
rect 13829 9605 13863 9639
rect 14749 9605 14783 9639
rect 17785 9605 17819 9639
rect 22661 9605 22695 9639
rect 1961 9537 1995 9571
rect 2605 9537 2639 9571
rect 4261 9537 4295 9571
rect 5733 9537 5767 9571
rect 8309 9537 8343 9571
rect 9045 9537 9079 9571
rect 11437 9537 11471 9571
rect 14289 9537 14323 9571
rect 21925 9537 21959 9571
rect 23121 9537 23155 9571
rect 2697 9469 2731 9503
rect 3985 9469 4019 9503
rect 6377 9469 6411 9503
rect 10149 9469 10183 9503
rect 11161 9469 11195 9503
rect 12633 9469 12667 9503
rect 13645 9469 13679 9503
rect 15393 9469 15427 9503
rect 15485 9469 15519 9503
rect 15741 9469 15775 9503
rect 18797 9469 18831 9503
rect 19064 9469 19098 9503
rect 21649 9469 21683 9503
rect 22109 9469 22143 9503
rect 22385 9469 22419 9503
rect 23489 9469 23523 9503
rect 24041 9469 24075 9503
rect 5733 9401 5767 9435
rect 5825 9401 5859 9435
rect 7205 9401 7239 9435
rect 7389 9401 7423 9435
rect 7481 9401 7515 9435
rect 8769 9401 8803 9435
rect 8953 9401 8987 9435
rect 9781 9401 9815 9435
rect 14289 9401 14323 9435
rect 14381 9401 14415 9435
rect 21833 9401 21867 9435
rect 23747 9401 23781 9435
rect 24225 9401 24259 9435
rect 24317 9401 24351 9435
rect 2605 9333 2639 9367
rect 3065 9333 3099 9367
rect 3525 9333 3559 9367
rect 4169 9333 4203 9367
rect 5089 9333 5123 9367
rect 6285 9333 6319 9367
rect 6377 9333 6411 9367
rect 6561 9333 6595 9367
rect 10609 9333 10643 9367
rect 11345 9333 11379 9367
rect 12817 9333 12851 9367
rect 13277 9333 13311 9367
rect 18613 9333 18647 9367
rect 20177 9333 20211 9367
rect 21355 9333 21389 9367
rect 22109 9333 22143 9367
rect 25053 9605 25087 9639
rect 25973 9537 26007 9571
rect 25237 9469 25271 9503
rect 25513 9401 25547 9435
rect 24501 9333 24535 9367
rect 24685 9333 24719 9367
rect 26341 9333 26375 9367
rect 2145 9129 2179 9163
rect 3709 9129 3743 9163
rect 4629 9129 4663 9163
rect 9873 9129 9907 9163
rect 10333 9129 10367 9163
rect 13369 9129 13403 9163
rect 16957 9129 16991 9163
rect 17509 9129 17543 9163
rect 18429 9129 18463 9163
rect 19533 9129 19567 9163
rect 20361 9129 20395 9163
rect 21833 9129 21867 9163
rect 24593 9129 24627 9163
rect 25329 9129 25363 9163
rect 2973 9061 3007 9095
rect 4445 9061 4479 9095
rect 10977 9061 11011 9095
rect 11069 9061 11103 9095
rect 15844 9061 15878 9095
rect 19073 9061 19107 9095
rect 19165 9061 19199 9095
rect 20729 9061 20763 9095
rect 21465 9061 21499 9095
rect 21557 9061 21591 9095
rect 3065 8993 3099 9027
rect 5089 8993 5123 9027
rect 5908 8993 5942 9027
rect 7573 8993 7607 9027
rect 8493 8993 8527 9027
rect 11989 8993 12023 9027
rect 12245 8993 12279 9027
rect 15025 8993 15059 9027
rect 15577 8993 15611 9027
rect 18889 8993 18923 9027
rect 21281 8993 21315 9027
rect 1409 8925 1443 8959
rect 2881 8925 2915 8959
rect 4721 8925 4755 8959
rect 5641 8925 5675 8959
rect 9413 8925 9447 8959
rect 10977 8925 11011 8959
rect 4169 8857 4203 8891
rect 8677 8857 8711 8891
rect 10517 8857 10551 8891
rect 14381 8857 14415 8891
rect 21005 8857 21039 8891
rect 22569 9061 22603 9095
rect 25697 9061 25731 9095
rect 22661 8993 22695 9027
rect 22928 8993 22962 9027
rect 25145 8993 25179 9027
rect 26065 8925 26099 8959
rect 24961 8857 24995 8891
rect 2513 8789 2547 8823
rect 5549 8789 5583 8823
rect 7021 8789 7055 8823
rect 7941 8789 7975 8823
rect 8309 8789 8343 8823
rect 9045 8789 9079 8823
rect 11437 8789 11471 8823
rect 11805 8789 11839 8823
rect 14013 8789 14047 8823
rect 14657 8789 14691 8823
rect 17969 8789 18003 8823
rect 18613 8789 18647 8823
rect 19993 8789 20027 8823
rect 21833 8789 21867 8823
rect 22017 8789 22051 8823
rect 24041 8789 24075 8823
rect 2421 8585 2455 8619
rect 3801 8585 3835 8619
rect 5273 8585 5307 8619
rect 5641 8585 5675 8619
rect 6929 8585 6963 8619
rect 11345 8585 11379 8619
rect 14381 8585 14415 8619
rect 15577 8585 15611 8619
rect 15761 8585 15795 8619
rect 17049 8585 17083 8619
rect 17877 8585 17911 8619
rect 20085 8585 20119 8619
rect 21281 8585 21315 8619
rect 23765 8585 23799 8619
rect 24685 8585 24719 8619
rect 25881 8585 25915 8619
rect 26157 8585 26191 8619
rect 2237 8517 2271 8551
rect 3985 8517 4019 8551
rect 4997 8517 5031 8551
rect 6101 8517 6135 8551
rect 8861 8517 8895 8551
rect 13829 8517 13863 8551
rect 16681 8517 16715 8551
rect 17417 8517 17451 8551
rect 20821 8517 20855 8551
rect 21005 8517 21039 8551
rect 23489 8517 23523 8551
rect 25053 8517 25087 8551
rect 25421 8517 25455 8551
rect 1869 8449 1903 8483
rect 2881 8449 2915 8483
rect 3433 8449 3467 8483
rect 7297 8449 7331 8483
rect 9045 8449 9079 8483
rect 11161 8449 11195 8483
rect 12449 8449 12483 8483
rect 15209 8449 15243 8483
rect 16313 8449 16347 8483
rect 4261 8381 4295 8415
rect 5457 8381 5491 8415
rect 6653 8381 6687 8415
rect 7481 8381 7515 8415
rect 11069 8381 11103 8415
rect 2881 8313 2915 8347
rect 2973 8313 3007 8347
rect 4537 8313 4571 8347
rect 7941 8313 7975 8347
rect 8493 8313 8527 8347
rect 9290 8313 9324 8347
rect 18705 8381 18739 8415
rect 18972 8381 19006 8415
rect 21557 8381 21591 8415
rect 22201 8381 22235 8415
rect 25237 8381 25271 8415
rect 11805 8313 11839 8347
rect 12173 8313 12207 8347
rect 12694 8313 12728 8347
rect 14749 8313 14783 8347
rect 16037 8313 16071 8347
rect 16221 8313 16255 8347
rect 20821 8313 20855 8347
rect 21833 8313 21867 8347
rect 23121 8313 23155 8347
rect 24041 8313 24075 8347
rect 24225 8313 24259 8347
rect 24317 8313 24351 8347
rect 4445 8245 4479 8279
rect 7389 8245 7423 8279
rect 10425 8245 10459 8279
rect 11161 8245 11195 8279
rect 18521 8245 18555 8279
rect 21741 8245 21775 8279
rect 22753 8245 22787 8279
rect 1961 8041 1995 8075
rect 5089 8041 5123 8075
rect 9137 8041 9171 8075
rect 12081 8041 12115 8075
rect 12541 8041 12575 8075
rect 15025 8041 15059 8075
rect 15761 8041 15795 8075
rect 18981 8041 19015 8075
rect 19349 8041 19383 8075
rect 19993 8041 20027 8075
rect 20913 8041 20947 8075
rect 21741 8041 21775 8075
rect 24225 8041 24259 8075
rect 24961 8041 24995 8075
rect 25789 8041 25823 8075
rect 26249 8041 26283 8075
rect 2973 7973 3007 8007
rect 4629 7973 4663 8007
rect 7380 7973 7414 8007
rect 10140 7973 10174 8007
rect 16589 7973 16623 8007
rect 18429 7973 18463 8007
rect 22192 7973 22226 8007
rect 25421 7973 25455 8007
rect 2789 7905 2823 7939
rect 5825 7905 5859 7939
rect 12633 7905 12667 7939
rect 12900 7905 12934 7939
rect 18521 7905 18555 7939
rect 19441 7905 19475 7939
rect 20729 7905 20763 7939
rect 23857 7905 23891 7939
rect 1409 7837 1443 7871
rect 3065 7837 3099 7871
rect 4629 7837 4663 7871
rect 4721 7837 4755 7871
rect 6101 7837 6135 7871
rect 7113 7837 7147 7871
rect 9873 7837 9907 7871
rect 16589 7837 16623 7871
rect 16681 7837 16715 7871
rect 18429 7837 18463 7871
rect 21925 7837 21959 7871
rect 24869 7837 24903 7871
rect 25053 7837 25087 7871
rect 2513 7769 2547 7803
rect 4169 7769 4203 7803
rect 11253 7769 11287 7803
rect 14013 7769 14047 7803
rect 19625 7769 19659 7803
rect 24501 7769 24535 7803
rect 2329 7701 2363 7735
rect 3525 7701 3559 7735
rect 3893 7701 3927 7735
rect 5641 7701 5675 7735
rect 6929 7701 6963 7735
rect 8493 7701 8527 7735
rect 9413 7701 9447 7735
rect 14657 7701 14691 7735
rect 16129 7701 16163 7735
rect 17049 7701 17083 7735
rect 17417 7701 17451 7735
rect 17969 7701 18003 7735
rect 21465 7701 21499 7735
rect 23305 7701 23339 7735
rect 2237 7497 2271 7531
rect 4905 7497 4939 7531
rect 6285 7497 6319 7531
rect 6561 7497 6595 7531
rect 9413 7497 9447 7531
rect 10701 7497 10735 7531
rect 11069 7497 11103 7531
rect 12265 7497 12299 7531
rect 16405 7497 16439 7531
rect 16957 7497 16991 7531
rect 18245 7497 18279 7531
rect 18705 7497 18739 7531
rect 21097 7497 21131 7531
rect 21741 7497 21775 7531
rect 22753 7497 22787 7531
rect 23489 7497 23523 7531
rect 24685 7497 24719 7531
rect 25053 7497 25087 7531
rect 25421 7497 25455 7531
rect 10333 7429 10367 7463
rect 13001 7429 13035 7463
rect 13553 7429 13587 7463
rect 18981 7429 19015 7463
rect 23765 7429 23799 7463
rect 5457 7361 5491 7395
rect 5825 7361 5859 7395
rect 6837 7361 6871 7395
rect 9229 7361 9263 7395
rect 9965 7361 9999 7395
rect 12449 7361 12483 7395
rect 14841 7361 14875 7395
rect 15025 7361 15059 7395
rect 19165 7361 19199 7395
rect 21465 7361 21499 7395
rect 22109 7361 22143 7395
rect 22293 7361 22327 7395
rect 24225 7361 24259 7395
rect 24317 7361 24351 7395
rect 26249 7361 26283 7395
rect 1869 7293 1903 7327
rect 2329 7293 2363 7327
rect 4629 7293 4663 7327
rect 5181 7293 5215 7327
rect 7104 7293 7138 7327
rect 9689 7293 9723 7327
rect 11241 7293 11275 7327
rect 14105 7293 14139 7327
rect 18061 7293 18095 7327
rect 23121 7293 23155 7327
rect 25237 7293 25271 7327
rect 2574 7225 2608 7259
rect 5365 7225 5399 7259
rect 9873 7225 9907 7259
rect 11897 7225 11931 7259
rect 13829 7225 13863 7259
rect 15270 7225 15304 7259
rect 19410 7225 19444 7259
rect 22201 7225 22235 7259
rect 24225 7225 24259 7259
rect 3709 7157 3743 7191
rect 4353 7157 4387 7191
rect 8217 7157 8251 7191
rect 8861 7157 8895 7191
rect 11437 7157 11471 7191
rect 13369 7157 13403 7191
rect 14013 7157 14047 7191
rect 14565 7157 14599 7191
rect 17417 7157 17451 7191
rect 17877 7157 17911 7191
rect 20545 7157 20579 7191
rect 25789 7157 25823 7191
rect 7665 6953 7699 6987
rect 8401 6953 8435 6987
rect 14473 6953 14507 6987
rect 15117 6953 15151 6987
rect 22385 6953 22419 6987
rect 2973 6885 3007 6919
rect 5273 6885 5307 6919
rect 6837 6885 6871 6919
rect 10241 6885 10275 6919
rect 15945 6885 15979 6919
rect 16405 6885 16439 6919
rect 21465 6885 21499 6919
rect 23029 6885 23063 6919
rect 23121 6885 23155 6919
rect 24593 6885 24627 6919
rect 1409 6817 1443 6851
rect 2329 6817 2363 6851
rect 7389 6817 7423 6851
rect 11069 6817 11103 6851
rect 11437 6817 11471 6851
rect 12541 6817 12575 6851
rect 12808 6817 12842 6851
rect 15761 6817 15795 6851
rect 16957 6817 16991 6851
rect 17224 6817 17258 6851
rect 19257 6817 19291 6851
rect 19717 6817 19751 6851
rect 21925 6817 21959 6851
rect 23489 6817 23523 6851
rect 23857 6817 23891 6851
rect 24685 6817 24719 6851
rect 25421 6817 25455 6851
rect 26249 6817 26283 6851
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 5273 6749 5307 6783
rect 5365 6749 5399 6783
rect 5825 6749 5859 6783
rect 6745 6749 6779 6783
rect 6929 6749 6963 6783
rect 8309 6749 8343 6783
rect 8493 6749 8527 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 16037 6749 16071 6783
rect 19625 6749 19659 6783
rect 21465 6749 21499 6783
rect 21557 6749 21591 6783
rect 23029 6749 23063 6783
rect 24593 6749 24627 6783
rect 25789 6749 25823 6783
rect 2513 6681 2547 6715
rect 6193 6681 6227 6715
rect 7941 6681 7975 6715
rect 19901 6681 19935 6715
rect 21005 6681 21039 6715
rect 22569 6681 22603 6715
rect 24133 6681 24167 6715
rect 1869 6613 1903 6647
rect 3433 6613 3467 6647
rect 3893 6613 3927 6647
rect 4353 6613 4387 6647
rect 4813 6613 4847 6647
rect 6377 6613 6411 6647
rect 8953 6613 8987 6647
rect 9505 6613 9539 6647
rect 9781 6613 9815 6647
rect 10701 6613 10735 6647
rect 11621 6613 11655 6647
rect 12081 6613 12115 6647
rect 12449 6613 12483 6647
rect 13921 6613 13955 6647
rect 15485 6613 15519 6647
rect 16865 6613 16899 6647
rect 18337 6613 18371 6647
rect 20269 6613 20303 6647
rect 20637 6613 20671 6647
rect 25053 6613 25087 6647
rect 4445 6409 4479 6443
rect 6929 6409 6963 6443
rect 7941 6409 7975 6443
rect 8585 6409 8619 6443
rect 10149 6409 10183 6443
rect 10793 6409 10827 6443
rect 11805 6409 11839 6443
rect 12265 6409 12299 6443
rect 13001 6409 13035 6443
rect 14841 6409 14875 6443
rect 15853 6409 15887 6443
rect 19533 6409 19567 6443
rect 20913 6409 20947 6443
rect 25421 6409 25455 6443
rect 6009 6341 6043 6375
rect 16221 6341 16255 6375
rect 16497 6341 16531 6375
rect 18153 6341 18187 6375
rect 19717 6341 19751 6375
rect 21281 6341 21315 6375
rect 23857 6341 23891 6375
rect 1777 6273 1811 6307
rect 1869 6273 1903 6307
rect 4905 6273 4939 6307
rect 7389 6273 7423 6307
rect 8769 6273 8803 6307
rect 11161 6273 11195 6307
rect 16865 6273 16899 6307
rect 18613 6273 18647 6307
rect 19165 6273 19199 6307
rect 20269 6273 20303 6307
rect 21833 6273 21867 6307
rect 24041 6273 24075 6307
rect 25973 6273 26007 6307
rect 2136 6205 2170 6239
rect 4261 6205 4295 6239
rect 4997 6205 5031 6239
rect 11253 6205 11287 6239
rect 13461 6205 13495 6239
rect 17049 6205 17083 6239
rect 17785 6205 17819 6239
rect 19993 6205 20027 6239
rect 21557 6205 21591 6239
rect 4905 6137 4939 6171
rect 7481 6137 7515 6171
rect 9014 6137 9048 6171
rect 13277 6137 13311 6171
rect 13728 6137 13762 6171
rect 16957 6137 16991 6171
rect 18705 6137 18739 6171
rect 20177 6137 20211 6171
rect 21741 6137 21775 6171
rect 22569 6137 22603 6171
rect 24286 6137 24320 6171
rect 3249 6069 3283 6103
rect 3893 6069 3927 6103
rect 5457 6069 5491 6103
rect 6285 6069 6319 6103
rect 7389 6069 7423 6103
rect 8309 6069 8343 6103
rect 11437 6069 11471 6103
rect 12449 6069 12483 6103
rect 15393 6069 15427 6103
rect 17509 6069 17543 6103
rect 18613 6069 18647 6103
rect 22937 6069 22971 6103
rect 23489 6069 23523 6103
rect 26341 6069 26375 6103
rect 1961 5865 1995 5899
rect 2513 5865 2547 5899
rect 2789 5865 2823 5899
rect 8861 5865 8895 5899
rect 10241 5865 10275 5899
rect 11327 5865 11361 5899
rect 12541 5865 12575 5899
rect 13553 5865 13587 5899
rect 14749 5865 14783 5899
rect 15117 5865 15151 5899
rect 16313 5865 16347 5899
rect 17601 5865 17635 5899
rect 17969 5865 18003 5899
rect 19073 5865 19107 5899
rect 19901 5865 19935 5899
rect 20729 5865 20763 5899
rect 21189 5865 21223 5899
rect 22661 5865 22695 5899
rect 23213 5865 23247 5899
rect 23581 5865 23615 5899
rect 24317 5865 24351 5899
rect 25881 5865 25915 5899
rect 1777 5797 1811 5831
rect 2053 5797 2087 5831
rect 4690 5797 4724 5831
rect 10057 5797 10091 5831
rect 10793 5797 10827 5831
rect 11621 5797 11655 5831
rect 11805 5797 11839 5831
rect 14197 5797 14231 5831
rect 14289 5797 14323 5831
rect 17049 5797 17083 5831
rect 17141 5797 17175 5831
rect 18613 5797 18647 5831
rect 7196 5729 7230 5763
rect 10333 5729 10367 5763
rect 15393 5729 15427 5763
rect 15945 5729 15979 5763
rect 16865 5729 16899 5763
rect 19717 5729 19751 5763
rect 21537 5729 21571 5763
rect 24133 5729 24167 5763
rect 25329 5729 25363 5763
rect 2973 5661 3007 5695
rect 4445 5661 4479 5695
rect 6929 5661 6963 5695
rect 11897 5661 11931 5695
rect 14197 5661 14231 5695
rect 18613 5661 18647 5695
rect 18705 5661 18739 5695
rect 21281 5661 21315 5695
rect 24409 5661 24443 5695
rect 25145 5661 25179 5695
rect 1501 5593 1535 5627
rect 9781 5593 9815 5627
rect 13737 5593 13771 5627
rect 15577 5593 15611 5627
rect 18153 5593 18187 5627
rect 19625 5593 19659 5627
rect 24869 5593 24903 5627
rect 3525 5525 3559 5559
rect 3893 5525 3927 5559
rect 4261 5525 4295 5559
rect 5825 5525 5859 5559
rect 6377 5525 6411 5559
rect 6745 5525 6779 5559
rect 8309 5525 8343 5559
rect 9321 5525 9355 5559
rect 11069 5525 11103 5559
rect 12909 5525 12943 5559
rect 16589 5525 16623 5559
rect 20269 5525 20303 5559
rect 23857 5525 23891 5559
rect 25513 5525 25547 5559
rect 26249 5525 26283 5559
rect 1501 5321 1535 5355
rect 2513 5321 2547 5355
rect 4353 5321 4387 5355
rect 5273 5321 5307 5355
rect 6929 5321 6963 5355
rect 10057 5321 10091 5355
rect 11345 5321 11379 5355
rect 11621 5321 11655 5355
rect 13737 5321 13771 5355
rect 14105 5321 14139 5355
rect 17509 5321 17543 5355
rect 17877 5321 17911 5355
rect 18153 5321 18187 5355
rect 19717 5321 19751 5355
rect 21373 5321 21407 5355
rect 22017 5321 22051 5355
rect 23121 5321 23155 5355
rect 23765 5321 23799 5355
rect 25973 5321 26007 5355
rect 8493 5253 8527 5287
rect 12541 5253 12575 5287
rect 19441 5253 19475 5287
rect 1961 5185 1995 5219
rect 2973 5185 3007 5219
rect 5733 5185 5767 5219
rect 7941 5185 7975 5219
rect 9045 5185 9079 5219
rect 10425 5185 10459 5219
rect 13001 5185 13035 5219
rect 14381 5185 14415 5219
rect 18521 5185 18555 5219
rect 18705 5185 18739 5219
rect 19993 5185 20027 5219
rect 24317 5185 24351 5219
rect 24777 5185 24811 5219
rect 25513 5185 25547 5219
rect 3240 5117 3274 5151
rect 5457 5117 5491 5151
rect 7481 5117 7515 5151
rect 9781 5117 9815 5151
rect 10609 5117 10643 5151
rect 12265 5117 12299 5151
rect 16865 5117 16899 5151
rect 20260 5117 20294 5151
rect 22477 5117 22511 5151
rect 25053 5117 25087 5151
rect 25237 5117 25271 5151
rect 2053 5049 2087 5083
rect 4997 5049 5031 5083
rect 7205 5049 7239 5083
rect 8309 5049 8343 5083
rect 8769 5049 8803 5083
rect 8953 5049 8987 5083
rect 13093 5049 13127 5083
rect 14648 5049 14682 5083
rect 16497 5049 16531 5083
rect 18613 5049 18647 5083
rect 22293 5049 22327 5083
rect 24041 5049 24075 5083
rect 1961 4981 1995 5015
rect 2881 4981 2915 5015
rect 6285 4981 6319 5015
rect 6561 4981 6595 5015
rect 7389 4981 7423 5015
rect 10517 4981 10551 5015
rect 13001 4981 13035 5015
rect 15761 4981 15795 5015
rect 17049 4981 17083 5015
rect 22661 4981 22695 5015
rect 23489 4981 23523 5015
rect 24225 4981 24259 5015
rect 26341 4981 26375 5015
rect 2145 4777 2179 4811
rect 5089 4777 5123 4811
rect 5733 4777 5767 4811
rect 6377 4777 6411 4811
rect 6929 4777 6963 4811
rect 8585 4777 8619 4811
rect 9137 4777 9171 4811
rect 9413 4777 9447 4811
rect 11253 4777 11287 4811
rect 11621 4777 11655 4811
rect 12633 4777 12667 4811
rect 14657 4777 14691 4811
rect 15853 4777 15887 4811
rect 16589 4777 16623 4811
rect 19717 4777 19751 4811
rect 22293 4777 22327 4811
rect 23857 4777 23891 4811
rect 24593 4777 24627 4811
rect 25789 4777 25823 4811
rect 26249 4777 26283 4811
rect 2789 4709 2823 4743
rect 2881 4709 2915 4743
rect 4629 4709 4663 4743
rect 7941 4709 7975 4743
rect 10057 4709 10091 4743
rect 10241 4709 10275 4743
rect 10333 4709 10367 4743
rect 10793 4709 10827 4743
rect 13553 4709 13587 4743
rect 14197 4709 14231 4743
rect 14289 4709 14323 4743
rect 15669 4709 15703 4743
rect 18604 4709 18638 4743
rect 21465 4709 21499 4743
rect 22845 4709 22879 4743
rect 23029 4709 23063 4743
rect 23121 4709 23155 4743
rect 6193 4641 6227 4675
rect 8401 4641 8435 4675
rect 8677 4641 8711 4675
rect 16957 4641 16991 4675
rect 18153 4641 18187 4675
rect 18337 4641 18371 4675
rect 24685 4641 24719 4675
rect 2789 4573 2823 4607
rect 4629 4573 4663 4607
rect 4721 4573 4755 4607
rect 6469 4573 6503 4607
rect 12633 4573 12667 4607
rect 12725 4573 12759 4607
rect 14197 4573 14231 4607
rect 15945 4573 15979 4607
rect 17141 4573 17175 4607
rect 21465 4573 21499 4607
rect 21557 4573 21591 4607
rect 21925 4573 21959 4607
rect 24593 4573 24627 4607
rect 2329 4505 2363 4539
rect 5917 4505 5951 4539
rect 8125 4505 8159 4539
rect 9781 4505 9815 4539
rect 12173 4505 12207 4539
rect 13737 4505 13771 4539
rect 15393 4505 15427 4539
rect 21005 4505 21039 4539
rect 24133 4505 24167 4539
rect 25053 4505 25087 4539
rect 1685 4437 1719 4471
rect 3433 4437 3467 4471
rect 3893 4437 3927 4471
rect 4169 4437 4203 4471
rect 7297 4437 7331 4471
rect 13185 4437 13219 4471
rect 15025 4437 15059 4471
rect 17785 4437 17819 4471
rect 20637 4437 20671 4471
rect 22569 4437 22603 4471
rect 25421 4437 25455 4471
rect 2145 4233 2179 4267
rect 3249 4233 3283 4267
rect 5457 4233 5491 4267
rect 6377 4233 6411 4267
rect 7113 4233 7147 4267
rect 8493 4233 8527 4267
rect 9045 4233 9079 4267
rect 12173 4233 12207 4267
rect 12725 4233 12759 4267
rect 13461 4233 13495 4267
rect 14381 4233 14415 4267
rect 14749 4233 14783 4267
rect 17417 4233 17451 4267
rect 21649 4233 21683 4267
rect 22017 4233 22051 4267
rect 22937 4233 22971 4267
rect 23765 4233 23799 4267
rect 3985 4165 4019 4199
rect 8769 4165 8803 4199
rect 10057 4165 10091 4199
rect 23213 4165 23247 4199
rect 2697 4097 2731 4131
rect 8033 4097 8067 4131
rect 9597 4097 9631 4131
rect 10977 4097 11011 4131
rect 11161 4097 11195 4131
rect 11805 4097 11839 4131
rect 13277 4097 13311 4131
rect 13829 4097 13863 4131
rect 14013 4097 14047 4131
rect 20269 4097 20303 4131
rect 20361 4097 20395 4131
rect 22293 4097 22327 4131
rect 25789 4097 25823 4131
rect 2421 4029 2455 4063
rect 4077 4029 4111 4063
rect 4333 4029 4367 4063
rect 6009 4029 6043 4063
rect 7665 4029 7699 4063
rect 9321 4029 9355 4063
rect 10591 4029 10625 4063
rect 14933 4029 14967 4063
rect 15189 4029 15223 4063
rect 16865 4029 16899 4063
rect 17877 4029 17911 4063
rect 18061 4029 18095 4063
rect 18317 4029 18351 4063
rect 2605 3961 2639 3995
rect 3617 3961 3651 3995
rect 7389 3961 7423 3995
rect 9505 3961 9539 3995
rect 13921 3961 13955 3995
rect 21189 4029 21223 4063
rect 22109 4029 22143 4063
rect 24041 4029 24075 4063
rect 25145 4029 25179 4063
rect 25237 4029 25271 4063
rect 20619 3961 20653 3995
rect 20913 3961 20947 3995
rect 24225 3961 24259 3995
rect 24317 3961 24351 3995
rect 1685 3893 1719 3927
rect 7573 3893 7607 3927
rect 10425 3893 10459 3927
rect 11069 3893 11103 3927
rect 16313 3893 16347 3927
rect 19441 3893 19475 3927
rect 19993 3893 20027 3927
rect 20269 3893 20303 3927
rect 21097 3893 21131 3927
rect 24685 3893 24719 3927
rect 25421 3893 25455 3927
rect 26249 3893 26283 3927
rect 5641 3689 5675 3723
rect 6285 3689 6319 3723
rect 10609 3689 10643 3723
rect 13461 3689 13495 3723
rect 14933 3689 14967 3723
rect 15853 3689 15887 3723
rect 17141 3689 17175 3723
rect 17509 3689 17543 3723
rect 18705 3689 18739 3723
rect 19809 3689 19843 3723
rect 20729 3689 20763 3723
rect 21925 3689 21959 3723
rect 22385 3689 22419 3723
rect 23029 3689 23063 3723
rect 23765 3689 23799 3723
rect 25421 3689 25455 3723
rect 26249 3689 26283 3723
rect 1685 3621 1719 3655
rect 2973 3621 3007 3655
rect 3249 3621 3283 3655
rect 3801 3621 3835 3655
rect 4528 3621 4562 3655
rect 14105 3621 14139 3655
rect 15669 3621 15703 3655
rect 15945 3621 15979 3655
rect 18061 3621 18095 3655
rect 18245 3621 18279 3655
rect 18337 3621 18371 3655
rect 21465 3621 21499 3655
rect 21557 3621 21591 3655
rect 24593 3621 24627 3655
rect 2789 3553 2823 3587
rect 4261 3553 4295 3587
rect 7021 3553 7055 3587
rect 7288 3553 7322 3587
rect 9781 3553 9815 3587
rect 10793 3553 10827 3587
rect 11325 3553 11359 3587
rect 14657 3553 14691 3587
rect 16865 3553 16899 3587
rect 19625 3553 19659 3587
rect 21281 3553 21315 3587
rect 23121 3553 23155 3587
rect 25789 3553 25823 3587
rect 3065 3485 3099 3519
rect 3249 3485 3283 3519
rect 10057 3485 10091 3519
rect 11069 3485 11103 3519
rect 13093 3485 13127 3519
rect 14105 3485 14139 3519
rect 14197 3485 14231 3519
rect 19901 3485 19935 3519
rect 20361 3485 20395 3519
rect 23029 3485 23063 3519
rect 24593 3485 24627 3519
rect 24685 3485 24719 3519
rect 25053 3485 25087 3519
rect 2513 3417 2547 3451
rect 10793 3417 10827 3451
rect 10885 3417 10919 3451
rect 13645 3417 13679 3451
rect 15393 3417 15427 3451
rect 17785 3417 17819 3451
rect 19349 3417 19383 3451
rect 21005 3417 21039 3451
rect 24133 3417 24167 3451
rect 2237 3349 2271 3383
rect 3525 3349 3559 3383
rect 6929 3349 6963 3383
rect 8401 3349 8435 3383
rect 9321 3349 9355 3383
rect 12449 3349 12483 3383
rect 16497 3349 16531 3383
rect 19073 3349 19107 3383
rect 22569 3349 22603 3383
rect 1501 3145 1535 3179
rect 2881 3145 2915 3179
rect 3801 3145 3835 3179
rect 4077 3145 4111 3179
rect 5641 3145 5675 3179
rect 6285 3145 6319 3179
rect 6929 3145 6963 3179
rect 7849 3145 7883 3179
rect 8401 3145 8435 3179
rect 8769 3145 8803 3179
rect 14381 3145 14415 3179
rect 14749 3145 14783 3179
rect 16865 3145 16899 3179
rect 17325 3145 17359 3179
rect 17693 3145 17727 3179
rect 18153 3145 18187 3179
rect 22569 3145 22603 3179
rect 23213 3145 23247 3179
rect 24685 3145 24719 3179
rect 26341 3145 26375 3179
rect 9045 3077 9079 3111
rect 16313 3077 16347 3111
rect 19717 3077 19751 3111
rect 21281 3077 21315 3111
rect 23765 3077 23799 3111
rect 1961 3009 1995 3043
rect 3249 3009 3283 3043
rect 4261 3009 4295 3043
rect 7481 3009 7515 3043
rect 9229 3009 9263 3043
rect 14933 3009 14967 3043
rect 18613 3009 18647 3043
rect 20177 3009 20211 3043
rect 21649 3009 21683 3043
rect 21833 3009 21867 3043
rect 24225 3009 24259 3043
rect 24317 3009 24351 3043
rect 25053 3009 25087 3043
rect 25421 3009 25455 3043
rect 2973 2941 3007 2975
rect 6653 2941 6687 2975
rect 9485 2941 9519 2975
rect 12081 2941 12115 2975
rect 12449 2941 12483 2975
rect 12716 2941 12750 2975
rect 20269 2941 20303 2975
rect 22845 2941 22879 2975
rect 25237 2941 25271 2975
rect 25973 2941 26007 2975
rect 2053 2873 2087 2907
rect 4506 2873 4540 2907
rect 7205 2873 7239 2907
rect 11897 2873 11931 2907
rect 15200 2873 15234 2907
rect 18613 2873 18647 2907
rect 18705 2873 18739 2907
rect 19165 2873 19199 2907
rect 19441 2873 19475 2907
rect 20177 2873 20211 2907
rect 20913 2873 20947 2907
rect 21741 2873 21775 2907
rect 24225 2873 24259 2907
rect 1961 2805 1995 2839
rect 2513 2805 2547 2839
rect 7389 2805 7423 2839
rect 10609 2805 10643 2839
rect 11161 2805 11195 2839
rect 12081 2805 12115 2839
rect 12173 2805 12207 2839
rect 13829 2805 13863 2839
rect 1961 2601 1995 2635
rect 2421 2601 2455 2635
rect 3801 2601 3835 2635
rect 5457 2601 5491 2635
rect 9597 2601 9631 2635
rect 11437 2601 11471 2635
rect 12449 2601 12483 2635
rect 16865 2601 16899 2635
rect 19809 2601 19843 2635
rect 22477 2601 22511 2635
rect 23765 2601 23799 2635
rect 25145 2601 25179 2635
rect 2053 2533 2087 2567
rect 4445 2533 4479 2567
rect 4629 2533 4663 2567
rect 4721 2533 4755 2567
rect 5089 2533 5123 2567
rect 6653 2533 6687 2567
rect 14381 2533 14415 2567
rect 14473 2533 14507 2567
rect 14841 2533 14875 2567
rect 18061 2533 18095 2567
rect 18705 2533 18739 2567
rect 18889 2533 18923 2567
rect 21741 2533 21775 2567
rect 24593 2533 24627 2567
rect 24685 2533 24719 2567
rect 1777 2465 1811 2499
rect 2881 2465 2915 2499
rect 3525 2465 3559 2499
rect 5733 2465 5767 2499
rect 7205 2465 7239 2499
rect 7472 2465 7506 2499
rect 10057 2465 10091 2499
rect 10324 2465 10358 2499
rect 11989 2465 12023 2499
rect 12725 2465 12759 2499
rect 15301 2465 15335 2499
rect 15752 2465 15786 2499
rect 19533 2465 19567 2499
rect 19993 2465 20027 2499
rect 21833 2465 21867 2499
rect 22753 2465 22787 2499
rect 23305 2465 23339 2499
rect 26065 2465 26099 2499
rect 2973 2397 3007 2431
rect 6285 2397 6319 2431
rect 9229 2397 9263 2431
rect 14289 2397 14323 2431
rect 15485 2397 15519 2431
rect 18981 2397 19015 2431
rect 20637 2397 20671 2431
rect 21741 2397 21775 2431
rect 24593 2397 24627 2431
rect 25421 2397 25455 2431
rect 25605 2397 25639 2431
rect 1501 2329 1535 2363
rect 4169 2329 4203 2363
rect 5917 2329 5951 2363
rect 21281 2329 21315 2363
rect 22937 2329 22971 2363
rect 24133 2329 24167 2363
rect 26433 2329 26467 2363
rect 8585 2261 8619 2295
rect 12909 2261 12943 2295
rect 13277 2261 13311 2295
rect 13645 2261 13679 2295
rect 13921 2261 13955 2295
rect 17693 2261 17727 2295
rect 18429 2261 18463 2295
rect 20177 2261 20211 2295
rect 20913 2261 20947 2295
<< metal1 >>
rect 10778 26800 10784 26852
rect 10836 26840 10842 26852
rect 17586 26840 17592 26852
rect 10836 26812 17592 26840
rect 10836 26800 10842 26812
rect 17586 26800 17592 26812
rect 17644 26800 17650 26852
rect 12437 26775 12495 26781
rect 12437 26741 12449 26775
rect 12483 26772 12495 26775
rect 25222 26772 25228 26784
rect 12483 26744 25228 26772
rect 12483 26741 12495 26744
rect 12437 26735 12495 26741
rect 25222 26732 25228 26744
rect 25280 26732 25286 26784
rect 7558 26664 7564 26716
rect 7616 26704 7622 26716
rect 9582 26704 9588 26716
rect 7616 26676 9588 26704
rect 7616 26664 7622 26676
rect 9582 26664 9588 26676
rect 9640 26664 9646 26716
rect 12069 26639 12127 26645
rect 12069 26605 12081 26639
rect 12115 26636 12127 26639
rect 12434 26636 12440 26648
rect 12115 26608 12440 26636
rect 12115 26605 12127 26608
rect 12069 26599 12127 26605
rect 12434 26596 12440 26608
rect 12492 26636 12498 26648
rect 19426 26636 19432 26648
rect 12492 26608 19432 26636
rect 12492 26596 12498 26608
rect 19426 26596 19432 26608
rect 19484 26596 19490 26648
rect 7558 26528 7564 26580
rect 7616 26568 7622 26580
rect 20806 26568 20812 26580
rect 7616 26540 20812 26568
rect 7616 26528 7622 26540
rect 20806 26528 20812 26540
rect 20864 26528 20870 26580
rect 11698 26460 11704 26512
rect 11756 26500 11762 26512
rect 24762 26500 24768 26512
rect 11756 26472 24768 26500
rect 11756 26460 11762 26472
rect 24762 26460 24768 26472
rect 24820 26460 24826 26512
rect 12161 26435 12219 26441
rect 12161 26401 12173 26435
rect 12207 26432 12219 26435
rect 13170 26432 13176 26444
rect 12207 26404 13176 26432
rect 12207 26401 12219 26404
rect 12161 26395 12219 26401
rect 13170 26392 13176 26404
rect 13228 26392 13234 26444
rect 11514 26324 11520 26376
rect 11572 26364 11578 26376
rect 12437 26367 12495 26373
rect 12437 26364 12449 26367
rect 11572 26336 12449 26364
rect 11572 26324 11578 26336
rect 12437 26333 12449 26336
rect 12483 26333 12495 26367
rect 12437 26327 12495 26333
rect 13354 26324 13360 26376
rect 13412 26364 13418 26376
rect 16022 26364 16028 26376
rect 13412 26336 16028 26364
rect 13412 26324 13418 26336
rect 16022 26324 16028 26336
rect 16080 26324 16086 26376
rect 4338 26256 4344 26308
rect 4396 26296 4402 26308
rect 20438 26296 20444 26308
rect 4396 26268 20444 26296
rect 4396 26256 4402 26268
rect 20438 26256 20444 26268
rect 20496 26256 20502 26308
rect 1302 26188 1308 26240
rect 1360 26228 1366 26240
rect 12437 26231 12495 26237
rect 12437 26228 12449 26231
rect 1360 26200 12449 26228
rect 1360 26188 1366 26200
rect 12437 26197 12449 26200
rect 12483 26197 12495 26231
rect 12437 26191 12495 26197
rect 14458 26188 14464 26240
rect 14516 26228 14522 26240
rect 19889 26231 19947 26237
rect 19889 26228 19901 26231
rect 14516 26200 19901 26228
rect 14516 26188 14522 26200
rect 19889 26197 19901 26200
rect 19935 26197 19947 26231
rect 19889 26191 19947 26197
rect 19981 26231 20039 26237
rect 19981 26197 19993 26231
rect 20027 26228 20039 26231
rect 25498 26228 25504 26240
rect 20027 26200 25504 26228
rect 20027 26197 20039 26200
rect 19981 26191 20039 26197
rect 25498 26188 25504 26200
rect 25556 26188 25562 26240
rect 4706 26120 4712 26172
rect 4764 26160 4770 26172
rect 9858 26160 9864 26172
rect 4764 26132 9864 26160
rect 4764 26120 4770 26132
rect 9858 26120 9864 26132
rect 9916 26120 9922 26172
rect 10042 26120 10048 26172
rect 10100 26160 10106 26172
rect 21542 26160 21548 26172
rect 10100 26132 21548 26160
rect 10100 26120 10106 26132
rect 21542 26120 21548 26132
rect 21600 26120 21606 26172
rect 7742 26052 7748 26104
rect 7800 26092 7806 26104
rect 17034 26092 17040 26104
rect 7800 26064 17040 26092
rect 7800 26052 7806 26064
rect 17034 26052 17040 26064
rect 17092 26052 17098 26104
rect 18874 26052 18880 26104
rect 18932 26092 18938 26104
rect 24302 26092 24308 26104
rect 18932 26064 24308 26092
rect 18932 26052 18938 26064
rect 24302 26052 24308 26064
rect 24360 26052 24366 26104
rect 3050 25984 3056 26036
rect 3108 26024 3114 26036
rect 7653 26027 7711 26033
rect 7653 26024 7665 26027
rect 3108 25996 7665 26024
rect 3108 25984 3114 25996
rect 7653 25993 7665 25996
rect 7699 25993 7711 26027
rect 7653 25987 7711 25993
rect 8754 25984 8760 26036
rect 8812 26024 8818 26036
rect 19794 26024 19800 26036
rect 8812 25996 19800 26024
rect 8812 25984 8818 25996
rect 19794 25984 19800 25996
rect 19852 25984 19858 26036
rect 19889 26027 19947 26033
rect 19889 25993 19901 26027
rect 19935 26024 19947 26027
rect 26050 26024 26056 26036
rect 19935 25996 26056 26024
rect 19935 25993 19947 25996
rect 19889 25987 19947 25993
rect 26050 25984 26056 25996
rect 26108 25984 26114 26036
rect 6914 25916 6920 25968
rect 6972 25956 6978 25968
rect 13906 25956 13912 25968
rect 6972 25928 13912 25956
rect 6972 25916 6978 25928
rect 13906 25916 13912 25928
rect 13964 25916 13970 25968
rect 15654 25916 15660 25968
rect 15712 25956 15718 25968
rect 17773 25959 17831 25965
rect 17773 25956 17785 25959
rect 15712 25928 17785 25956
rect 15712 25916 15718 25928
rect 17773 25925 17785 25928
rect 17819 25925 17831 25959
rect 17773 25919 17831 25925
rect 17862 25916 17868 25968
rect 17920 25956 17926 25968
rect 19981 25959 20039 25965
rect 19981 25956 19993 25959
rect 17920 25928 19993 25956
rect 17920 25916 17926 25928
rect 19981 25925 19993 25928
rect 20027 25925 20039 25959
rect 19981 25919 20039 25925
rect 1946 25848 1952 25900
rect 2004 25888 2010 25900
rect 2004 25860 5856 25888
rect 2004 25848 2010 25860
rect 5828 25820 5856 25860
rect 7282 25848 7288 25900
rect 7340 25888 7346 25900
rect 23198 25888 23204 25900
rect 7340 25860 12296 25888
rect 7340 25848 7346 25860
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 5828 25792 12173 25820
rect 12161 25789 12173 25792
rect 12207 25789 12219 25823
rect 12161 25783 12219 25789
rect 12069 25755 12127 25761
rect 12069 25752 12081 25755
rect 7576 25724 12081 25752
rect 842 25644 848 25696
rect 900 25684 906 25696
rect 7576 25684 7604 25724
rect 12069 25721 12081 25724
rect 12115 25721 12127 25755
rect 12268 25752 12296 25860
rect 17696 25860 23204 25888
rect 12437 25823 12495 25829
rect 12437 25789 12449 25823
rect 12483 25820 12495 25823
rect 14550 25820 14556 25832
rect 12483 25792 14556 25820
rect 12483 25789 12495 25792
rect 12437 25783 12495 25789
rect 14550 25780 14556 25792
rect 14608 25780 14614 25832
rect 14734 25780 14740 25832
rect 14792 25820 14798 25832
rect 17696 25820 17724 25860
rect 23198 25848 23204 25860
rect 23256 25848 23262 25900
rect 14792 25792 17724 25820
rect 17773 25823 17831 25829
rect 14792 25780 14798 25792
rect 17773 25789 17785 25823
rect 17819 25820 17831 25823
rect 23750 25820 23756 25832
rect 17819 25792 23756 25820
rect 17819 25789 17831 25792
rect 17773 25783 17831 25789
rect 23750 25780 23756 25792
rect 23808 25780 23814 25832
rect 18690 25752 18696 25764
rect 12268 25724 18696 25752
rect 12069 25715 12127 25721
rect 18690 25712 18696 25724
rect 18748 25712 18754 25764
rect 18782 25712 18788 25764
rect 18840 25752 18846 25764
rect 27614 25752 27620 25764
rect 18840 25724 27620 25752
rect 18840 25712 18846 25724
rect 27614 25712 27620 25724
rect 27672 25712 27678 25764
rect 900 25656 7604 25684
rect 7653 25687 7711 25693
rect 900 25644 906 25656
rect 7653 25653 7665 25687
rect 7699 25684 7711 25687
rect 9950 25684 9956 25696
rect 7699 25656 9956 25684
rect 7699 25653 7711 25656
rect 7653 25647 7711 25653
rect 9950 25644 9956 25656
rect 10008 25644 10014 25696
rect 11422 25644 11428 25696
rect 11480 25684 11486 25696
rect 22094 25684 22100 25696
rect 11480 25656 22100 25684
rect 11480 25644 11486 25656
rect 22094 25644 22100 25656
rect 22152 25644 22158 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 7653 25483 7711 25489
rect 7653 25449 7665 25483
rect 7699 25480 7711 25483
rect 7742 25480 7748 25492
rect 7699 25452 7748 25480
rect 7699 25449 7711 25452
rect 7653 25443 7711 25449
rect 7742 25440 7748 25452
rect 7800 25440 7806 25492
rect 8754 25480 8760 25492
rect 8715 25452 8760 25480
rect 8754 25440 8760 25452
rect 8812 25440 8818 25492
rect 10042 25480 10048 25492
rect 10003 25452 10048 25480
rect 10042 25440 10048 25452
rect 10100 25440 10106 25492
rect 11054 25440 11060 25492
rect 11112 25480 11118 25492
rect 11517 25483 11575 25489
rect 11517 25480 11529 25483
rect 11112 25452 11529 25480
rect 11112 25440 11118 25452
rect 11517 25449 11529 25452
rect 11563 25480 11575 25483
rect 13078 25480 13084 25492
rect 11563 25452 13084 25480
rect 11563 25449 11575 25452
rect 11517 25443 11575 25449
rect 13078 25440 13084 25452
rect 13136 25480 13142 25492
rect 14090 25480 14096 25492
rect 13136 25452 14096 25480
rect 13136 25440 13142 25452
rect 14090 25440 14096 25452
rect 14148 25440 14154 25492
rect 14461 25483 14519 25489
rect 14461 25449 14473 25483
rect 14507 25480 14519 25483
rect 14734 25480 14740 25492
rect 14507 25452 14740 25480
rect 14507 25449 14519 25452
rect 14461 25443 14519 25449
rect 14734 25440 14740 25452
rect 14792 25440 14798 25492
rect 14918 25480 14924 25492
rect 14879 25452 14924 25480
rect 14918 25440 14924 25452
rect 14976 25440 14982 25492
rect 15562 25440 15568 25492
rect 15620 25480 15626 25492
rect 18782 25480 18788 25492
rect 15620 25452 18788 25480
rect 15620 25440 15626 25452
rect 18782 25440 18788 25452
rect 18840 25440 18846 25492
rect 19705 25483 19763 25489
rect 19705 25449 19717 25483
rect 19751 25480 19763 25483
rect 20898 25480 20904 25492
rect 19751 25452 20904 25480
rect 19751 25449 19763 25452
rect 19705 25443 19763 25449
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 21913 25483 21971 25489
rect 21913 25449 21925 25483
rect 21959 25480 21971 25483
rect 24762 25480 24768 25492
rect 21959 25452 24768 25480
rect 21959 25449 21971 25452
rect 21913 25443 21971 25449
rect 24762 25440 24768 25452
rect 24820 25440 24826 25492
rect 6270 25372 6276 25424
rect 6328 25412 6334 25424
rect 10778 25412 10784 25424
rect 6328 25384 10784 25412
rect 6328 25372 6334 25384
rect 10778 25372 10784 25384
rect 10836 25372 10842 25424
rect 12437 25415 12495 25421
rect 12437 25381 12449 25415
rect 12483 25412 12495 25415
rect 13173 25415 13231 25421
rect 13173 25412 13185 25415
rect 12483 25384 13185 25412
rect 12483 25381 12495 25384
rect 12437 25375 12495 25381
rect 13173 25381 13185 25384
rect 13219 25412 13231 25415
rect 13262 25412 13268 25424
rect 13219 25384 13268 25412
rect 13219 25381 13231 25384
rect 13173 25375 13231 25381
rect 13262 25372 13268 25384
rect 13320 25372 13326 25424
rect 14826 25372 14832 25424
rect 14884 25412 14890 25424
rect 15838 25412 15844 25424
rect 14884 25384 15844 25412
rect 14884 25372 14890 25384
rect 15838 25372 15844 25384
rect 15896 25372 15902 25424
rect 16025 25415 16083 25421
rect 16025 25381 16037 25415
rect 16071 25381 16083 25415
rect 24854 25412 24860 25424
rect 16025 25375 16083 25381
rect 17052 25384 24860 25412
rect 7469 25347 7527 25353
rect 7469 25313 7481 25347
rect 7515 25344 7527 25347
rect 7742 25344 7748 25356
rect 7515 25316 7748 25344
rect 7515 25313 7527 25316
rect 7469 25307 7527 25313
rect 7742 25304 7748 25316
rect 7800 25304 7806 25356
rect 8573 25347 8631 25353
rect 8573 25313 8585 25347
rect 8619 25344 8631 25347
rect 9030 25344 9036 25356
rect 8619 25316 9036 25344
rect 8619 25313 8631 25316
rect 8573 25307 8631 25313
rect 9030 25304 9036 25316
rect 9088 25304 9094 25356
rect 9861 25347 9919 25353
rect 9861 25313 9873 25347
rect 9907 25344 9919 25347
rect 10962 25344 10968 25356
rect 9907 25316 10968 25344
rect 9907 25313 9919 25316
rect 9861 25307 9919 25313
rect 10962 25304 10968 25316
rect 11020 25304 11026 25356
rect 11330 25344 11336 25356
rect 11243 25316 11336 25344
rect 11330 25304 11336 25316
rect 11388 25344 11394 25356
rect 11790 25344 11796 25356
rect 11388 25316 11796 25344
rect 11388 25304 11394 25316
rect 11790 25304 11796 25316
rect 11848 25304 11854 25356
rect 12526 25304 12532 25356
rect 12584 25344 12590 25356
rect 12989 25347 13047 25353
rect 12989 25344 13001 25347
rect 12584 25316 13001 25344
rect 12584 25304 12590 25316
rect 12989 25313 13001 25316
rect 13035 25344 13047 25347
rect 13354 25344 13360 25356
rect 13035 25316 13360 25344
rect 13035 25313 13047 25316
rect 12989 25307 13047 25313
rect 13354 25304 13360 25316
rect 13412 25304 13418 25356
rect 14182 25304 14188 25356
rect 14240 25344 14246 25356
rect 14277 25347 14335 25353
rect 14277 25344 14289 25347
rect 14240 25316 14289 25344
rect 14240 25304 14246 25316
rect 14277 25313 14289 25316
rect 14323 25313 14335 25347
rect 14277 25307 14335 25313
rect 14366 25304 14372 25356
rect 14424 25344 14430 25356
rect 15470 25344 15476 25356
rect 14424 25316 15476 25344
rect 14424 25304 14430 25316
rect 15470 25304 15476 25316
rect 15528 25344 15534 25356
rect 16040 25344 16068 25375
rect 15528 25316 16068 25344
rect 15528 25304 15534 25316
rect 6454 25236 6460 25288
rect 6512 25276 6518 25288
rect 9585 25279 9643 25285
rect 6512 25248 9352 25276
rect 6512 25236 6518 25248
rect 8202 25168 8208 25220
rect 8260 25208 8266 25220
rect 9324 25208 9352 25248
rect 9585 25245 9597 25279
rect 9631 25276 9643 25279
rect 10042 25276 10048 25288
rect 9631 25248 10048 25276
rect 9631 25245 9643 25248
rect 9585 25239 9643 25245
rect 10042 25236 10048 25248
rect 10100 25236 10106 25288
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 10778 25276 10784 25288
rect 10551 25248 10784 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 10873 25279 10931 25285
rect 10873 25245 10885 25279
rect 10919 25276 10931 25279
rect 11609 25279 11667 25285
rect 11609 25276 11621 25279
rect 10919 25248 11621 25276
rect 10919 25245 10931 25248
rect 10873 25239 10931 25245
rect 11609 25245 11621 25248
rect 11655 25276 11667 25279
rect 12802 25276 12808 25288
rect 11655 25248 12808 25276
rect 11655 25245 11667 25248
rect 11609 25239 11667 25245
rect 12802 25236 12808 25248
rect 12860 25276 12866 25288
rect 13265 25279 13323 25285
rect 13265 25276 13277 25279
rect 12860 25248 13277 25276
rect 12860 25236 12866 25248
rect 13265 25245 13277 25248
rect 13311 25276 13323 25279
rect 15289 25279 15347 25285
rect 15289 25276 15301 25279
rect 13311 25248 15301 25276
rect 13311 25245 13323 25248
rect 13265 25239 13323 25245
rect 15289 25245 15301 25248
rect 15335 25276 15347 25279
rect 16117 25279 16175 25285
rect 16117 25276 16129 25279
rect 15335 25248 16129 25276
rect 15335 25245 15347 25248
rect 15289 25239 15347 25245
rect 16117 25245 16129 25248
rect 16163 25276 16175 25279
rect 16666 25276 16672 25288
rect 16163 25248 16672 25276
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 16666 25236 16672 25248
rect 16724 25236 16730 25288
rect 17052 25276 17080 25384
rect 24854 25372 24860 25384
rect 24912 25372 24918 25424
rect 17129 25347 17187 25353
rect 17129 25313 17141 25347
rect 17175 25344 17187 25347
rect 18417 25347 18475 25353
rect 17175 25316 17540 25344
rect 17175 25313 17187 25316
rect 17129 25307 17187 25313
rect 17052 25248 17356 25276
rect 8260 25180 9260 25208
rect 9324 25180 12848 25208
rect 8260 25168 8266 25180
rect 6638 25140 6644 25152
rect 6599 25112 6644 25140
rect 6638 25100 6644 25112
rect 6696 25100 6702 25152
rect 7377 25143 7435 25149
rect 7377 25109 7389 25143
rect 7423 25140 7435 25143
rect 7834 25140 7840 25152
rect 7423 25112 7840 25140
rect 7423 25109 7435 25112
rect 7377 25103 7435 25109
rect 7834 25100 7840 25112
rect 7892 25100 7898 25152
rect 8018 25140 8024 25152
rect 7979 25112 8024 25140
rect 8018 25100 8024 25112
rect 8076 25100 8082 25152
rect 8386 25140 8392 25152
rect 8347 25112 8392 25140
rect 8386 25100 8392 25112
rect 8444 25100 8450 25152
rect 9232 25149 9260 25180
rect 9217 25143 9275 25149
rect 9217 25109 9229 25143
rect 9263 25140 9275 25143
rect 9674 25140 9680 25152
rect 9263 25112 9680 25140
rect 9263 25109 9275 25112
rect 9217 25103 9275 25109
rect 9674 25100 9680 25112
rect 9732 25100 9738 25152
rect 11057 25143 11115 25149
rect 11057 25109 11069 25143
rect 11103 25140 11115 25143
rect 11977 25143 12035 25149
rect 11977 25140 11989 25143
rect 11103 25112 11989 25140
rect 11103 25109 11115 25112
rect 11057 25103 11115 25109
rect 11977 25109 11989 25112
rect 12023 25140 12035 25143
rect 12526 25140 12532 25152
rect 12023 25112 12532 25140
rect 12023 25109 12035 25112
rect 11977 25103 12035 25109
rect 12526 25100 12532 25112
rect 12584 25100 12590 25152
rect 12710 25140 12716 25152
rect 12671 25112 12716 25140
rect 12710 25100 12716 25112
rect 12768 25100 12774 25152
rect 12820 25140 12848 25180
rect 12986 25168 12992 25220
rect 13044 25208 13050 25220
rect 17328 25217 17356 25248
rect 17512 25220 17540 25316
rect 18417 25313 18429 25347
rect 18463 25344 18475 25347
rect 18506 25344 18512 25356
rect 18463 25316 18512 25344
rect 18463 25313 18475 25316
rect 18417 25307 18475 25313
rect 18506 25304 18512 25316
rect 18564 25304 18570 25356
rect 19518 25344 19524 25356
rect 19479 25316 19524 25344
rect 19518 25304 19524 25316
rect 19576 25304 19582 25356
rect 21266 25304 21272 25356
rect 21324 25344 21330 25356
rect 21729 25347 21787 25353
rect 21729 25344 21741 25347
rect 21324 25316 21741 25344
rect 21324 25304 21330 25316
rect 21729 25313 21741 25316
rect 21775 25313 21787 25347
rect 21729 25307 21787 25313
rect 22833 25347 22891 25353
rect 22833 25313 22845 25347
rect 22879 25344 22891 25347
rect 23014 25344 23020 25356
rect 22879 25316 23020 25344
rect 22879 25313 22891 25316
rect 22833 25307 22891 25313
rect 23014 25304 23020 25316
rect 23072 25304 23078 25356
rect 24118 25304 24124 25356
rect 24176 25344 24182 25356
rect 24581 25347 24639 25353
rect 24581 25344 24593 25347
rect 24176 25316 24593 25344
rect 24176 25304 24182 25316
rect 24581 25313 24593 25316
rect 24627 25313 24639 25347
rect 24581 25307 24639 25313
rect 25314 25276 25320 25288
rect 18616 25248 25320 25276
rect 13725 25211 13783 25217
rect 13725 25208 13737 25211
rect 13044 25180 13737 25208
rect 13044 25168 13050 25180
rect 13725 25177 13737 25180
rect 13771 25208 13783 25211
rect 15565 25211 15623 25217
rect 15565 25208 15577 25211
rect 13771 25180 15577 25208
rect 13771 25177 13783 25180
rect 13725 25171 13783 25177
rect 15565 25177 15577 25180
rect 15611 25177 15623 25211
rect 15565 25171 15623 25177
rect 17313 25211 17371 25217
rect 17313 25177 17325 25211
rect 17359 25177 17371 25211
rect 17313 25171 17371 25177
rect 17494 25168 17500 25220
rect 17552 25208 17558 25220
rect 18616 25217 18644 25248
rect 25314 25236 25320 25248
rect 25372 25236 25378 25288
rect 18601 25211 18659 25217
rect 17552 25180 18368 25208
rect 17552 25168 17558 25180
rect 13814 25140 13820 25152
rect 12820 25112 13820 25140
rect 13814 25100 13820 25112
rect 13872 25100 13878 25152
rect 13998 25140 14004 25152
rect 13959 25112 14004 25140
rect 13998 25100 14004 25112
rect 14056 25100 14062 25152
rect 14366 25100 14372 25152
rect 14424 25140 14430 25152
rect 16022 25140 16028 25152
rect 14424 25112 16028 25140
rect 14424 25100 14430 25112
rect 16022 25100 16028 25112
rect 16080 25100 16086 25152
rect 17865 25143 17923 25149
rect 17865 25109 17877 25143
rect 17911 25140 17923 25143
rect 18230 25140 18236 25152
rect 17911 25112 18236 25140
rect 17911 25109 17923 25112
rect 17865 25103 17923 25109
rect 18230 25100 18236 25112
rect 18288 25100 18294 25152
rect 18340 25140 18368 25180
rect 18601 25177 18613 25211
rect 18647 25177 18659 25211
rect 22370 25208 22376 25220
rect 18601 25171 18659 25177
rect 18708 25180 22376 25208
rect 18708 25140 18736 25180
rect 22370 25168 22376 25180
rect 22428 25168 22434 25220
rect 23017 25211 23075 25217
rect 23017 25177 23029 25211
rect 23063 25208 23075 25211
rect 24670 25208 24676 25220
rect 23063 25180 24676 25208
rect 23063 25177 23075 25180
rect 23017 25171 23075 25177
rect 24670 25168 24676 25180
rect 24728 25168 24734 25220
rect 18340 25112 18736 25140
rect 19426 25100 19432 25152
rect 19484 25140 19490 25152
rect 20070 25140 20076 25152
rect 19484 25112 20076 25140
rect 19484 25100 19490 25112
rect 20070 25100 20076 25112
rect 20128 25100 20134 25152
rect 20533 25143 20591 25149
rect 20533 25109 20545 25143
rect 20579 25140 20591 25143
rect 20622 25140 20628 25152
rect 20579 25112 20628 25140
rect 20579 25109 20591 25112
rect 20533 25103 20591 25109
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 21453 25143 21511 25149
rect 21453 25109 21465 25143
rect 21499 25140 21511 25143
rect 21634 25140 21640 25152
rect 21499 25112 21640 25140
rect 21499 25109 21511 25112
rect 21453 25103 21511 25109
rect 21634 25100 21640 25112
rect 21692 25100 21698 25152
rect 22278 25140 22284 25152
rect 22239 25112 22284 25140
rect 22278 25100 22284 25112
rect 22336 25100 22342 25152
rect 23658 25140 23664 25152
rect 23619 25112 23664 25140
rect 23658 25100 23664 25112
rect 23716 25100 23722 25152
rect 24762 25140 24768 25152
rect 24723 25112 24768 25140
rect 24762 25100 24768 25112
rect 24820 25100 24826 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 6086 24896 6092 24948
rect 6144 24936 6150 24948
rect 11422 24936 11428 24948
rect 6144 24908 11192 24936
rect 11383 24908 11428 24936
rect 6144 24896 6150 24908
rect 1670 24828 1676 24880
rect 1728 24868 1734 24880
rect 7377 24871 7435 24877
rect 7377 24868 7389 24871
rect 1728 24840 7389 24868
rect 1728 24828 1734 24840
rect 7377 24837 7389 24840
rect 7423 24868 7435 24871
rect 7653 24871 7711 24877
rect 7653 24868 7665 24871
rect 7423 24840 7665 24868
rect 7423 24837 7435 24840
rect 7377 24831 7435 24837
rect 7653 24837 7665 24840
rect 7699 24837 7711 24871
rect 7653 24831 7711 24837
rect 8938 24828 8944 24880
rect 8996 24868 9002 24880
rect 11054 24868 11060 24880
rect 8996 24840 10916 24868
rect 11015 24840 11060 24868
rect 8996 24828 9002 24840
rect 6914 24760 6920 24812
rect 6972 24800 6978 24812
rect 7745 24803 7803 24809
rect 7745 24800 7757 24803
rect 6972 24772 7757 24800
rect 6972 24760 6978 24772
rect 7745 24769 7757 24772
rect 7791 24800 7803 24803
rect 8389 24803 8447 24809
rect 8389 24800 8401 24803
rect 7791 24772 8401 24800
rect 7791 24769 7803 24772
rect 7745 24763 7803 24769
rect 8389 24769 8401 24772
rect 8435 24769 8447 24803
rect 10888 24800 10916 24840
rect 11054 24828 11060 24840
rect 11112 24828 11118 24880
rect 11164 24868 11192 24908
rect 11422 24896 11428 24908
rect 11480 24896 11486 24948
rect 15930 24936 15936 24948
rect 11532 24908 15936 24936
rect 11532 24868 11560 24908
rect 15930 24896 15936 24908
rect 15988 24896 15994 24948
rect 17494 24936 17500 24948
rect 17455 24908 17500 24936
rect 17494 24896 17500 24908
rect 17552 24896 17558 24948
rect 19978 24896 19984 24948
rect 20036 24936 20042 24948
rect 24210 24936 24216 24948
rect 20036 24908 24216 24936
rect 20036 24896 20042 24908
rect 24210 24896 24216 24908
rect 24268 24896 24274 24948
rect 11164 24840 11560 24868
rect 11790 24828 11796 24880
rect 11848 24868 11854 24880
rect 12253 24871 12311 24877
rect 12253 24868 12265 24871
rect 11848 24840 12265 24868
rect 11848 24828 11854 24840
rect 12253 24837 12265 24840
rect 12299 24868 12311 24871
rect 13630 24868 13636 24880
rect 12299 24840 13636 24868
rect 12299 24837 12311 24840
rect 12253 24831 12311 24837
rect 13630 24828 13636 24840
rect 13688 24828 13694 24880
rect 13814 24828 13820 24880
rect 13872 24868 13878 24880
rect 15562 24868 15568 24880
rect 13872 24840 15568 24868
rect 13872 24828 13878 24840
rect 15562 24828 15568 24840
rect 15620 24828 15626 24880
rect 15654 24828 15660 24880
rect 15712 24828 15718 24880
rect 16114 24828 16120 24880
rect 16172 24868 16178 24880
rect 20254 24868 20260 24880
rect 16172 24840 20260 24868
rect 16172 24828 16178 24840
rect 20254 24828 20260 24840
rect 20312 24868 20318 24880
rect 20312 24840 20484 24868
rect 20312 24828 20318 24840
rect 11330 24800 11336 24812
rect 10888 24772 11336 24800
rect 8389 24763 8447 24769
rect 11330 24760 11336 24772
rect 11388 24760 11394 24812
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24800 13047 24803
rect 13078 24800 13084 24812
rect 13035 24772 13084 24800
rect 13035 24769 13047 24772
rect 12989 24763 13047 24769
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 14090 24760 14096 24812
rect 14148 24800 14154 24812
rect 15197 24803 15255 24809
rect 15197 24800 15209 24803
rect 14148 24772 15209 24800
rect 14148 24760 14154 24772
rect 15197 24769 15209 24772
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 6641 24735 6699 24741
rect 6641 24701 6653 24735
rect 6687 24732 6699 24735
rect 6730 24732 6736 24744
rect 6687 24704 6736 24732
rect 6687 24701 6699 24704
rect 6641 24695 6699 24701
rect 6730 24692 6736 24704
rect 6788 24732 6794 24744
rect 6825 24735 6883 24741
rect 6825 24732 6837 24735
rect 6788 24704 6837 24732
rect 6788 24692 6794 24704
rect 6825 24701 6837 24704
rect 6871 24701 6883 24735
rect 6825 24695 6883 24701
rect 8018 24692 8024 24744
rect 8076 24732 8082 24744
rect 9401 24735 9459 24741
rect 8076 24704 8616 24732
rect 8076 24692 8082 24704
rect 6273 24667 6331 24673
rect 6273 24633 6285 24667
rect 6319 24664 6331 24667
rect 7098 24664 7104 24676
rect 6319 24636 7104 24664
rect 6319 24633 6331 24636
rect 6273 24627 6331 24633
rect 7098 24624 7104 24636
rect 7156 24624 7162 24676
rect 7653 24667 7711 24673
rect 7653 24633 7665 24667
rect 7699 24664 7711 24667
rect 8478 24664 8484 24676
rect 7699 24636 8484 24664
rect 7699 24633 7711 24636
rect 7653 24627 7711 24633
rect 8478 24624 8484 24636
rect 8536 24624 8542 24676
rect 8588 24673 8616 24704
rect 9401 24701 9413 24735
rect 9447 24732 9459 24735
rect 11241 24735 11299 24741
rect 9447 24704 10180 24732
rect 9447 24701 9459 24704
rect 9401 24695 9459 24701
rect 10152 24676 10180 24704
rect 11241 24701 11253 24735
rect 11287 24732 11299 24735
rect 13998 24732 14004 24744
rect 11287 24704 11652 24732
rect 13959 24704 14004 24732
rect 11287 24701 11299 24704
rect 11241 24695 11299 24701
rect 8573 24667 8631 24673
rect 8573 24633 8585 24667
rect 8619 24664 8631 24667
rect 8754 24664 8760 24676
rect 8619 24636 8760 24664
rect 8619 24633 8631 24636
rect 8573 24627 8631 24633
rect 8754 24624 8760 24636
rect 8812 24624 8818 24676
rect 9858 24664 9864 24676
rect 9819 24636 9864 24664
rect 9858 24624 9864 24636
rect 9916 24624 9922 24676
rect 10134 24664 10140 24676
rect 10095 24636 10140 24664
rect 10134 24624 10140 24636
rect 10192 24624 10198 24676
rect 11624 24608 11652 24704
rect 13998 24692 14004 24704
rect 14056 24692 14062 24744
rect 15212 24676 15240 24763
rect 15286 24760 15292 24812
rect 15344 24800 15350 24812
rect 15672 24800 15700 24828
rect 20456 24809 20484 24840
rect 23014 24828 23020 24880
rect 23072 24868 23078 24880
rect 25130 24868 25136 24880
rect 23072 24840 25136 24868
rect 23072 24828 23078 24840
rect 25130 24828 25136 24840
rect 25188 24828 25194 24880
rect 15344 24772 15700 24800
rect 20441 24803 20499 24809
rect 15344 24760 15350 24772
rect 20441 24769 20453 24803
rect 20487 24769 20499 24803
rect 22186 24800 22192 24812
rect 22099 24772 22192 24800
rect 20441 24763 20499 24769
rect 22186 24760 22192 24772
rect 22244 24800 22250 24812
rect 22649 24803 22707 24809
rect 22649 24800 22661 24803
rect 22244 24772 22661 24800
rect 22244 24760 22250 24772
rect 22649 24769 22661 24772
rect 22695 24769 22707 24803
rect 22649 24763 22707 24769
rect 15378 24692 15384 24744
rect 15436 24732 15442 24744
rect 15749 24735 15807 24741
rect 15749 24732 15761 24735
rect 15436 24704 15761 24732
rect 15436 24692 15442 24704
rect 15749 24701 15761 24704
rect 15795 24732 15807 24735
rect 16390 24732 16396 24744
rect 15795 24704 16396 24732
rect 15795 24701 15807 24704
rect 15749 24695 15807 24701
rect 16390 24692 16396 24704
rect 16448 24692 16454 24744
rect 18046 24692 18052 24744
rect 18104 24732 18110 24744
rect 18877 24735 18935 24741
rect 18877 24732 18889 24735
rect 18104 24704 18889 24732
rect 18104 24692 18110 24704
rect 18877 24701 18889 24704
rect 18923 24732 18935 24735
rect 19429 24735 19487 24741
rect 19429 24732 19441 24735
rect 18923 24704 19441 24732
rect 18923 24701 18935 24704
rect 18877 24695 18935 24701
rect 19429 24701 19441 24704
rect 19475 24701 19487 24735
rect 19429 24695 19487 24701
rect 20070 24692 20076 24744
rect 20128 24692 20134 24744
rect 23474 24692 23480 24744
rect 23532 24732 23538 24744
rect 24118 24732 24124 24744
rect 23532 24704 24124 24732
rect 23532 24692 23538 24704
rect 24118 24692 24124 24704
rect 24176 24692 24182 24744
rect 25038 24692 25044 24744
rect 25096 24732 25102 24744
rect 25225 24735 25283 24741
rect 25225 24732 25237 24735
rect 25096 24704 25237 24732
rect 25096 24692 25102 24704
rect 25225 24701 25237 24704
rect 25271 24732 25283 24735
rect 25777 24735 25835 24741
rect 25777 24732 25789 24735
rect 25271 24704 25789 24732
rect 25271 24701 25283 24704
rect 25225 24695 25283 24701
rect 25777 24701 25789 24704
rect 25823 24701 25835 24735
rect 25777 24695 25835 24701
rect 12986 24664 12992 24676
rect 12947 24636 12992 24664
rect 12986 24624 12992 24636
rect 13044 24624 13050 24676
rect 13078 24624 13084 24676
rect 13136 24664 13142 24676
rect 13817 24667 13875 24673
rect 13817 24664 13829 24667
rect 13136 24636 13829 24664
rect 13136 24624 13142 24636
rect 13817 24633 13829 24636
rect 13863 24633 13875 24667
rect 14274 24664 14280 24676
rect 14235 24636 14280 24664
rect 13817 24627 13875 24633
rect 14274 24624 14280 24636
rect 14332 24624 14338 24676
rect 15194 24664 15200 24676
rect 15107 24636 15200 24664
rect 15194 24624 15200 24636
rect 15252 24664 15258 24676
rect 15933 24667 15991 24673
rect 15933 24664 15945 24667
rect 15252 24636 15945 24664
rect 15252 24624 15258 24636
rect 15933 24633 15945 24636
rect 15979 24633 15991 24667
rect 15933 24627 15991 24633
rect 16025 24667 16083 24673
rect 16025 24633 16037 24667
rect 16071 24664 16083 24667
rect 16761 24667 16819 24673
rect 16761 24664 16773 24667
rect 16071 24636 16773 24664
rect 16071 24633 16083 24636
rect 16025 24627 16083 24633
rect 16761 24633 16773 24636
rect 16807 24664 16819 24667
rect 16850 24664 16856 24676
rect 16807 24636 16856 24664
rect 16807 24633 16819 24636
rect 16761 24627 16819 24633
rect 16850 24624 16856 24636
rect 16908 24624 16914 24676
rect 16945 24667 17003 24673
rect 16945 24633 16957 24667
rect 16991 24664 17003 24667
rect 17862 24664 17868 24676
rect 16991 24636 17868 24664
rect 16991 24633 17003 24636
rect 16945 24627 17003 24633
rect 17862 24624 17868 24636
rect 17920 24624 17926 24676
rect 20088 24664 20116 24692
rect 20622 24664 20628 24676
rect 20088 24636 20300 24664
rect 20583 24636 20628 24664
rect 4706 24556 4712 24608
rect 4764 24596 4770 24608
rect 4801 24599 4859 24605
rect 4801 24596 4813 24599
rect 4764 24568 4813 24596
rect 4764 24556 4770 24568
rect 4801 24565 4813 24568
rect 4847 24565 4859 24599
rect 5258 24596 5264 24608
rect 5219 24568 5264 24596
rect 4801 24559 4859 24565
rect 5258 24556 5264 24568
rect 5316 24556 5322 24608
rect 5534 24596 5540 24608
rect 5495 24568 5540 24596
rect 5534 24556 5540 24568
rect 5592 24556 5598 24608
rect 7006 24596 7012 24608
rect 6967 24568 7012 24596
rect 7006 24556 7012 24568
rect 7064 24556 7070 24608
rect 7466 24556 7472 24608
rect 7524 24596 7530 24608
rect 8003 24599 8061 24605
rect 8003 24596 8015 24599
rect 7524 24568 8015 24596
rect 7524 24556 7530 24568
rect 8003 24565 8015 24568
rect 8049 24565 8061 24599
rect 9030 24596 9036 24608
rect 8991 24568 9036 24596
rect 8003 24559 8061 24565
rect 9030 24556 9036 24568
rect 9088 24556 9094 24608
rect 9582 24605 9588 24608
rect 9575 24599 9588 24605
rect 9575 24565 9587 24599
rect 9640 24596 9646 24608
rect 10042 24596 10048 24608
rect 9640 24568 9675 24596
rect 10003 24568 10048 24596
rect 9575 24559 9588 24565
rect 9582 24556 9588 24559
rect 9640 24556 9646 24568
rect 10042 24556 10048 24568
rect 10100 24556 10106 24608
rect 10597 24599 10655 24605
rect 10597 24565 10609 24599
rect 10643 24596 10655 24599
rect 10962 24596 10968 24608
rect 10643 24568 10968 24596
rect 10643 24565 10655 24568
rect 10597 24559 10655 24565
rect 10962 24556 10968 24568
rect 11020 24556 11026 24608
rect 11606 24556 11612 24608
rect 11664 24596 11670 24608
rect 12526 24605 12532 24608
rect 11793 24599 11851 24605
rect 11793 24596 11805 24599
rect 11664 24568 11805 24596
rect 11664 24556 11670 24568
rect 11793 24565 11805 24568
rect 11839 24565 11851 24599
rect 11793 24559 11851 24565
rect 12519 24599 12532 24605
rect 12519 24565 12531 24599
rect 12584 24596 12590 24608
rect 12584 24568 12619 24596
rect 12519 24559 12532 24565
rect 12526 24556 12532 24559
rect 12584 24556 12590 24568
rect 13354 24556 13360 24608
rect 13412 24596 13418 24608
rect 13449 24599 13507 24605
rect 13449 24596 13461 24599
rect 13412 24568 13461 24596
rect 13412 24556 13418 24568
rect 13449 24565 13461 24568
rect 13495 24565 13507 24599
rect 13449 24559 13507 24565
rect 14182 24556 14188 24608
rect 14240 24596 14246 24608
rect 14737 24599 14795 24605
rect 14737 24596 14749 24599
rect 14240 24568 14749 24596
rect 14240 24556 14246 24568
rect 14737 24565 14749 24568
rect 14783 24565 14795 24599
rect 14737 24559 14795 24565
rect 15463 24599 15521 24605
rect 15463 24565 15475 24599
rect 15509 24596 15521 24599
rect 15654 24596 15660 24608
rect 15509 24568 15660 24596
rect 15509 24565 15521 24568
rect 15463 24559 15521 24565
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 17773 24599 17831 24605
rect 17773 24565 17785 24599
rect 17819 24596 17831 24599
rect 18322 24596 18328 24608
rect 17819 24568 18328 24596
rect 17819 24565 17831 24568
rect 17773 24559 17831 24565
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 18506 24596 18512 24608
rect 18467 24568 18512 24596
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 19058 24596 19064 24608
rect 19019 24568 19064 24596
rect 19058 24556 19064 24568
rect 19116 24556 19122 24608
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 20070 24605 20076 24608
rect 19797 24599 19855 24605
rect 19797 24596 19809 24599
rect 19484 24568 19809 24596
rect 19484 24556 19490 24568
rect 19797 24565 19809 24568
rect 19843 24565 19855 24599
rect 19797 24559 19855 24565
rect 20063 24599 20076 24605
rect 20063 24565 20075 24599
rect 20128 24596 20134 24608
rect 20272 24596 20300 24636
rect 20622 24624 20628 24636
rect 20680 24624 20686 24676
rect 21177 24667 21235 24673
rect 21177 24633 21189 24667
rect 21223 24664 21235 24667
rect 21711 24667 21769 24673
rect 21223 24636 21680 24664
rect 21223 24633 21235 24636
rect 21177 24627 21235 24633
rect 20533 24599 20591 24605
rect 20533 24596 20545 24599
rect 20128 24568 20163 24596
rect 20272 24568 20545 24596
rect 20063 24559 20076 24565
rect 20070 24556 20076 24559
rect 20128 24556 20134 24568
rect 20533 24565 20545 24568
rect 20579 24565 20591 24599
rect 20533 24559 20591 24565
rect 21266 24556 21272 24608
rect 21324 24596 21330 24608
rect 21453 24599 21511 24605
rect 21453 24596 21465 24599
rect 21324 24568 21465 24596
rect 21324 24556 21330 24568
rect 21453 24565 21465 24568
rect 21499 24565 21511 24599
rect 21652 24596 21680 24636
rect 21711 24633 21723 24667
rect 21757 24664 21769 24667
rect 22002 24664 22008 24676
rect 21757 24636 22008 24664
rect 21757 24633 21769 24636
rect 21711 24627 21769 24633
rect 22002 24624 22008 24636
rect 22060 24624 22066 24676
rect 22278 24664 22284 24676
rect 22239 24636 22284 24664
rect 22278 24624 22284 24636
rect 22336 24624 22342 24676
rect 22922 24624 22928 24676
rect 22980 24664 22986 24676
rect 23658 24664 23664 24676
rect 22980 24636 23664 24664
rect 22980 24624 22986 24636
rect 23658 24624 23664 24636
rect 23716 24664 23722 24676
rect 24029 24667 24087 24673
rect 24029 24664 24041 24667
rect 23716 24636 24041 24664
rect 23716 24624 23722 24636
rect 24029 24633 24041 24636
rect 24075 24633 24087 24667
rect 24029 24627 24087 24633
rect 21818 24596 21824 24608
rect 21652 24568 21824 24596
rect 21453 24559 21511 24565
rect 21818 24556 21824 24568
rect 21876 24596 21882 24608
rect 22189 24599 22247 24605
rect 22189 24596 22201 24599
rect 21876 24568 22201 24596
rect 21876 24556 21882 24568
rect 22189 24565 22201 24568
rect 22235 24565 22247 24599
rect 22296 24596 22324 24624
rect 23017 24599 23075 24605
rect 23017 24596 23029 24599
rect 22296 24568 23029 24596
rect 22189 24559 22247 24565
rect 23017 24565 23029 24568
rect 23063 24596 23075 24599
rect 23290 24596 23296 24608
rect 23063 24568 23296 24596
rect 23063 24565 23075 24568
rect 23017 24559 23075 24565
rect 23290 24556 23296 24568
rect 23348 24556 23354 24608
rect 23474 24596 23480 24608
rect 23435 24568 23480 24596
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 23750 24605 23756 24608
rect 23743 24599 23756 24605
rect 23743 24565 23755 24599
rect 23808 24596 23814 24608
rect 24136 24596 24164 24692
rect 24302 24664 24308 24676
rect 24263 24636 24308 24664
rect 24302 24624 24308 24636
rect 24360 24624 24366 24676
rect 24213 24599 24271 24605
rect 24213 24596 24225 24599
rect 23808 24568 23843 24596
rect 24136 24568 24225 24596
rect 23743 24559 23756 24565
rect 23750 24556 23756 24559
rect 23808 24556 23814 24568
rect 24213 24565 24225 24568
rect 24259 24596 24271 24599
rect 24673 24599 24731 24605
rect 24673 24596 24685 24599
rect 24259 24568 24685 24596
rect 24259 24565 24271 24568
rect 24213 24559 24271 24565
rect 24673 24565 24685 24568
rect 24719 24565 24731 24599
rect 25406 24596 25412 24608
rect 25367 24568 25412 24596
rect 24673 24559 24731 24565
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1578 24392 1584 24404
rect 1539 24364 1584 24392
rect 1578 24352 1584 24364
rect 1636 24352 1642 24404
rect 5997 24395 6055 24401
rect 5997 24361 6009 24395
rect 6043 24392 6055 24395
rect 6086 24392 6092 24404
rect 6043 24364 6092 24392
rect 6043 24361 6055 24364
rect 5997 24355 6055 24361
rect 6086 24352 6092 24364
rect 6144 24352 6150 24404
rect 6454 24392 6460 24404
rect 6415 24364 6460 24392
rect 6454 24352 6460 24364
rect 6512 24352 6518 24404
rect 7101 24395 7159 24401
rect 7101 24361 7113 24395
rect 7147 24392 7159 24395
rect 7282 24392 7288 24404
rect 7147 24364 7288 24392
rect 7147 24361 7159 24364
rect 7101 24355 7159 24361
rect 7282 24352 7288 24364
rect 7340 24352 7346 24404
rect 10505 24395 10563 24401
rect 10505 24361 10517 24395
rect 10551 24392 10563 24395
rect 11238 24392 11244 24404
rect 10551 24364 11244 24392
rect 10551 24361 10563 24364
rect 10505 24355 10563 24361
rect 11238 24352 11244 24364
rect 11296 24392 11302 24404
rect 12526 24392 12532 24404
rect 11296 24364 12532 24392
rect 11296 24352 11302 24364
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 12710 24352 12716 24404
rect 12768 24392 12774 24404
rect 14921 24395 14979 24401
rect 14921 24392 14933 24395
rect 12768 24364 14933 24392
rect 12768 24352 12774 24364
rect 14921 24361 14933 24364
rect 14967 24361 14979 24395
rect 15470 24392 15476 24404
rect 15431 24364 15476 24392
rect 14921 24355 14979 24361
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 15838 24392 15844 24404
rect 15799 24364 15844 24392
rect 15838 24352 15844 24364
rect 15896 24392 15902 24404
rect 16114 24392 16120 24404
rect 15896 24364 16120 24392
rect 15896 24352 15902 24364
rect 16114 24352 16120 24364
rect 16172 24352 16178 24404
rect 16850 24352 16856 24404
rect 16908 24392 16914 24404
rect 18782 24392 18788 24404
rect 16908 24364 18788 24392
rect 16908 24352 16914 24364
rect 18782 24352 18788 24364
rect 18840 24352 18846 24404
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 19978 24392 19984 24404
rect 19935 24364 19984 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 20254 24392 20260 24404
rect 20215 24364 20260 24392
rect 20254 24352 20260 24364
rect 20312 24352 20318 24404
rect 22925 24395 22983 24401
rect 22925 24361 22937 24395
rect 22971 24392 22983 24395
rect 23014 24392 23020 24404
rect 22971 24364 23020 24392
rect 22971 24361 22983 24364
rect 22925 24355 22983 24361
rect 23014 24352 23020 24364
rect 23072 24352 23078 24404
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 2222 24256 2228 24268
rect 1443 24228 2228 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 2222 24216 2228 24228
rect 2280 24216 2286 24268
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6472 24256 6500 24352
rect 8573 24327 8631 24333
rect 8573 24293 8585 24327
rect 8619 24324 8631 24327
rect 8846 24324 8852 24336
rect 8619 24296 8852 24324
rect 8619 24293 8631 24296
rect 8573 24287 8631 24293
rect 8846 24284 8852 24296
rect 8904 24284 8910 24336
rect 13446 24284 13452 24336
rect 13504 24324 13510 24336
rect 13725 24327 13783 24333
rect 13725 24324 13737 24327
rect 13504 24296 13737 24324
rect 13504 24284 13510 24296
rect 13725 24293 13737 24296
rect 13771 24293 13783 24327
rect 13725 24287 13783 24293
rect 16761 24327 16819 24333
rect 16761 24293 16773 24327
rect 16807 24324 16819 24327
rect 16942 24324 16948 24336
rect 16807 24296 16948 24324
rect 16807 24293 16819 24296
rect 16761 24287 16819 24293
rect 16942 24284 16948 24296
rect 17000 24324 17006 24336
rect 17221 24327 17279 24333
rect 17221 24324 17233 24327
rect 17000 24296 17233 24324
rect 17000 24284 17006 24296
rect 17221 24293 17233 24296
rect 17267 24293 17279 24327
rect 18322 24324 18328 24336
rect 18283 24296 18328 24324
rect 17221 24287 17279 24293
rect 18322 24284 18328 24296
rect 18380 24284 18386 24336
rect 21082 24284 21088 24336
rect 21140 24324 21146 24336
rect 22005 24327 22063 24333
rect 22005 24324 22017 24327
rect 21140 24296 22017 24324
rect 21140 24284 21146 24296
rect 22005 24293 22017 24296
rect 22051 24293 22063 24327
rect 22005 24287 22063 24293
rect 22830 24284 22836 24336
rect 22888 24324 22894 24336
rect 23661 24327 23719 24333
rect 23661 24324 23673 24327
rect 22888 24296 23673 24324
rect 22888 24284 22894 24296
rect 23661 24293 23673 24296
rect 23707 24293 23719 24327
rect 23661 24287 23719 24293
rect 6914 24256 6920 24268
rect 5859 24228 6500 24256
rect 6875 24228 6920 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 6914 24216 6920 24228
rect 6972 24216 6978 24268
rect 7742 24216 7748 24268
rect 7800 24256 7806 24268
rect 7929 24259 7987 24265
rect 7929 24256 7941 24259
rect 7800 24228 7941 24256
rect 7800 24216 7806 24228
rect 7929 24225 7941 24228
rect 7975 24256 7987 24259
rect 8018 24256 8024 24268
rect 7975 24228 8024 24256
rect 7975 24225 7987 24228
rect 7929 24219 7987 24225
rect 8018 24216 8024 24228
rect 8076 24216 8082 24268
rect 8294 24216 8300 24268
rect 8352 24256 8358 24268
rect 8389 24259 8447 24265
rect 8389 24256 8401 24259
rect 8352 24228 8401 24256
rect 8352 24216 8358 24228
rect 8389 24225 8401 24228
rect 8435 24225 8447 24259
rect 10864 24259 10922 24265
rect 10864 24256 10876 24259
rect 8389 24219 8447 24225
rect 10428 24228 10876 24256
rect 4525 24191 4583 24197
rect 4525 24157 4537 24191
rect 4571 24188 4583 24191
rect 5166 24188 5172 24200
rect 4571 24160 5172 24188
rect 4571 24157 4583 24160
rect 4525 24151 4583 24157
rect 5166 24148 5172 24160
rect 5224 24148 5230 24200
rect 5261 24191 5319 24197
rect 5261 24157 5273 24191
rect 5307 24188 5319 24191
rect 6178 24188 6184 24200
rect 5307 24160 6184 24188
rect 5307 24157 5319 24160
rect 5261 24151 5319 24157
rect 6178 24148 6184 24160
rect 6236 24148 6242 24200
rect 8665 24191 8723 24197
rect 8665 24188 8677 24191
rect 7760 24160 8677 24188
rect 4893 24123 4951 24129
rect 4893 24089 4905 24123
rect 4939 24120 4951 24123
rect 5350 24120 5356 24132
rect 4939 24092 5356 24120
rect 4939 24089 4951 24092
rect 4893 24083 4951 24089
rect 5350 24080 5356 24092
rect 5408 24080 5414 24132
rect 7760 24064 7788 24160
rect 8665 24157 8677 24160
rect 8711 24188 8723 24191
rect 10428 24188 10456 24228
rect 10864 24225 10876 24228
rect 10910 24256 10922 24259
rect 11422 24256 11428 24268
rect 10910 24228 11428 24256
rect 10910 24225 10922 24228
rect 10864 24219 10922 24225
rect 11422 24216 11428 24228
rect 11480 24216 11486 24268
rect 11974 24216 11980 24268
rect 12032 24256 12038 24268
rect 13541 24259 13599 24265
rect 13541 24256 13553 24259
rect 12032 24228 13553 24256
rect 12032 24216 12038 24228
rect 10594 24188 10600 24200
rect 8711 24160 10456 24188
rect 10555 24160 10600 24188
rect 8711 24157 8723 24160
rect 8665 24151 8723 24157
rect 10594 24148 10600 24160
rect 10652 24148 10658 24200
rect 12434 24148 12440 24200
rect 12492 24188 12498 24200
rect 12894 24188 12900 24200
rect 12492 24160 12900 24188
rect 12492 24148 12498 24160
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 8113 24123 8171 24129
rect 8113 24089 8125 24123
rect 8159 24120 8171 24123
rect 8202 24120 8208 24132
rect 8159 24092 8208 24120
rect 8159 24089 8171 24092
rect 8113 24083 8171 24089
rect 8202 24080 8208 24092
rect 8260 24080 8266 24132
rect 12713 24123 12771 24129
rect 12713 24089 12725 24123
rect 12759 24120 12771 24123
rect 12802 24120 12808 24132
rect 12759 24092 12808 24120
rect 12759 24089 12771 24092
rect 12713 24083 12771 24089
rect 12802 24080 12808 24092
rect 12860 24080 12866 24132
rect 13262 24120 13268 24132
rect 13223 24092 13268 24120
rect 13262 24080 13268 24092
rect 13320 24080 13326 24132
rect 13464 24120 13492 24228
rect 13541 24225 13553 24228
rect 13587 24225 13599 24259
rect 14550 24256 14556 24268
rect 14511 24228 14556 24256
rect 13541 24219 13599 24225
rect 14550 24216 14556 24228
rect 14608 24216 14614 24268
rect 16574 24216 16580 24268
rect 16632 24256 16638 24268
rect 16853 24259 16911 24265
rect 16853 24256 16865 24259
rect 16632 24228 16865 24256
rect 16632 24216 16638 24228
rect 16853 24225 16865 24228
rect 16899 24225 16911 24259
rect 19702 24256 19708 24268
rect 19663 24228 19708 24256
rect 16853 24219 16911 24225
rect 19702 24216 19708 24228
rect 19760 24216 19766 24268
rect 23290 24216 23296 24268
rect 23348 24256 23354 24268
rect 23753 24259 23811 24265
rect 23753 24256 23765 24259
rect 23348 24228 23765 24256
rect 23348 24216 23354 24228
rect 23753 24225 23765 24228
rect 23799 24256 23811 24259
rect 24302 24256 24308 24268
rect 23799 24228 24308 24256
rect 23799 24225 23811 24228
rect 23753 24219 23811 24225
rect 24302 24216 24308 24228
rect 24360 24256 24366 24268
rect 24489 24259 24547 24265
rect 24489 24256 24501 24259
rect 24360 24228 24501 24256
rect 24360 24216 24366 24228
rect 24489 24225 24501 24228
rect 24535 24225 24547 24259
rect 24489 24219 24547 24225
rect 24673 24259 24731 24265
rect 24673 24225 24685 24259
rect 24719 24256 24731 24259
rect 24946 24256 24952 24268
rect 24719 24228 24952 24256
rect 24719 24225 24731 24228
rect 24673 24219 24731 24225
rect 24946 24216 24952 24228
rect 25004 24216 25010 24268
rect 13817 24191 13875 24197
rect 13817 24157 13829 24191
rect 13863 24157 13875 24191
rect 13817 24151 13875 24157
rect 13538 24120 13544 24132
rect 13464 24092 13544 24120
rect 13538 24080 13544 24092
rect 13596 24080 13602 24132
rect 13832 24120 13860 24151
rect 16206 24148 16212 24200
rect 16264 24188 16270 24200
rect 16669 24191 16727 24197
rect 16669 24188 16681 24191
rect 16264 24160 16681 24188
rect 16264 24148 16270 24160
rect 16669 24157 16681 24160
rect 16715 24188 16727 24191
rect 18046 24188 18052 24200
rect 16715 24160 18052 24188
rect 16715 24157 16727 24160
rect 16669 24151 16727 24157
rect 18046 24148 18052 24160
rect 18104 24148 18110 24200
rect 18230 24188 18236 24200
rect 18143 24160 18236 24188
rect 18230 24148 18236 24160
rect 18288 24148 18294 24200
rect 18414 24188 18420 24200
rect 18375 24160 18420 24188
rect 18414 24148 18420 24160
rect 18472 24148 18478 24200
rect 21910 24188 21916 24200
rect 21871 24160 21916 24188
rect 21910 24148 21916 24160
rect 21968 24148 21974 24200
rect 22094 24148 22100 24200
rect 22152 24188 22158 24200
rect 22152 24160 22197 24188
rect 22152 24148 22158 24160
rect 23382 24148 23388 24200
rect 23440 24188 23446 24200
rect 23569 24191 23627 24197
rect 23569 24188 23581 24191
rect 23440 24160 23581 24188
rect 23440 24148 23446 24160
rect 23569 24157 23581 24160
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 14277 24123 14335 24129
rect 14277 24120 14289 24123
rect 13832 24092 14289 24120
rect 5721 24055 5779 24061
rect 5721 24021 5733 24055
rect 5767 24052 5779 24055
rect 6546 24052 6552 24064
rect 5767 24024 6552 24052
rect 5767 24021 5779 24024
rect 5721 24015 5779 24021
rect 6546 24012 6552 24024
rect 6604 24012 6610 24064
rect 6822 24052 6828 24064
rect 6783 24024 6828 24052
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 7561 24055 7619 24061
rect 7561 24021 7573 24055
rect 7607 24052 7619 24055
rect 7742 24052 7748 24064
rect 7607 24024 7748 24052
rect 7607 24021 7619 24024
rect 7561 24015 7619 24021
rect 7742 24012 7748 24024
rect 7800 24012 7806 24064
rect 9122 24052 9128 24064
rect 9083 24024 9128 24052
rect 9122 24012 9128 24024
rect 9180 24012 9186 24064
rect 9490 24052 9496 24064
rect 9451 24024 9496 24052
rect 9490 24012 9496 24024
rect 9548 24012 9554 24064
rect 9858 24052 9864 24064
rect 9819 24024 9864 24052
rect 9858 24012 9864 24024
rect 9916 24012 9922 24064
rect 11974 24052 11980 24064
rect 11935 24024 11980 24052
rect 11974 24012 11980 24024
rect 12032 24012 12038 24064
rect 13081 24055 13139 24061
rect 13081 24021 13093 24055
rect 13127 24052 13139 24055
rect 13832 24052 13860 24092
rect 14277 24089 14289 24092
rect 14323 24120 14335 24123
rect 14734 24120 14740 24132
rect 14323 24092 14740 24120
rect 14323 24089 14335 24092
rect 14277 24083 14335 24089
rect 14734 24080 14740 24092
rect 14792 24080 14798 24132
rect 18248 24120 18276 24148
rect 18690 24120 18696 24132
rect 18248 24092 18696 24120
rect 18690 24080 18696 24092
rect 18748 24080 18754 24132
rect 21361 24123 21419 24129
rect 21361 24089 21373 24123
rect 21407 24120 21419 24123
rect 21818 24120 21824 24132
rect 21407 24092 21824 24120
rect 21407 24089 21419 24092
rect 21361 24083 21419 24089
rect 21818 24080 21824 24092
rect 21876 24080 21882 24132
rect 16298 24052 16304 24064
rect 13127 24024 13860 24052
rect 16259 24024 16304 24052
rect 13127 24021 13139 24024
rect 13081 24015 13139 24021
rect 16298 24012 16304 24024
rect 16356 24012 16362 24064
rect 17586 24052 17592 24064
rect 17547 24024 17592 24052
rect 17586 24012 17592 24024
rect 17644 24012 17650 24064
rect 17865 24055 17923 24061
rect 17865 24021 17877 24055
rect 17911 24052 17923 24055
rect 18230 24052 18236 24064
rect 17911 24024 18236 24052
rect 17911 24021 17923 24024
rect 17865 24015 17923 24021
rect 18230 24012 18236 24024
rect 18288 24012 18294 24064
rect 19150 24052 19156 24064
rect 19111 24024 19156 24052
rect 19150 24012 19156 24024
rect 19208 24012 19214 24064
rect 19518 24052 19524 24064
rect 19479 24024 19524 24052
rect 19518 24012 19524 24024
rect 19576 24012 19582 24064
rect 20714 24052 20720 24064
rect 20675 24024 20720 24052
rect 20714 24012 20720 24024
rect 20772 24012 20778 24064
rect 21542 24052 21548 24064
rect 21503 24024 21548 24052
rect 21542 24012 21548 24024
rect 21600 24012 21606 24064
rect 22554 24052 22560 24064
rect 22515 24024 22560 24052
rect 22554 24012 22560 24024
rect 22612 24012 22618 24064
rect 23198 24052 23204 24064
rect 23159 24024 23204 24052
rect 23198 24012 23204 24024
rect 23256 24012 23262 24064
rect 24118 24052 24124 24064
rect 24079 24024 24124 24052
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 24762 24012 24768 24064
rect 24820 24052 24826 24064
rect 24857 24055 24915 24061
rect 24857 24052 24869 24055
rect 24820 24024 24869 24052
rect 24820 24012 24826 24024
rect 24857 24021 24869 24024
rect 24903 24021 24915 24055
rect 24857 24015 24915 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1394 23808 1400 23860
rect 1452 23848 1458 23860
rect 1581 23851 1639 23857
rect 1581 23848 1593 23851
rect 1452 23820 1593 23848
rect 1452 23808 1458 23820
rect 1581 23817 1593 23820
rect 1627 23817 1639 23851
rect 1581 23811 1639 23817
rect 5813 23851 5871 23857
rect 5813 23817 5825 23851
rect 5859 23848 5871 23851
rect 6270 23848 6276 23860
rect 5859 23820 6276 23848
rect 5859 23817 5871 23820
rect 5813 23811 5871 23817
rect 6270 23808 6276 23820
rect 6328 23808 6334 23860
rect 7558 23848 7564 23860
rect 7519 23820 7564 23848
rect 7558 23808 7564 23820
rect 7616 23808 7622 23860
rect 8202 23808 8208 23860
rect 8260 23848 8266 23860
rect 9030 23848 9036 23860
rect 8260 23820 9036 23848
rect 8260 23808 8266 23820
rect 9030 23808 9036 23820
rect 9088 23848 9094 23860
rect 12342 23848 12348 23860
rect 9088 23820 12348 23848
rect 9088 23808 9094 23820
rect 12342 23808 12348 23820
rect 12400 23808 12406 23860
rect 12526 23848 12532 23860
rect 12487 23820 12532 23848
rect 12526 23808 12532 23820
rect 12584 23808 12590 23860
rect 14550 23808 14556 23860
rect 14608 23848 14614 23860
rect 15565 23851 15623 23857
rect 14608 23820 15148 23848
rect 14608 23808 14614 23820
rect 11422 23780 11428 23792
rect 11335 23752 11428 23780
rect 11422 23740 11428 23752
rect 11480 23780 11486 23792
rect 12802 23780 12808 23792
rect 11480 23752 12808 23780
rect 11480 23740 11486 23752
rect 12802 23740 12808 23752
rect 12860 23740 12866 23792
rect 15120 23780 15148 23820
rect 15565 23817 15577 23851
rect 15611 23848 15623 23851
rect 15746 23848 15752 23860
rect 15611 23820 15752 23848
rect 15611 23817 15623 23820
rect 15565 23811 15623 23817
rect 15746 23808 15752 23820
rect 15804 23808 15810 23860
rect 18138 23848 18144 23860
rect 18099 23820 18144 23848
rect 18138 23808 18144 23820
rect 18196 23808 18202 23860
rect 18966 23808 18972 23860
rect 19024 23848 19030 23860
rect 19153 23851 19211 23857
rect 19153 23848 19165 23851
rect 19024 23820 19165 23848
rect 19024 23808 19030 23820
rect 19153 23817 19165 23820
rect 19199 23817 19211 23851
rect 19613 23851 19671 23857
rect 19613 23848 19625 23851
rect 19153 23811 19211 23817
rect 19260 23820 19625 23848
rect 15120 23752 18920 23780
rect 7377 23715 7435 23721
rect 7377 23681 7389 23715
rect 7423 23712 7435 23715
rect 8018 23712 8024 23724
rect 7423 23684 8024 23712
rect 7423 23681 7435 23684
rect 7377 23675 7435 23681
rect 8018 23672 8024 23684
rect 8076 23672 8082 23724
rect 11974 23672 11980 23724
rect 12032 23712 12038 23724
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 12032 23684 12081 23712
rect 12032 23672 12038 23684
rect 12069 23681 12081 23684
rect 12115 23712 12127 23715
rect 13078 23712 13084 23724
rect 12115 23684 13084 23712
rect 12115 23681 12127 23684
rect 12069 23675 12127 23681
rect 13078 23672 13084 23684
rect 13136 23672 13142 23724
rect 17497 23715 17555 23721
rect 17497 23681 17509 23715
rect 17543 23712 17555 23715
rect 18414 23712 18420 23724
rect 17543 23684 18420 23712
rect 17543 23681 17555 23684
rect 17497 23675 17555 23681
rect 18414 23672 18420 23684
rect 18472 23672 18478 23724
rect 18693 23715 18751 23721
rect 18693 23681 18705 23715
rect 18739 23712 18751 23715
rect 18782 23712 18788 23724
rect 18739 23684 18788 23712
rect 18739 23681 18751 23684
rect 18693 23675 18751 23681
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 1443 23616 2452 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 2424 23520 2452 23616
rect 4614 23604 4620 23656
rect 4672 23644 4678 23656
rect 5077 23647 5135 23653
rect 5077 23644 5089 23647
rect 4672 23616 5089 23644
rect 4672 23604 4678 23616
rect 5077 23613 5089 23616
rect 5123 23613 5135 23647
rect 5077 23607 5135 23613
rect 5629 23647 5687 23653
rect 5629 23613 5641 23647
rect 5675 23644 5687 23647
rect 9030 23644 9036 23656
rect 5675 23616 6408 23644
rect 8991 23616 9036 23644
rect 5675 23613 5687 23616
rect 5629 23607 5687 23613
rect 3605 23579 3663 23585
rect 3605 23545 3617 23579
rect 3651 23576 3663 23579
rect 3970 23576 3976 23588
rect 3651 23548 3976 23576
rect 3651 23545 3663 23548
rect 3605 23539 3663 23545
rect 3970 23536 3976 23548
rect 4028 23536 4034 23588
rect 4341 23579 4399 23585
rect 4341 23545 4353 23579
rect 4387 23576 4399 23579
rect 4798 23576 4804 23588
rect 4387 23548 4804 23576
rect 4387 23545 4399 23548
rect 4341 23539 4399 23545
rect 4798 23536 4804 23548
rect 4856 23536 4862 23588
rect 5537 23579 5595 23585
rect 5537 23545 5549 23579
rect 5583 23576 5595 23579
rect 6270 23576 6276 23588
rect 5583 23548 6276 23576
rect 5583 23545 5595 23548
rect 5537 23539 5595 23545
rect 6270 23536 6276 23548
rect 6328 23536 6334 23588
rect 2041 23511 2099 23517
rect 2041 23477 2053 23511
rect 2087 23508 2099 23511
rect 2222 23508 2228 23520
rect 2087 23480 2228 23508
rect 2087 23477 2099 23480
rect 2041 23471 2099 23477
rect 2222 23468 2228 23480
rect 2280 23468 2286 23520
rect 2406 23508 2412 23520
rect 2367 23480 2412 23508
rect 2406 23468 2412 23480
rect 2464 23468 2470 23520
rect 3234 23508 3240 23520
rect 3195 23480 3240 23508
rect 3234 23468 3240 23480
rect 3292 23468 3298 23520
rect 3786 23468 3792 23520
rect 3844 23508 3850 23520
rect 3881 23511 3939 23517
rect 3881 23508 3893 23511
rect 3844 23480 3893 23508
rect 3844 23468 3850 23480
rect 3881 23477 3893 23480
rect 3927 23477 3939 23511
rect 3881 23471 3939 23477
rect 4709 23511 4767 23517
rect 4709 23477 4721 23511
rect 4755 23508 4767 23511
rect 4890 23508 4896 23520
rect 4755 23480 4896 23508
rect 4755 23477 4767 23480
rect 4709 23471 4767 23477
rect 4890 23468 4896 23480
rect 4948 23468 4954 23520
rect 6181 23511 6239 23517
rect 6181 23477 6193 23511
rect 6227 23508 6239 23511
rect 6380 23508 6408 23616
rect 9030 23604 9036 23616
rect 9088 23604 9094 23656
rect 9122 23604 9128 23656
rect 9180 23644 9186 23656
rect 9289 23647 9347 23653
rect 9289 23644 9301 23647
rect 9180 23616 9301 23644
rect 9180 23604 9186 23616
rect 9289 23613 9301 23616
rect 9335 23613 9347 23647
rect 9289 23607 9347 23613
rect 10134 23604 10140 23656
rect 10192 23604 10198 23656
rect 10594 23604 10600 23656
rect 10652 23644 10658 23656
rect 11057 23647 11115 23653
rect 11057 23644 11069 23647
rect 10652 23616 11069 23644
rect 10652 23604 10658 23616
rect 11057 23613 11069 23616
rect 11103 23644 11115 23647
rect 11103 23616 12480 23644
rect 11103 23613 11115 23616
rect 11057 23607 11115 23613
rect 6641 23579 6699 23585
rect 6641 23545 6653 23579
rect 6687 23576 6699 23579
rect 6914 23576 6920 23588
rect 6687 23548 6920 23576
rect 6687 23545 6699 23548
rect 6641 23539 6699 23545
rect 6914 23536 6920 23548
rect 6972 23576 6978 23588
rect 7374 23576 7380 23588
rect 6972 23548 7380 23576
rect 6972 23536 6978 23548
rect 7374 23536 7380 23548
rect 7432 23536 7438 23588
rect 7742 23536 7748 23588
rect 7800 23576 7806 23588
rect 8113 23579 8171 23585
rect 8113 23576 8125 23579
rect 7800 23548 8125 23576
rect 7800 23536 7806 23548
rect 8113 23545 8125 23548
rect 8159 23545 8171 23579
rect 8113 23539 8171 23545
rect 6730 23508 6736 23520
rect 6227 23480 6736 23508
rect 6227 23477 6239 23480
rect 6181 23471 6239 23477
rect 6730 23468 6736 23480
rect 6788 23468 6794 23520
rect 7558 23468 7564 23520
rect 7616 23508 7622 23520
rect 8021 23511 8079 23517
rect 8021 23508 8033 23511
rect 7616 23480 8033 23508
rect 7616 23468 7622 23480
rect 8021 23477 8033 23480
rect 8067 23477 8079 23511
rect 8021 23471 8079 23477
rect 8294 23468 8300 23520
rect 8352 23508 8358 23520
rect 8481 23511 8539 23517
rect 8481 23508 8493 23511
rect 8352 23480 8493 23508
rect 8352 23468 8358 23480
rect 8481 23477 8493 23480
rect 8527 23477 8539 23511
rect 8846 23508 8852 23520
rect 8807 23480 8852 23508
rect 8481 23471 8539 23477
rect 8846 23468 8852 23480
rect 8904 23468 8910 23520
rect 9674 23468 9680 23520
rect 9732 23508 9738 23520
rect 10152 23508 10180 23604
rect 11885 23579 11943 23585
rect 11885 23545 11897 23579
rect 11931 23576 11943 23579
rect 12342 23576 12348 23588
rect 11931 23548 12348 23576
rect 11931 23545 11943 23548
rect 11885 23539 11943 23545
rect 12342 23536 12348 23548
rect 12400 23536 12406 23588
rect 10413 23511 10471 23517
rect 10413 23508 10425 23511
rect 9732 23480 10425 23508
rect 9732 23468 9738 23480
rect 10413 23477 10425 23480
rect 10459 23477 10471 23511
rect 10413 23471 10471 23477
rect 11146 23468 11152 23520
rect 11204 23508 11210 23520
rect 12069 23511 12127 23517
rect 12069 23508 12081 23511
rect 11204 23480 12081 23508
rect 11204 23468 11210 23480
rect 12069 23477 12081 23480
rect 12115 23508 12127 23511
rect 12161 23511 12219 23517
rect 12161 23508 12173 23511
rect 12115 23480 12173 23508
rect 12115 23477 12127 23480
rect 12069 23471 12127 23477
rect 12161 23477 12173 23480
rect 12207 23477 12219 23511
rect 12452 23508 12480 23616
rect 12618 23604 12624 23656
rect 12676 23644 12682 23656
rect 12805 23647 12863 23653
rect 12805 23644 12817 23647
rect 12676 23616 12817 23644
rect 12676 23604 12682 23616
rect 12805 23613 12817 23616
rect 12851 23613 12863 23647
rect 13446 23644 13452 23656
rect 13407 23616 13452 23644
rect 12805 23607 12863 23613
rect 13446 23604 13452 23616
rect 13504 23604 13510 23656
rect 14185 23647 14243 23653
rect 14185 23644 14197 23647
rect 14016 23616 14197 23644
rect 12710 23536 12716 23588
rect 12768 23576 12774 23588
rect 12989 23579 13047 23585
rect 12989 23576 13001 23579
rect 12768 23548 13001 23576
rect 12768 23536 12774 23548
rect 12989 23545 13001 23548
rect 13035 23545 13047 23579
rect 12989 23539 13047 23545
rect 13262 23536 13268 23588
rect 13320 23576 13326 23588
rect 13538 23576 13544 23588
rect 13320 23548 13544 23576
rect 13320 23536 13326 23548
rect 13538 23536 13544 23548
rect 13596 23536 13602 23588
rect 13446 23508 13452 23520
rect 12452 23480 13452 23508
rect 12161 23471 12219 23477
rect 13446 23468 13452 23480
rect 13504 23508 13510 23520
rect 14016 23517 14044 23616
rect 14185 23613 14197 23616
rect 14231 23613 14243 23647
rect 14185 23607 14243 23613
rect 16482 23604 16488 23656
rect 16540 23644 16546 23656
rect 16669 23647 16727 23653
rect 16669 23644 16681 23647
rect 16540 23616 16681 23644
rect 16540 23604 16546 23616
rect 16669 23613 16681 23616
rect 16715 23644 16727 23647
rect 17586 23644 17592 23656
rect 16715 23616 17592 23644
rect 16715 23613 16727 23616
rect 16669 23607 16727 23613
rect 17586 23604 17592 23616
rect 17644 23604 17650 23656
rect 18322 23604 18328 23656
rect 18380 23644 18386 23656
rect 18708 23644 18736 23675
rect 18782 23672 18788 23684
rect 18840 23672 18846 23724
rect 18892 23712 18920 23752
rect 19058 23740 19064 23792
rect 19116 23780 19122 23792
rect 19260 23780 19288 23820
rect 19613 23817 19625 23820
rect 19659 23848 19671 23851
rect 19702 23848 19708 23860
rect 19659 23820 19708 23848
rect 19659 23817 19671 23820
rect 19613 23811 19671 23817
rect 19702 23808 19708 23820
rect 19760 23808 19766 23860
rect 21177 23851 21235 23857
rect 21177 23817 21189 23851
rect 21223 23848 21235 23851
rect 22094 23848 22100 23860
rect 21223 23820 22100 23848
rect 21223 23817 21235 23820
rect 21177 23811 21235 23817
rect 22094 23808 22100 23820
rect 22152 23848 22158 23860
rect 22557 23851 22615 23857
rect 22557 23848 22569 23851
rect 22152 23820 22569 23848
rect 22152 23808 22158 23820
rect 22557 23817 22569 23820
rect 22603 23817 22615 23851
rect 22830 23848 22836 23860
rect 22791 23820 22836 23848
rect 22557 23811 22615 23817
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 25682 23848 25688 23860
rect 25643 23820 25688 23848
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 19116 23752 19288 23780
rect 19797 23783 19855 23789
rect 19116 23740 19122 23752
rect 19797 23749 19809 23783
rect 19843 23780 19855 23783
rect 20806 23780 20812 23792
rect 19843 23752 20812 23780
rect 19843 23749 19855 23752
rect 19797 23743 19855 23749
rect 20806 23740 20812 23752
rect 20864 23740 20870 23792
rect 21358 23780 21364 23792
rect 21319 23752 21364 23780
rect 21358 23740 21364 23752
rect 21416 23740 21422 23792
rect 23474 23780 23480 23792
rect 21468 23752 23480 23780
rect 21468 23712 21496 23752
rect 23474 23740 23480 23752
rect 23532 23740 23538 23792
rect 24026 23780 24032 23792
rect 23987 23752 24032 23780
rect 24026 23740 24032 23752
rect 24084 23740 24090 23792
rect 21818 23712 21824 23724
rect 18892 23684 21496 23712
rect 21744 23684 21824 23712
rect 18380 23616 18736 23644
rect 18380 23604 18386 23616
rect 18966 23604 18972 23656
rect 19024 23644 19030 23656
rect 20073 23647 20131 23653
rect 20073 23644 20085 23647
rect 19024 23616 20085 23644
rect 19024 23604 19030 23616
rect 20073 23613 20085 23616
rect 20119 23613 20131 23647
rect 21634 23644 21640 23656
rect 21595 23616 21640 23644
rect 20073 23607 20131 23613
rect 21634 23604 21640 23616
rect 21692 23604 21698 23656
rect 14452 23579 14510 23585
rect 14452 23545 14464 23579
rect 14498 23576 14510 23579
rect 14734 23576 14740 23588
rect 14498 23548 14740 23576
rect 14498 23545 14510 23548
rect 14452 23539 14510 23545
rect 14734 23536 14740 23548
rect 14792 23536 14798 23588
rect 15286 23536 15292 23588
rect 15344 23576 15350 23588
rect 15746 23576 15752 23588
rect 15344 23548 15752 23576
rect 15344 23536 15350 23548
rect 15746 23536 15752 23548
rect 15804 23536 15810 23588
rect 16945 23579 17003 23585
rect 16945 23576 16957 23579
rect 16684 23548 16957 23576
rect 16684 23520 16712 23548
rect 16945 23545 16957 23548
rect 16991 23545 17003 23579
rect 16945 23539 17003 23545
rect 18138 23536 18144 23588
rect 18196 23576 18202 23588
rect 18417 23579 18475 23585
rect 18417 23576 18429 23579
rect 18196 23548 18429 23576
rect 18196 23536 18202 23548
rect 18417 23545 18429 23548
rect 18463 23545 18475 23579
rect 18598 23576 18604 23588
rect 18559 23548 18604 23576
rect 18417 23539 18475 23545
rect 18598 23536 18604 23548
rect 18656 23536 18662 23588
rect 20346 23576 20352 23588
rect 20307 23548 20352 23576
rect 20346 23536 20352 23548
rect 20404 23536 20410 23588
rect 14001 23511 14059 23517
rect 14001 23508 14013 23511
rect 13504 23480 14013 23508
rect 13504 23468 13510 23480
rect 14001 23477 14013 23480
rect 14047 23477 14059 23511
rect 16206 23508 16212 23520
rect 16167 23480 16212 23508
rect 14001 23471 14059 23477
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 16666 23468 16672 23520
rect 16724 23468 16730 23520
rect 17865 23511 17923 23517
rect 17865 23477 17877 23511
rect 17911 23508 17923 23511
rect 18616 23508 18644 23536
rect 17911 23480 18644 23508
rect 17911 23477 17923 23480
rect 17865 23471 17923 23477
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 20257 23511 20315 23517
rect 20257 23508 20269 23511
rect 20036 23480 20269 23508
rect 20036 23468 20042 23480
rect 20257 23477 20269 23480
rect 20303 23477 20315 23511
rect 20257 23471 20315 23477
rect 20809 23511 20867 23517
rect 20809 23477 20821 23511
rect 20855 23508 20867 23511
rect 21082 23508 21088 23520
rect 20855 23480 21088 23508
rect 20855 23477 20867 23480
rect 20809 23471 20867 23477
rect 21082 23468 21088 23480
rect 21140 23468 21146 23520
rect 21744 23508 21772 23684
rect 21818 23672 21824 23684
rect 21876 23712 21882 23724
rect 21913 23715 21971 23721
rect 21913 23712 21925 23715
rect 21876 23684 21925 23712
rect 21876 23672 21882 23684
rect 21913 23681 21925 23684
rect 21959 23681 21971 23715
rect 21913 23675 21971 23681
rect 24210 23672 24216 23724
rect 24268 23712 24274 23724
rect 24581 23715 24639 23721
rect 24581 23712 24593 23715
rect 24268 23684 24593 23712
rect 24268 23672 24274 23684
rect 24581 23681 24593 23684
rect 24627 23681 24639 23715
rect 24581 23675 24639 23681
rect 22554 23644 22560 23656
rect 21836 23616 22560 23644
rect 21836 23585 21864 23616
rect 22554 23604 22560 23616
rect 22612 23604 22618 23656
rect 25498 23644 25504 23656
rect 25459 23616 25504 23644
rect 25498 23604 25504 23616
rect 25556 23644 25562 23656
rect 26053 23647 26111 23653
rect 26053 23644 26065 23647
rect 25556 23616 26065 23644
rect 25556 23604 25562 23616
rect 26053 23613 26065 23616
rect 26099 23613 26111 23647
rect 26053 23607 26111 23613
rect 21821 23579 21879 23585
rect 21821 23545 21833 23579
rect 21867 23545 21879 23579
rect 22094 23576 22100 23588
rect 21821 23539 21879 23545
rect 21928 23548 22100 23576
rect 21928 23508 21956 23548
rect 22094 23536 22100 23548
rect 22152 23536 22158 23588
rect 22830 23536 22836 23588
rect 22888 23576 22894 23588
rect 23109 23579 23167 23585
rect 23109 23576 23121 23579
rect 22888 23548 23121 23576
rect 22888 23536 22894 23548
rect 23109 23545 23121 23548
rect 23155 23576 23167 23579
rect 23382 23576 23388 23588
rect 23155 23548 23388 23576
rect 23155 23545 23167 23548
rect 23109 23539 23167 23545
rect 23382 23536 23388 23548
rect 23440 23536 23446 23588
rect 23474 23536 23480 23588
rect 23532 23576 23538 23588
rect 24118 23576 24124 23588
rect 23532 23548 24124 23576
rect 23532 23536 23538 23548
rect 24118 23536 24124 23548
rect 24176 23576 24182 23588
rect 24305 23579 24363 23585
rect 24305 23576 24317 23579
rect 24176 23548 24317 23576
rect 24176 23536 24182 23548
rect 24305 23545 24317 23548
rect 24351 23545 24363 23579
rect 24305 23539 24363 23545
rect 21744 23480 21956 23508
rect 22186 23468 22192 23520
rect 22244 23508 22250 23520
rect 22373 23511 22431 23517
rect 22373 23508 22385 23511
rect 22244 23480 22385 23508
rect 22244 23468 22250 23480
rect 22373 23477 22385 23480
rect 22419 23477 22431 23511
rect 22373 23471 22431 23477
rect 22557 23511 22615 23517
rect 22557 23477 22569 23511
rect 22603 23508 22615 23511
rect 23014 23508 23020 23520
rect 22603 23480 23020 23508
rect 22603 23477 22615 23480
rect 22557 23471 22615 23477
rect 23014 23468 23020 23480
rect 23072 23468 23078 23520
rect 23934 23468 23940 23520
rect 23992 23508 23998 23520
rect 24489 23511 24547 23517
rect 24489 23508 24501 23511
rect 23992 23480 24501 23508
rect 23992 23468 23998 23480
rect 24489 23477 24501 23480
rect 24535 23477 24547 23511
rect 24946 23508 24952 23520
rect 24907 23480 24952 23508
rect 24489 23471 24547 23477
rect 24946 23468 24952 23480
rect 25004 23468 25010 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1486 23264 1492 23316
rect 1544 23304 1550 23316
rect 1581 23307 1639 23313
rect 1581 23304 1593 23307
rect 1544 23276 1593 23304
rect 1544 23264 1550 23276
rect 1581 23273 1593 23276
rect 1627 23273 1639 23307
rect 1581 23267 1639 23273
rect 5537 23307 5595 23313
rect 5537 23273 5549 23307
rect 5583 23304 5595 23307
rect 5626 23304 5632 23316
rect 5583 23276 5632 23304
rect 5583 23273 5595 23276
rect 5537 23267 5595 23273
rect 5626 23264 5632 23276
rect 5684 23264 5690 23316
rect 11057 23307 11115 23313
rect 11057 23273 11069 23307
rect 11103 23273 11115 23307
rect 11057 23267 11115 23273
rect 6546 23196 6552 23248
rect 6604 23236 6610 23248
rect 7009 23239 7067 23245
rect 7009 23236 7021 23239
rect 6604 23208 7021 23236
rect 6604 23196 6610 23208
rect 7009 23205 7021 23208
rect 7055 23205 7067 23239
rect 8386 23236 8392 23248
rect 8347 23208 8392 23236
rect 7009 23199 7067 23205
rect 8386 23196 8392 23208
rect 8444 23196 8450 23248
rect 8570 23236 8576 23248
rect 8531 23208 8576 23236
rect 8570 23196 8576 23208
rect 8628 23196 8634 23248
rect 8665 23239 8723 23245
rect 8665 23205 8677 23239
rect 8711 23236 8723 23239
rect 8754 23236 8760 23248
rect 8711 23208 8760 23236
rect 8711 23205 8723 23208
rect 8665 23199 8723 23205
rect 8754 23196 8760 23208
rect 8812 23236 8818 23248
rect 9122 23236 9128 23248
rect 8812 23208 9128 23236
rect 8812 23196 8818 23208
rect 9122 23196 9128 23208
rect 9180 23236 9186 23248
rect 11072 23236 11100 23267
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 12805 23307 12863 23313
rect 12805 23304 12817 23307
rect 12492 23276 12817 23304
rect 12492 23264 12498 23276
rect 12805 23273 12817 23276
rect 12851 23273 12863 23307
rect 13262 23304 13268 23316
rect 13223 23276 13268 23304
rect 12805 23267 12863 23273
rect 13262 23264 13268 23276
rect 13320 23264 13326 23316
rect 15930 23264 15936 23316
rect 15988 23304 15994 23316
rect 16206 23304 16212 23316
rect 15988 23276 16212 23304
rect 15988 23264 15994 23276
rect 16206 23264 16212 23276
rect 16264 23264 16270 23316
rect 16393 23307 16451 23313
rect 16393 23273 16405 23307
rect 16439 23304 16451 23307
rect 16574 23304 16580 23316
rect 16439 23276 16580 23304
rect 16439 23273 16451 23276
rect 16393 23267 16451 23273
rect 16574 23264 16580 23276
rect 16632 23264 16638 23316
rect 18138 23304 18144 23316
rect 18099 23276 18144 23304
rect 18138 23264 18144 23276
rect 18196 23264 18202 23316
rect 19334 23264 19340 23316
rect 19392 23304 19398 23316
rect 20070 23304 20076 23316
rect 19392 23276 20076 23304
rect 19392 23264 19398 23276
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 20165 23307 20223 23313
rect 20165 23273 20177 23307
rect 20211 23304 20223 23307
rect 20346 23304 20352 23316
rect 20211 23276 20352 23304
rect 20211 23273 20223 23276
rect 20165 23267 20223 23273
rect 20346 23264 20352 23276
rect 20404 23264 20410 23316
rect 20714 23264 20720 23316
rect 20772 23304 20778 23316
rect 21450 23304 21456 23316
rect 20772 23276 21456 23304
rect 20772 23264 20778 23276
rect 21450 23264 21456 23276
rect 21508 23264 21514 23316
rect 21910 23304 21916 23316
rect 21871 23276 21916 23304
rect 21910 23264 21916 23276
rect 21968 23264 21974 23316
rect 22823 23307 22881 23313
rect 22823 23273 22835 23307
rect 22869 23304 22881 23307
rect 24854 23304 24860 23316
rect 22869 23276 24716 23304
rect 24815 23276 24860 23304
rect 22869 23273 22881 23276
rect 22823 23267 22881 23273
rect 11422 23236 11428 23248
rect 9180 23208 11428 23236
rect 9180 23196 9186 23208
rect 11422 23196 11428 23208
rect 11480 23196 11486 23248
rect 15470 23196 15476 23248
rect 15528 23236 15534 23248
rect 15657 23239 15715 23245
rect 15657 23236 15669 23239
rect 15528 23208 15669 23236
rect 15528 23196 15534 23208
rect 15657 23205 15669 23208
rect 15703 23205 15715 23239
rect 15838 23236 15844 23248
rect 15799 23208 15844 23236
rect 15657 23199 15715 23205
rect 15838 23196 15844 23208
rect 15896 23196 15902 23248
rect 17402 23236 17408 23248
rect 17363 23208 17408 23236
rect 17402 23196 17408 23208
rect 17460 23196 17466 23248
rect 17954 23196 17960 23248
rect 18012 23236 18018 23248
rect 18785 23239 18843 23245
rect 18785 23236 18797 23239
rect 18012 23208 18797 23236
rect 18012 23196 18018 23208
rect 18785 23205 18797 23208
rect 18831 23236 18843 23239
rect 18874 23236 18880 23248
rect 18831 23208 18880 23236
rect 18831 23205 18843 23208
rect 18785 23199 18843 23205
rect 18874 23196 18880 23208
rect 18932 23196 18938 23248
rect 18966 23196 18972 23248
rect 19024 23236 19030 23248
rect 23293 23239 23351 23245
rect 19024 23208 19069 23236
rect 19024 23196 19030 23208
rect 23293 23205 23305 23239
rect 23339 23236 23351 23239
rect 23566 23236 23572 23248
rect 23339 23208 23572 23236
rect 23339 23205 23351 23208
rect 23293 23199 23351 23205
rect 23566 23196 23572 23208
rect 23624 23196 23630 23248
rect 24688 23245 24716 23276
rect 24854 23264 24860 23276
rect 24912 23304 24918 23316
rect 25317 23307 25375 23313
rect 25317 23304 25329 23307
rect 24912 23276 25329 23304
rect 24912 23264 24918 23276
rect 25317 23273 25329 23276
rect 25363 23273 25375 23307
rect 25317 23267 25375 23273
rect 24673 23239 24731 23245
rect 24673 23205 24685 23239
rect 24719 23205 24731 23239
rect 24673 23199 24731 23205
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23137 1455 23171
rect 1397 23131 1455 23137
rect 2501 23171 2559 23177
rect 2501 23137 2513 23171
rect 2547 23168 2559 23171
rect 2774 23168 2780 23180
rect 2547 23140 2780 23168
rect 2547 23137 2559 23140
rect 2501 23131 2559 23137
rect 1412 23100 1440 23131
rect 2774 23128 2780 23140
rect 2832 23128 2838 23180
rect 4982 23128 4988 23180
rect 5040 23168 5046 23180
rect 5353 23171 5411 23177
rect 5353 23168 5365 23171
rect 5040 23140 5365 23168
rect 5040 23128 5046 23140
rect 5353 23137 5365 23140
rect 5399 23137 5411 23171
rect 5353 23131 5411 23137
rect 6914 23128 6920 23180
rect 6972 23168 6978 23180
rect 7101 23171 7159 23177
rect 7101 23168 7113 23171
rect 6972 23140 7113 23168
rect 6972 23128 6978 23140
rect 7101 23137 7113 23140
rect 7147 23137 7159 23171
rect 7101 23131 7159 23137
rect 9944 23171 10002 23177
rect 9944 23137 9956 23171
rect 9990 23168 10002 23171
rect 10226 23168 10232 23180
rect 9990 23140 10232 23168
rect 9990 23137 10002 23140
rect 9944 23131 10002 23137
rect 10226 23128 10232 23140
rect 10284 23168 10290 23180
rect 11146 23168 11152 23180
rect 10284 23140 11152 23168
rect 10284 23128 10290 23140
rect 11146 23128 11152 23140
rect 11204 23128 11210 23180
rect 12158 23128 12164 23180
rect 12216 23168 12222 23180
rect 12621 23171 12679 23177
rect 12621 23168 12633 23171
rect 12216 23140 12633 23168
rect 12216 23128 12222 23140
rect 12621 23137 12633 23140
rect 12667 23137 12679 23171
rect 13906 23168 13912 23180
rect 13867 23140 13912 23168
rect 12621 23131 12679 23137
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 17497 23171 17555 23177
rect 17497 23168 17509 23171
rect 16684 23140 17509 23168
rect 1762 23100 1768 23112
rect 1412 23072 1768 23100
rect 1762 23060 1768 23072
rect 1820 23060 1826 23112
rect 4525 23103 4583 23109
rect 4525 23069 4537 23103
rect 4571 23100 4583 23103
rect 5074 23100 5080 23112
rect 4571 23072 5080 23100
rect 4571 23069 4583 23072
rect 4525 23063 4583 23069
rect 5074 23060 5080 23072
rect 5132 23060 5138 23112
rect 7006 23100 7012 23112
rect 6967 23072 7012 23100
rect 7006 23060 7012 23072
rect 7064 23060 7070 23112
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 9088 23072 9137 23100
rect 9088 23060 9094 23072
rect 9125 23069 9137 23072
rect 9171 23100 9183 23103
rect 9677 23103 9735 23109
rect 9677 23100 9689 23103
rect 9171 23072 9689 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9677 23069 9689 23072
rect 9723 23069 9735 23103
rect 9677 23063 9735 23069
rect 12897 23103 12955 23109
rect 12897 23069 12909 23103
rect 12943 23100 12955 23103
rect 12943 23072 13768 23100
rect 12943 23069 12955 23072
rect 12897 23063 12955 23069
rect 2958 22992 2964 23044
rect 3016 23032 3022 23044
rect 3421 23035 3479 23041
rect 3421 23032 3433 23035
rect 3016 23004 3433 23032
rect 3016 22992 3022 23004
rect 3421 23001 3433 23004
rect 3467 23001 3479 23035
rect 3421 22995 3479 23001
rect 6365 23035 6423 23041
rect 6365 23001 6377 23035
rect 6411 23032 6423 23035
rect 6822 23032 6828 23044
rect 6411 23004 6828 23032
rect 6411 23001 6423 23004
rect 6365 22995 6423 23001
rect 6822 22992 6828 23004
rect 6880 22992 6886 23044
rect 7282 22992 7288 23044
rect 7340 23032 7346 23044
rect 7742 23032 7748 23044
rect 7340 23004 7748 23032
rect 7340 22992 7346 23004
rect 7742 22992 7748 23004
rect 7800 23032 7806 23044
rect 7837 23035 7895 23041
rect 7837 23032 7849 23035
rect 7800 23004 7849 23032
rect 7800 22992 7806 23004
rect 7837 23001 7849 23004
rect 7883 23001 7895 23035
rect 8110 23032 8116 23044
rect 8071 23004 8116 23032
rect 7837 22995 7895 23001
rect 1946 22964 1952 22976
rect 1907 22936 1952 22964
rect 1946 22924 1952 22936
rect 2004 22924 2010 22976
rect 2314 22964 2320 22976
rect 2275 22936 2320 22964
rect 2314 22924 2320 22936
rect 2372 22924 2378 22976
rect 2406 22924 2412 22976
rect 2464 22964 2470 22976
rect 2685 22967 2743 22973
rect 2685 22964 2697 22967
rect 2464 22936 2697 22964
rect 2464 22924 2470 22936
rect 2685 22933 2697 22936
rect 2731 22933 2743 22967
rect 3050 22964 3056 22976
rect 3011 22936 3056 22964
rect 2685 22927 2743 22933
rect 3050 22924 3056 22936
rect 3108 22924 3114 22976
rect 3142 22924 3148 22976
rect 3200 22964 3206 22976
rect 3789 22967 3847 22973
rect 3789 22964 3801 22967
rect 3200 22936 3801 22964
rect 3200 22924 3206 22936
rect 3789 22933 3801 22936
rect 3835 22933 3847 22967
rect 3789 22927 3847 22933
rect 4522 22924 4528 22976
rect 4580 22964 4586 22976
rect 4801 22967 4859 22973
rect 4801 22964 4813 22967
rect 4580 22936 4813 22964
rect 4580 22924 4586 22936
rect 4801 22933 4813 22936
rect 4847 22933 4859 22967
rect 4801 22927 4859 22933
rect 5261 22967 5319 22973
rect 5261 22933 5273 22967
rect 5307 22964 5319 22967
rect 5442 22964 5448 22976
rect 5307 22936 5448 22964
rect 5307 22933 5319 22936
rect 5261 22927 5319 22933
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 5997 22967 6055 22973
rect 5997 22933 6009 22967
rect 6043 22964 6055 22967
rect 6086 22964 6092 22976
rect 6043 22936 6092 22964
rect 6043 22933 6055 22936
rect 5997 22927 6055 22933
rect 6086 22924 6092 22936
rect 6144 22924 6150 22976
rect 6454 22924 6460 22976
rect 6512 22964 6518 22976
rect 6549 22967 6607 22973
rect 6549 22964 6561 22967
rect 6512 22936 6561 22964
rect 6512 22924 6518 22936
rect 6549 22933 6561 22936
rect 6595 22933 6607 22967
rect 7558 22964 7564 22976
rect 7519 22936 7564 22964
rect 6549 22927 6607 22933
rect 7558 22924 7564 22936
rect 7616 22924 7622 22976
rect 7852 22964 7880 22995
rect 8110 22992 8116 23004
rect 8168 22992 8174 23044
rect 9030 22964 9036 22976
rect 7852 22936 9036 22964
rect 9030 22924 9036 22936
rect 9088 22924 9094 22976
rect 9122 22924 9128 22976
rect 9180 22964 9186 22976
rect 9306 22964 9312 22976
rect 9180 22936 9312 22964
rect 9180 22924 9186 22936
rect 9306 22924 9312 22936
rect 9364 22924 9370 22976
rect 9493 22967 9551 22973
rect 9493 22933 9505 22967
rect 9539 22964 9551 22967
rect 9582 22964 9588 22976
rect 9539 22936 9588 22964
rect 9539 22933 9551 22936
rect 9493 22927 9551 22933
rect 9582 22924 9588 22936
rect 9640 22924 9646 22976
rect 9692 22964 9720 23063
rect 12250 22992 12256 23044
rect 12308 23032 12314 23044
rect 12345 23035 12403 23041
rect 12345 23032 12357 23035
rect 12308 23004 12357 23032
rect 12308 22992 12314 23004
rect 12345 23001 12357 23004
rect 12391 23001 12403 23035
rect 12345 22995 12403 23001
rect 13740 22976 13768 23072
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 14093 23103 14151 23109
rect 14093 23100 14105 23103
rect 13872 23072 14105 23100
rect 13872 23060 13878 23072
rect 14093 23069 14105 23072
rect 14139 23069 14151 23103
rect 14093 23063 14151 23069
rect 15933 23103 15991 23109
rect 15933 23069 15945 23103
rect 15979 23069 15991 23103
rect 15933 23063 15991 23069
rect 15102 23032 15108 23044
rect 15063 23004 15108 23032
rect 15102 22992 15108 23004
rect 15160 22992 15166 23044
rect 15378 23032 15384 23044
rect 15339 23004 15384 23032
rect 15378 22992 15384 23004
rect 15436 22992 15442 23044
rect 15948 22976 15976 23063
rect 10318 22964 10324 22976
rect 9692 22936 10324 22964
rect 10318 22924 10324 22936
rect 10376 22924 10382 22976
rect 11330 22924 11336 22976
rect 11388 22964 11394 22976
rect 11609 22967 11667 22973
rect 11609 22964 11621 22967
rect 11388 22936 11621 22964
rect 11388 22924 11394 22936
rect 11609 22933 11621 22936
rect 11655 22933 11667 22967
rect 11974 22964 11980 22976
rect 11935 22936 11980 22964
rect 11609 22927 11667 22933
rect 11974 22924 11980 22936
rect 12032 22924 12038 22976
rect 13722 22964 13728 22976
rect 13683 22936 13728 22964
rect 13722 22924 13728 22936
rect 13780 22924 13786 22976
rect 14642 22964 14648 22976
rect 14603 22936 14648 22964
rect 14642 22924 14648 22936
rect 14700 22924 14706 22976
rect 15930 22924 15936 22976
rect 15988 22964 15994 22976
rect 16684 22973 16712 23140
rect 17497 23137 17509 23140
rect 17543 23137 17555 23171
rect 17497 23131 17555 23137
rect 18506 23128 18512 23180
rect 18564 23168 18570 23180
rect 21818 23168 21824 23180
rect 18564 23140 21824 23168
rect 18564 23128 18570 23140
rect 21818 23128 21824 23140
rect 21876 23128 21882 23180
rect 22094 23128 22100 23180
rect 22152 23168 22158 23180
rect 23385 23171 23443 23177
rect 23385 23168 23397 23171
rect 22152 23140 23397 23168
rect 22152 23128 22158 23140
rect 23385 23137 23397 23140
rect 23431 23137 23443 23171
rect 24688 23168 24716 23199
rect 24854 23168 24860 23180
rect 24688 23140 24860 23168
rect 23385 23131 23443 23137
rect 24854 23128 24860 23140
rect 24912 23128 24918 23180
rect 17405 23103 17463 23109
rect 17405 23069 17417 23103
rect 17451 23100 17463 23103
rect 17678 23100 17684 23112
rect 17451 23072 17684 23100
rect 17451 23069 17463 23072
rect 17405 23063 17463 23069
rect 17678 23060 17684 23072
rect 17736 23060 17742 23112
rect 19061 23103 19119 23109
rect 19061 23100 19073 23103
rect 18064 23072 19073 23100
rect 16942 23032 16948 23044
rect 16903 23004 16948 23032
rect 16942 22992 16948 23004
rect 17000 22992 17006 23044
rect 18064 22976 18092 23072
rect 19061 23069 19073 23072
rect 19107 23069 19119 23103
rect 21358 23100 21364 23112
rect 21319 23072 21364 23100
rect 19061 23063 19119 23069
rect 21358 23060 21364 23072
rect 21416 23060 21422 23112
rect 21542 23100 21548 23112
rect 21503 23072 21548 23100
rect 21542 23060 21548 23072
rect 21600 23100 21606 23112
rect 22646 23100 22652 23112
rect 21600 23072 22652 23100
rect 21600 23060 21606 23072
rect 22646 23060 22652 23072
rect 22704 23060 22710 23112
rect 23293 23103 23351 23109
rect 23293 23069 23305 23103
rect 23339 23069 23351 23103
rect 24946 23100 24952 23112
rect 24907 23072 24952 23100
rect 23293 23063 23351 23069
rect 19794 23032 19800 23044
rect 19352 23004 19800 23032
rect 19352 22976 19380 23004
rect 19794 22992 19800 23004
rect 19852 22992 19858 23044
rect 20346 22992 20352 23044
rect 20404 23032 20410 23044
rect 20993 23035 21051 23041
rect 20404 23004 20668 23032
rect 20404 22992 20410 23004
rect 16669 22967 16727 22973
rect 16669 22964 16681 22967
rect 15988 22936 16681 22964
rect 15988 22924 15994 22936
rect 16669 22933 16681 22936
rect 16715 22933 16727 22967
rect 16669 22927 16727 22933
rect 18046 22924 18052 22976
rect 18104 22924 18110 22976
rect 18138 22924 18144 22976
rect 18196 22964 18202 22976
rect 18509 22967 18567 22973
rect 18509 22964 18521 22967
rect 18196 22936 18521 22964
rect 18196 22924 18202 22936
rect 18509 22933 18521 22936
rect 18555 22933 18567 22967
rect 18509 22927 18567 22933
rect 19334 22924 19340 22976
rect 19392 22924 19398 22976
rect 19426 22924 19432 22976
rect 19484 22964 19490 22976
rect 19705 22967 19763 22973
rect 19705 22964 19717 22967
rect 19484 22936 19717 22964
rect 19484 22924 19490 22936
rect 19705 22933 19717 22936
rect 19751 22964 19763 22967
rect 19978 22964 19984 22976
rect 19751 22936 19984 22964
rect 19751 22933 19763 22936
rect 19705 22927 19763 22933
rect 19978 22924 19984 22936
rect 20036 22924 20042 22976
rect 20530 22964 20536 22976
rect 20491 22936 20536 22964
rect 20530 22924 20536 22936
rect 20588 22924 20594 22976
rect 20640 22964 20668 23004
rect 20993 23001 21005 23035
rect 21039 23032 21051 23035
rect 21634 23032 21640 23044
rect 21039 23004 21640 23032
rect 21039 23001 21051 23004
rect 20993 22995 21051 23001
rect 21634 22992 21640 23004
rect 21692 22992 21698 23044
rect 23308 23032 23336 23063
rect 24946 23060 24952 23072
rect 25004 23060 25010 23112
rect 23750 23032 23756 23044
rect 23308 23004 23756 23032
rect 23750 22992 23756 23004
rect 23808 22992 23814 23044
rect 24118 22992 24124 23044
rect 24176 23032 24182 23044
rect 25685 23035 25743 23041
rect 25685 23032 25697 23035
rect 24176 23004 25697 23032
rect 24176 22992 24182 23004
rect 25685 23001 25697 23004
rect 25731 23001 25743 23035
rect 25685 22995 25743 23001
rect 21174 22964 21180 22976
rect 20640 22936 21180 22964
rect 21174 22924 21180 22936
rect 21232 22964 21238 22976
rect 22186 22964 22192 22976
rect 21232 22936 22192 22964
rect 21232 22924 21238 22936
rect 22186 22924 22192 22936
rect 22244 22924 22250 22976
rect 22557 22967 22615 22973
rect 22557 22933 22569 22967
rect 22603 22964 22615 22967
rect 22738 22964 22744 22976
rect 22603 22936 22744 22964
rect 22603 22933 22615 22936
rect 22557 22927 22615 22933
rect 22738 22924 22744 22936
rect 22796 22924 22802 22976
rect 23934 22964 23940 22976
rect 23895 22936 23940 22964
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 24397 22967 24455 22973
rect 24397 22933 24409 22967
rect 24443 22964 24455 22967
rect 24670 22964 24676 22976
rect 24443 22936 24676 22964
rect 24443 22933 24455 22936
rect 24397 22927 24455 22933
rect 24670 22924 24676 22936
rect 24728 22924 24734 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2682 22760 2688 22772
rect 2643 22732 2688 22760
rect 2682 22720 2688 22732
rect 2740 22720 2746 22772
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 7377 22763 7435 22769
rect 7377 22760 7389 22763
rect 6972 22732 7389 22760
rect 6972 22720 6978 22732
rect 7377 22729 7389 22732
rect 7423 22729 7435 22763
rect 7377 22723 7435 22729
rect 7745 22763 7803 22769
rect 7745 22729 7757 22763
rect 7791 22760 7803 22763
rect 8386 22760 8392 22772
rect 7791 22732 8392 22760
rect 7791 22729 7803 22732
rect 7745 22723 7803 22729
rect 8386 22720 8392 22732
rect 8444 22720 8450 22772
rect 8570 22720 8576 22772
rect 8628 22760 8634 22772
rect 9309 22763 9367 22769
rect 9309 22760 9321 22763
rect 8628 22732 9321 22760
rect 8628 22720 8634 22732
rect 9309 22729 9321 22732
rect 9355 22729 9367 22763
rect 9309 22723 9367 22729
rect 10042 22720 10048 22772
rect 10100 22760 10106 22772
rect 10873 22763 10931 22769
rect 10873 22760 10885 22763
rect 10100 22732 10885 22760
rect 10100 22720 10106 22732
rect 10873 22729 10885 22732
rect 10919 22729 10931 22763
rect 10873 22723 10931 22729
rect 11609 22763 11667 22769
rect 11609 22729 11621 22763
rect 11655 22760 11667 22763
rect 11790 22760 11796 22772
rect 11655 22732 11796 22760
rect 11655 22729 11667 22732
rect 11609 22723 11667 22729
rect 11790 22720 11796 22732
rect 11848 22720 11854 22772
rect 14734 22760 14740 22772
rect 14695 22732 14740 22760
rect 14734 22720 14740 22732
rect 14792 22720 14798 22772
rect 15470 22720 15476 22772
rect 15528 22760 15534 22772
rect 15657 22763 15715 22769
rect 15657 22760 15669 22763
rect 15528 22732 15669 22760
rect 15528 22720 15534 22732
rect 15657 22729 15669 22732
rect 15703 22729 15715 22763
rect 16482 22760 16488 22772
rect 16443 22732 16488 22760
rect 15657 22723 15715 22729
rect 16482 22720 16488 22732
rect 16540 22720 16546 22772
rect 17402 22760 17408 22772
rect 17363 22732 17408 22760
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 20073 22763 20131 22769
rect 20073 22729 20085 22763
rect 20119 22760 20131 22763
rect 21542 22760 21548 22772
rect 20119 22732 21548 22760
rect 20119 22729 20131 22732
rect 20073 22723 20131 22729
rect 21542 22720 21548 22732
rect 21600 22720 21606 22772
rect 23382 22760 23388 22772
rect 23343 22732 23388 22760
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 25130 22720 25136 22772
rect 25188 22760 25194 22772
rect 25188 22732 25452 22760
rect 25188 22720 25194 22732
rect 1578 22692 1584 22704
rect 1539 22664 1584 22692
rect 1578 22652 1584 22664
rect 1636 22652 1642 22704
rect 4062 22652 4068 22704
rect 4120 22692 4126 22704
rect 5261 22695 5319 22701
rect 5261 22692 5273 22695
rect 4120 22664 5273 22692
rect 4120 22652 4126 22664
rect 5261 22661 5273 22664
rect 5307 22661 5319 22695
rect 8754 22692 8760 22704
rect 5261 22655 5319 22661
rect 5368 22664 7052 22692
rect 8715 22664 8760 22692
rect 2409 22627 2467 22633
rect 2409 22593 2421 22627
rect 2455 22624 2467 22627
rect 4709 22627 4767 22633
rect 2455 22596 4660 22624
rect 2455 22593 2467 22596
rect 2409 22587 2467 22593
rect 1394 22556 1400 22568
rect 1355 22528 1400 22556
rect 1394 22516 1400 22528
rect 1452 22516 1458 22568
rect 2516 22565 2544 22596
rect 2501 22559 2559 22565
rect 2501 22525 2513 22559
rect 2547 22556 2559 22559
rect 3605 22559 3663 22565
rect 3605 22556 3617 22559
rect 2547 22528 2581 22556
rect 3436 22528 3617 22556
rect 2547 22525 2559 22528
rect 2501 22519 2559 22525
rect 2866 22448 2872 22500
rect 2924 22488 2930 22500
rect 3436 22497 3464 22528
rect 3605 22525 3617 22528
rect 3651 22525 3663 22559
rect 4632 22556 4660 22596
rect 4709 22593 4721 22627
rect 4755 22624 4767 22627
rect 4982 22624 4988 22636
rect 4755 22596 4988 22624
rect 4755 22593 4767 22596
rect 4709 22587 4767 22593
rect 4982 22584 4988 22596
rect 5040 22624 5046 22636
rect 5368 22624 5396 22664
rect 5040 22596 5396 22624
rect 5040 22584 5046 22596
rect 5442 22584 5448 22636
rect 5500 22624 5506 22636
rect 5721 22627 5779 22633
rect 5721 22624 5733 22627
rect 5500 22596 5733 22624
rect 5500 22584 5506 22596
rect 5721 22593 5733 22596
rect 5767 22624 5779 22627
rect 6454 22624 6460 22636
rect 5767 22596 6460 22624
rect 5767 22593 5779 22596
rect 5721 22587 5779 22593
rect 6454 22584 6460 22596
rect 6512 22584 6518 22636
rect 5626 22556 5632 22568
rect 4632 22528 5632 22556
rect 3605 22519 3663 22525
rect 5626 22516 5632 22528
rect 5684 22516 5690 22568
rect 5813 22559 5871 22565
rect 5813 22525 5825 22559
rect 5859 22556 5871 22559
rect 6914 22556 6920 22568
rect 5859 22528 6920 22556
rect 5859 22525 5871 22528
rect 5813 22519 5871 22525
rect 3421 22491 3479 22497
rect 3421 22488 3433 22491
rect 2924 22460 3433 22488
rect 2924 22448 2930 22460
rect 3421 22457 3433 22460
rect 3467 22457 3479 22491
rect 3421 22451 3479 22457
rect 4154 22448 4160 22500
rect 4212 22488 4218 22500
rect 4341 22491 4399 22497
rect 4341 22488 4353 22491
rect 4212 22460 4353 22488
rect 4212 22448 4218 22460
rect 4341 22457 4353 22460
rect 4387 22488 4399 22491
rect 5828 22488 5856 22519
rect 6914 22516 6920 22528
rect 6972 22516 6978 22568
rect 7024 22556 7052 22664
rect 8754 22652 8760 22664
rect 8812 22652 8818 22704
rect 16301 22695 16359 22701
rect 16301 22661 16313 22695
rect 16347 22692 16359 22695
rect 16758 22692 16764 22704
rect 16347 22664 16764 22692
rect 16347 22661 16359 22664
rect 16301 22655 16359 22661
rect 16758 22652 16764 22664
rect 16816 22692 16822 22704
rect 17678 22692 17684 22704
rect 16816 22664 17684 22692
rect 16816 22652 16822 22664
rect 17678 22652 17684 22664
rect 17736 22652 17742 22704
rect 19334 22652 19340 22704
rect 19392 22692 19398 22704
rect 19702 22692 19708 22704
rect 19392 22664 19708 22692
rect 19392 22652 19398 22664
rect 19702 22652 19708 22664
rect 19760 22652 19766 22704
rect 19794 22652 19800 22704
rect 19852 22692 19858 22704
rect 20625 22695 20683 22701
rect 20625 22692 20637 22695
rect 19852 22664 20637 22692
rect 19852 22652 19858 22664
rect 20625 22661 20637 22664
rect 20671 22661 20683 22695
rect 23750 22692 23756 22704
rect 23663 22664 23756 22692
rect 20625 22655 20683 22661
rect 23750 22652 23756 22664
rect 23808 22692 23814 22704
rect 24762 22692 24768 22704
rect 23808 22664 24768 22692
rect 23808 22652 23814 22664
rect 24762 22652 24768 22664
rect 24820 22652 24826 22704
rect 7098 22584 7104 22636
rect 7156 22624 7162 22636
rect 8018 22624 8024 22636
rect 7156 22596 8024 22624
rect 7156 22584 7162 22596
rect 8018 22584 8024 22596
rect 8076 22624 8082 22636
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 8076 22596 8125 22624
rect 8076 22584 8082 22596
rect 8113 22593 8125 22596
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 9769 22627 9827 22633
rect 9769 22593 9781 22627
rect 9815 22624 9827 22627
rect 10778 22624 10784 22636
rect 9815 22596 10784 22624
rect 9815 22593 9827 22596
rect 9769 22587 9827 22593
rect 10778 22584 10784 22596
rect 10836 22584 10842 22636
rect 11238 22624 11244 22636
rect 11199 22596 11244 22624
rect 11238 22584 11244 22596
rect 11296 22584 11302 22636
rect 11422 22624 11428 22636
rect 11383 22596 11428 22624
rect 11422 22584 11428 22596
rect 11480 22584 11486 22636
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22624 17095 22627
rect 17221 22627 17279 22633
rect 17221 22624 17233 22627
rect 17083 22596 17233 22624
rect 17083 22593 17095 22596
rect 17037 22587 17095 22593
rect 17221 22593 17233 22596
rect 17267 22593 17279 22627
rect 17221 22587 17279 22593
rect 20441 22627 20499 22633
rect 20441 22593 20453 22627
rect 20487 22624 20499 22627
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 20487 22596 21097 22624
rect 20487 22593 20499 22596
rect 20441 22587 20499 22593
rect 21085 22593 21097 22596
rect 21131 22624 21143 22627
rect 21266 22624 21272 22636
rect 21131 22596 21272 22624
rect 21131 22593 21143 22596
rect 21085 22587 21143 22593
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 22370 22624 22376 22636
rect 22331 22596 22376 22624
rect 22370 22584 22376 22596
rect 22428 22584 22434 22636
rect 24118 22624 24124 22636
rect 22480 22596 24124 22624
rect 7742 22556 7748 22568
rect 7024 22528 7748 22556
rect 7742 22516 7748 22528
rect 7800 22516 7806 22568
rect 8202 22516 8208 22568
rect 8260 22556 8266 22568
rect 8297 22559 8355 22565
rect 8297 22556 8309 22559
rect 8260 22528 8309 22556
rect 8260 22516 8266 22528
rect 8297 22525 8309 22528
rect 8343 22556 8355 22559
rect 9033 22559 9091 22565
rect 9033 22556 9045 22559
rect 8343 22528 9045 22556
rect 8343 22525 8355 22528
rect 8297 22519 8355 22525
rect 9033 22525 9045 22528
rect 9079 22556 9091 22559
rect 9861 22559 9919 22565
rect 9861 22556 9873 22559
rect 9079 22528 9873 22556
rect 9079 22525 9091 22528
rect 9033 22519 9091 22525
rect 9861 22525 9873 22528
rect 9907 22556 9919 22559
rect 10226 22556 10232 22568
rect 9907 22528 10232 22556
rect 9907 22525 9919 22528
rect 9861 22519 9919 22525
rect 10226 22516 10232 22528
rect 10284 22556 10290 22568
rect 10597 22559 10655 22565
rect 10597 22556 10609 22559
rect 10284 22528 10609 22556
rect 10284 22516 10290 22528
rect 10597 22525 10609 22528
rect 10643 22525 10655 22559
rect 12158 22556 12164 22568
rect 12119 22528 12164 22556
rect 10597 22519 10655 22525
rect 12158 22516 12164 22528
rect 12216 22516 12222 22568
rect 13357 22559 13415 22565
rect 13357 22556 13369 22559
rect 12636 22528 13369 22556
rect 9766 22488 9772 22500
rect 4387 22460 5856 22488
rect 9727 22460 9772 22488
rect 4387 22457 4399 22460
rect 4341 22451 4399 22457
rect 9766 22448 9772 22460
rect 9824 22448 9830 22500
rect 10318 22488 10324 22500
rect 10231 22460 10324 22488
rect 10318 22448 10324 22460
rect 10376 22488 10382 22500
rect 12636 22488 12664 22528
rect 13357 22525 13369 22528
rect 13403 22556 13415 22559
rect 13446 22556 13452 22568
rect 13403 22528 13452 22556
rect 13403 22525 13415 22528
rect 13357 22519 13415 22525
rect 13446 22516 13452 22528
rect 13504 22516 13510 22568
rect 14826 22516 14832 22568
rect 14884 22556 14890 22568
rect 14884 22528 17172 22556
rect 14884 22516 14890 22528
rect 10376 22460 12664 22488
rect 10376 22448 10382 22460
rect 1762 22380 1768 22432
rect 1820 22420 1826 22432
rect 1949 22423 2007 22429
rect 1949 22420 1961 22423
rect 1820 22392 1961 22420
rect 1820 22380 1826 22392
rect 1949 22389 1961 22392
rect 1995 22389 2007 22423
rect 1949 22383 2007 22389
rect 2774 22380 2780 22432
rect 2832 22420 2838 22432
rect 3053 22423 3111 22429
rect 3053 22420 3065 22423
rect 2832 22392 3065 22420
rect 2832 22380 2838 22392
rect 3053 22389 3065 22392
rect 3099 22389 3111 22423
rect 3053 22383 3111 22389
rect 3510 22380 3516 22432
rect 3568 22420 3574 22432
rect 3789 22423 3847 22429
rect 3789 22420 3801 22423
rect 3568 22392 3801 22420
rect 3568 22380 3574 22392
rect 3789 22389 3801 22392
rect 3835 22389 3847 22423
rect 3789 22383 3847 22389
rect 5077 22423 5135 22429
rect 5077 22389 5089 22423
rect 5123 22420 5135 22423
rect 5718 22420 5724 22432
rect 5123 22392 5724 22420
rect 5123 22389 5135 22392
rect 5077 22383 5135 22389
rect 5718 22380 5724 22392
rect 5776 22380 5782 22432
rect 6546 22420 6552 22432
rect 6507 22392 6552 22420
rect 6546 22380 6552 22392
rect 6604 22380 6610 22432
rect 7098 22420 7104 22432
rect 7059 22392 7104 22420
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 7834 22380 7840 22432
rect 7892 22420 7898 22432
rect 8205 22423 8263 22429
rect 8205 22420 8217 22423
rect 7892 22392 8217 22420
rect 7892 22380 7898 22392
rect 8205 22389 8217 22392
rect 8251 22389 8263 22423
rect 8205 22383 8263 22389
rect 11333 22423 11391 22429
rect 11333 22389 11345 22423
rect 11379 22420 11391 22423
rect 11609 22423 11667 22429
rect 11609 22420 11621 22423
rect 11379 22392 11621 22420
rect 11379 22389 11391 22392
rect 11333 22383 11391 22389
rect 11609 22389 11621 22392
rect 11655 22389 11667 22423
rect 11882 22420 11888 22432
rect 11843 22392 11888 22420
rect 11609 22383 11667 22389
rect 11882 22380 11888 22392
rect 11940 22380 11946 22432
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 12636 22420 12664 22460
rect 12713 22491 12771 22497
rect 12713 22457 12725 22491
rect 12759 22488 12771 22491
rect 13624 22491 13682 22497
rect 13624 22488 13636 22491
rect 12759 22460 13636 22488
rect 12759 22457 12771 22460
rect 12713 22451 12771 22457
rect 13624 22457 13636 22460
rect 13670 22488 13682 22491
rect 13722 22488 13728 22500
rect 13670 22460 13728 22488
rect 13670 22457 13682 22460
rect 13624 22451 13682 22457
rect 13722 22448 13728 22460
rect 13780 22448 13786 22500
rect 16482 22448 16488 22500
rect 16540 22488 16546 22500
rect 16761 22491 16819 22497
rect 16761 22488 16773 22491
rect 16540 22460 16773 22488
rect 16540 22448 16546 22460
rect 16761 22457 16773 22460
rect 16807 22457 16819 22491
rect 16761 22451 16819 22457
rect 16850 22448 16856 22500
rect 16908 22488 16914 22500
rect 16945 22491 17003 22497
rect 16945 22488 16957 22491
rect 16908 22460 16957 22488
rect 16908 22448 16914 22460
rect 16945 22457 16957 22460
rect 16991 22457 17003 22491
rect 17144 22488 17172 22528
rect 17494 22516 17500 22568
rect 17552 22556 17558 22568
rect 17773 22559 17831 22565
rect 17773 22556 17785 22559
rect 17552 22528 17785 22556
rect 17552 22516 17558 22528
rect 17773 22525 17785 22528
rect 17819 22556 17831 22559
rect 18049 22559 18107 22565
rect 18049 22556 18061 22559
rect 17819 22528 18061 22556
rect 17819 22525 17831 22528
rect 17773 22519 17831 22525
rect 18049 22525 18061 22528
rect 18095 22525 18107 22559
rect 18049 22519 18107 22525
rect 19334 22516 19340 22568
rect 19392 22556 19398 22568
rect 20257 22559 20315 22565
rect 20257 22556 20269 22559
rect 19392 22528 20269 22556
rect 19392 22516 19398 22528
rect 20257 22525 20269 22528
rect 20303 22525 20315 22559
rect 20257 22519 20315 22525
rect 20530 22516 20536 22568
rect 20588 22556 20594 22568
rect 21177 22559 21235 22565
rect 21177 22556 21189 22559
rect 20588 22528 21189 22556
rect 20588 22516 20594 22528
rect 21177 22525 21189 22528
rect 21223 22525 21235 22559
rect 22094 22556 22100 22568
rect 22007 22528 22100 22556
rect 21177 22519 21235 22525
rect 22094 22516 22100 22528
rect 22152 22556 22158 22568
rect 22480 22556 22508 22596
rect 24118 22584 24124 22596
rect 24176 22584 24182 22636
rect 24946 22584 24952 22636
rect 25004 22584 25010 22636
rect 25424 22633 25452 22732
rect 25409 22627 25467 22633
rect 25409 22593 25421 22627
rect 25455 22593 25467 22627
rect 25409 22587 25467 22593
rect 22152 22528 22508 22556
rect 22152 22516 22158 22528
rect 23842 22516 23848 22568
rect 23900 22556 23906 22568
rect 24673 22559 24731 22565
rect 24673 22556 24685 22559
rect 23900 22528 24685 22556
rect 23900 22516 23906 22528
rect 24673 22525 24685 22528
rect 24719 22556 24731 22559
rect 24964 22556 24992 22584
rect 25222 22556 25228 22568
rect 24719 22528 24992 22556
rect 25183 22528 25228 22556
rect 24719 22525 24731 22528
rect 24673 22519 24731 22525
rect 25222 22516 25228 22528
rect 25280 22556 25286 22568
rect 25961 22559 26019 22565
rect 25961 22556 25973 22559
rect 25280 22528 25973 22556
rect 25280 22516 25286 22528
rect 25961 22525 25973 22528
rect 26007 22525 26019 22559
rect 25961 22519 26019 22525
rect 17144 22460 18092 22488
rect 16945 22451 17003 22457
rect 13173 22423 13231 22429
rect 13173 22420 13185 22423
rect 12492 22392 13185 22420
rect 12492 22380 12498 22392
rect 13173 22389 13185 22392
rect 13219 22389 13231 22423
rect 13173 22383 13231 22389
rect 13262 22380 13268 22432
rect 13320 22420 13326 22432
rect 15289 22423 15347 22429
rect 15289 22420 15301 22423
rect 13320 22392 15301 22420
rect 13320 22380 13326 22392
rect 15289 22389 15301 22392
rect 15335 22420 15347 22423
rect 15838 22420 15844 22432
rect 15335 22392 15844 22420
rect 15335 22389 15347 22392
rect 15289 22383 15347 22389
rect 15838 22380 15844 22392
rect 15896 22380 15902 22432
rect 17218 22420 17224 22432
rect 17131 22392 17224 22420
rect 17218 22380 17224 22392
rect 17276 22420 17282 22432
rect 17862 22420 17868 22432
rect 17276 22392 17868 22420
rect 17276 22380 17282 22392
rect 17862 22380 17868 22392
rect 17920 22380 17926 22432
rect 18064 22420 18092 22460
rect 18230 22448 18236 22500
rect 18288 22497 18294 22500
rect 18288 22491 18352 22497
rect 18288 22457 18306 22491
rect 18340 22457 18352 22491
rect 20438 22488 20444 22500
rect 18288 22451 18352 22457
rect 18432 22460 20444 22488
rect 18288 22448 18294 22451
rect 18432 22420 18460 22460
rect 20438 22448 20444 22460
rect 20496 22448 20502 22500
rect 21358 22488 21364 22500
rect 20640 22460 21364 22488
rect 18064 22392 18460 22420
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19429 22423 19487 22429
rect 19429 22420 19441 22423
rect 19392 22392 19441 22420
rect 19392 22380 19398 22392
rect 19429 22389 19441 22392
rect 19475 22389 19487 22423
rect 19429 22383 19487 22389
rect 20257 22423 20315 22429
rect 20257 22389 20269 22423
rect 20303 22420 20315 22423
rect 20640 22420 20668 22460
rect 21358 22448 21364 22460
rect 21416 22488 21422 22500
rect 21545 22491 21603 22497
rect 21545 22488 21557 22491
rect 21416 22460 21557 22488
rect 21416 22448 21422 22460
rect 21545 22457 21557 22460
rect 21591 22457 21603 22491
rect 21545 22451 21603 22457
rect 23658 22448 23664 22500
rect 23716 22488 23722 22500
rect 24029 22491 24087 22497
rect 24029 22488 24041 22491
rect 23716 22460 24041 22488
rect 23716 22448 23722 22460
rect 24029 22457 24041 22460
rect 24075 22457 24087 22491
rect 24029 22451 24087 22457
rect 24305 22491 24363 22497
rect 24305 22457 24317 22491
rect 24351 22488 24363 22491
rect 25314 22488 25320 22500
rect 24351 22460 25320 22488
rect 24351 22457 24363 22460
rect 24305 22451 24363 22457
rect 25314 22448 25320 22460
rect 25372 22448 25378 22500
rect 20303 22392 20668 22420
rect 20303 22389 20315 22392
rect 20257 22383 20315 22389
rect 20714 22380 20720 22432
rect 20772 22420 20778 22432
rect 21085 22423 21143 22429
rect 21085 22420 21097 22423
rect 20772 22392 21097 22420
rect 20772 22380 20778 22392
rect 21085 22389 21097 22392
rect 21131 22389 21143 22423
rect 21085 22383 21143 22389
rect 22005 22423 22063 22429
rect 22005 22389 22017 22423
rect 22051 22420 22063 22423
rect 22186 22420 22192 22432
rect 22051 22392 22192 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 22186 22380 22192 22392
rect 22244 22380 22250 22432
rect 23109 22423 23167 22429
rect 23109 22389 23121 22423
rect 23155 22420 23167 22423
rect 23382 22420 23388 22432
rect 23155 22392 23388 22420
rect 23155 22389 23167 22392
rect 23109 22383 23167 22389
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 23474 22380 23480 22432
rect 23532 22420 23538 22432
rect 24213 22423 24271 22429
rect 24213 22420 24225 22423
rect 23532 22392 24225 22420
rect 23532 22380 23538 22392
rect 24213 22389 24225 22392
rect 24259 22389 24271 22423
rect 24213 22383 24271 22389
rect 24854 22380 24860 22432
rect 24912 22420 24918 22432
rect 25041 22423 25099 22429
rect 25041 22420 25053 22423
rect 24912 22392 25053 22420
rect 24912 22380 24918 22392
rect 25041 22389 25053 22392
rect 25087 22389 25099 22423
rect 25041 22383 25099 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1394 22176 1400 22228
rect 1452 22216 1458 22228
rect 1949 22219 2007 22225
rect 1949 22216 1961 22219
rect 1452 22188 1961 22216
rect 1452 22176 1458 22188
rect 1949 22185 1961 22188
rect 1995 22216 2007 22219
rect 2038 22216 2044 22228
rect 1995 22188 2044 22216
rect 1995 22185 2007 22188
rect 1949 22179 2007 22185
rect 2038 22176 2044 22188
rect 2096 22176 2102 22228
rect 5442 22216 5448 22228
rect 5403 22188 5448 22216
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 6539 22219 6597 22225
rect 6539 22185 6551 22219
rect 6585 22216 6597 22219
rect 7834 22216 7840 22228
rect 6585 22188 7840 22216
rect 6585 22185 6597 22188
rect 6539 22179 6597 22185
rect 7834 22176 7840 22188
rect 7892 22176 7898 22228
rect 11054 22176 11060 22228
rect 11112 22216 11118 22228
rect 12986 22216 12992 22228
rect 11112 22188 12992 22216
rect 11112 22176 11118 22188
rect 12986 22176 12992 22188
rect 13044 22176 13050 22228
rect 16485 22219 16543 22225
rect 16485 22185 16497 22219
rect 16531 22216 16543 22219
rect 17218 22216 17224 22228
rect 16531 22188 17224 22216
rect 16531 22185 16543 22188
rect 16485 22179 16543 22185
rect 17218 22176 17224 22188
rect 17276 22176 17282 22228
rect 17957 22219 18015 22225
rect 17957 22185 17969 22219
rect 18003 22216 18015 22219
rect 18230 22216 18236 22228
rect 18003 22188 18236 22216
rect 18003 22185 18015 22188
rect 17957 22179 18015 22185
rect 18230 22176 18236 22188
rect 18288 22176 18294 22228
rect 18340 22188 19288 22216
rect 4154 22108 4160 22160
rect 4212 22108 4218 22160
rect 7009 22151 7067 22157
rect 7009 22117 7021 22151
rect 7055 22148 7067 22151
rect 7190 22148 7196 22160
rect 7055 22120 7196 22148
rect 7055 22117 7067 22120
rect 7009 22111 7067 22117
rect 7190 22108 7196 22120
rect 7248 22108 7254 22160
rect 8573 22151 8631 22157
rect 8573 22148 8585 22151
rect 8303 22120 8585 22148
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22049 1455 22083
rect 2498 22080 2504 22092
rect 2459 22052 2504 22080
rect 1397 22043 1455 22049
rect 1412 22012 1440 22043
rect 2498 22040 2504 22052
rect 2556 22040 2562 22092
rect 3326 22040 3332 22092
rect 3384 22080 3390 22092
rect 4172 22080 4200 22108
rect 3384 22052 4200 22080
rect 6365 22083 6423 22089
rect 3384 22040 3390 22052
rect 6365 22049 6377 22083
rect 6411 22080 6423 22083
rect 7101 22083 7159 22089
rect 7101 22080 7113 22083
rect 6411 22052 7113 22080
rect 6411 22049 6423 22052
rect 6365 22043 6423 22049
rect 7101 22049 7113 22052
rect 7147 22080 7159 22083
rect 7282 22080 7288 22092
rect 7147 22052 7288 22080
rect 7147 22049 7159 22052
rect 7101 22043 7159 22049
rect 7282 22040 7288 22052
rect 7340 22040 7346 22092
rect 7745 22083 7803 22089
rect 7745 22049 7757 22083
rect 7791 22080 7803 22083
rect 8202 22080 8208 22092
rect 7791 22052 8208 22080
rect 7791 22049 7803 22052
rect 7745 22043 7803 22049
rect 8202 22040 8208 22052
rect 8260 22040 8266 22092
rect 1854 22012 1860 22024
rect 1412 21984 1860 22012
rect 1854 21972 1860 21984
rect 1912 21972 1918 22024
rect 3878 21972 3884 22024
rect 3936 22012 3942 22024
rect 4706 22012 4712 22024
rect 3936 21984 4712 22012
rect 3936 21972 3942 21984
rect 4706 21972 4712 21984
rect 4764 22012 4770 22024
rect 5353 22015 5411 22021
rect 5353 22012 5365 22015
rect 4764 21984 5365 22012
rect 4764 21972 4770 21984
rect 5353 21981 5365 21984
rect 5399 21981 5411 22015
rect 5534 22012 5540 22024
rect 5495 21984 5540 22012
rect 5353 21975 5411 21981
rect 5534 21972 5540 21984
rect 5592 21972 5598 22024
rect 7006 22012 7012 22024
rect 6967 21984 7012 22012
rect 7006 21972 7012 21984
rect 7064 21972 7070 22024
rect 7834 21972 7840 22024
rect 7892 22012 7898 22024
rect 8303 22012 8331 22120
rect 8573 22117 8585 22120
rect 8619 22117 8631 22151
rect 8573 22111 8631 22117
rect 9122 22108 9128 22160
rect 9180 22148 9186 22160
rect 9398 22148 9404 22160
rect 9180 22120 9404 22148
rect 9180 22108 9186 22120
rect 9398 22108 9404 22120
rect 9456 22108 9462 22160
rect 10226 22148 10232 22160
rect 10187 22120 10232 22148
rect 10226 22108 10232 22120
rect 10284 22108 10290 22160
rect 11241 22151 11299 22157
rect 11241 22117 11253 22151
rect 11287 22148 11299 22151
rect 11422 22148 11428 22160
rect 11287 22120 11428 22148
rect 11287 22117 11299 22120
rect 11241 22111 11299 22117
rect 11422 22108 11428 22120
rect 11480 22108 11486 22160
rect 12066 22108 12072 22160
rect 12124 22148 12130 22160
rect 12161 22151 12219 22157
rect 12161 22148 12173 22151
rect 12124 22120 12173 22148
rect 12124 22108 12130 22120
rect 12161 22117 12173 22120
rect 12207 22117 12219 22151
rect 12161 22111 12219 22117
rect 13679 22151 13737 22157
rect 13679 22117 13691 22151
rect 13725 22148 13737 22151
rect 13906 22148 13912 22160
rect 13725 22120 13912 22148
rect 13725 22117 13737 22120
rect 13679 22111 13737 22117
rect 13906 22108 13912 22120
rect 13964 22108 13970 22160
rect 17770 22148 17776 22160
rect 14016 22120 17776 22148
rect 8389 22083 8447 22089
rect 8389 22049 8401 22083
rect 8435 22080 8447 22083
rect 8846 22080 8852 22092
rect 8435 22052 8852 22080
rect 8435 22049 8447 22052
rect 8389 22043 8447 22049
rect 8588 22024 8616 22052
rect 8846 22040 8852 22052
rect 8904 22040 8910 22092
rect 8938 22040 8944 22092
rect 8996 22080 9002 22092
rect 9766 22080 9772 22092
rect 8996 22052 9772 22080
rect 8996 22040 9002 22052
rect 9766 22040 9772 22052
rect 9824 22080 9830 22092
rect 10321 22083 10379 22089
rect 10321 22080 10333 22083
rect 9824 22052 10333 22080
rect 9824 22040 9830 22052
rect 10321 22049 10333 22052
rect 10367 22049 10379 22083
rect 10321 22043 10379 22049
rect 10870 22040 10876 22092
rect 10928 22040 10934 22092
rect 11698 22040 11704 22092
rect 11756 22080 11762 22092
rect 11977 22083 12035 22089
rect 11977 22080 11989 22083
rect 11756 22052 11989 22080
rect 11756 22040 11762 22052
rect 11977 22049 11989 22052
rect 12023 22049 12035 22083
rect 11977 22043 12035 22049
rect 13538 22040 13544 22092
rect 13596 22080 13602 22092
rect 14016 22080 14044 22120
rect 17770 22108 17776 22120
rect 17828 22108 17834 22160
rect 18340 22148 18368 22188
rect 18874 22148 18880 22160
rect 18064 22120 18368 22148
rect 18835 22120 18880 22148
rect 18064 22092 18092 22120
rect 18874 22108 18880 22120
rect 18932 22108 18938 22160
rect 13596 22052 14044 22080
rect 15289 22083 15347 22089
rect 13596 22040 13602 22052
rect 15289 22049 15301 22083
rect 15335 22080 15347 22083
rect 15378 22080 15384 22092
rect 15335 22052 15384 22080
rect 15335 22049 15347 22052
rect 15289 22043 15347 22049
rect 15378 22040 15384 22052
rect 15436 22040 15442 22092
rect 15562 22080 15568 22092
rect 15523 22052 15568 22080
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 16844 22083 16902 22089
rect 16844 22049 16856 22083
rect 16890 22080 16902 22083
rect 17126 22080 17132 22092
rect 16890 22052 17132 22080
rect 16890 22049 16902 22052
rect 16844 22043 16902 22049
rect 17126 22040 17132 22052
rect 17184 22080 17190 22092
rect 18046 22080 18052 22092
rect 17184 22052 18052 22080
rect 17184 22040 17190 22052
rect 18046 22040 18052 22052
rect 18104 22040 18110 22092
rect 18601 22083 18659 22089
rect 18601 22049 18613 22083
rect 18647 22080 18659 22083
rect 18966 22080 18972 22092
rect 18647 22052 18972 22080
rect 18647 22049 18659 22052
rect 18601 22043 18659 22049
rect 18966 22040 18972 22052
rect 19024 22080 19030 22092
rect 19150 22080 19156 22092
rect 19024 22052 19156 22080
rect 19024 22040 19030 22052
rect 19150 22040 19156 22052
rect 19208 22040 19214 22092
rect 19260 22080 19288 22188
rect 20806 22176 20812 22228
rect 20864 22216 20870 22228
rect 21450 22216 21456 22228
rect 20864 22188 21456 22216
rect 20864 22176 20870 22188
rect 21450 22176 21456 22188
rect 21508 22176 21514 22228
rect 22296 22188 23704 22216
rect 19610 22148 19616 22160
rect 19571 22120 19616 22148
rect 19610 22108 19616 22120
rect 19668 22108 19674 22160
rect 20990 22157 20996 22160
rect 20975 22151 20996 22157
rect 20975 22117 20987 22151
rect 20975 22111 20996 22117
rect 20990 22108 20996 22111
rect 21048 22108 21054 22160
rect 21269 22151 21327 22157
rect 21269 22117 21281 22151
rect 21315 22148 21327 22151
rect 22296 22148 22324 22188
rect 21315 22120 22324 22148
rect 22373 22151 22431 22157
rect 21315 22117 21327 22120
rect 21269 22111 21327 22117
rect 22373 22117 22385 22151
rect 22419 22148 22431 22151
rect 23017 22151 23075 22157
rect 23017 22148 23029 22151
rect 22419 22120 23029 22148
rect 22419 22117 22431 22120
rect 22373 22111 22431 22117
rect 23017 22117 23029 22120
rect 23063 22148 23075 22151
rect 23382 22148 23388 22160
rect 23063 22120 23388 22148
rect 23063 22117 23075 22120
rect 23017 22111 23075 22117
rect 23382 22108 23388 22120
rect 23440 22108 23446 22160
rect 23676 22148 23704 22188
rect 23750 22176 23756 22228
rect 23808 22216 23814 22228
rect 24581 22219 24639 22225
rect 24581 22216 24593 22219
rect 23808 22188 24593 22216
rect 23808 22176 23814 22188
rect 24581 22185 24593 22188
rect 24627 22185 24639 22219
rect 25774 22216 25780 22228
rect 24581 22179 24639 22185
rect 24688 22188 25780 22216
rect 24210 22148 24216 22160
rect 23676 22120 24216 22148
rect 24210 22108 24216 22120
rect 24268 22148 24274 22160
rect 24688 22148 24716 22188
rect 25774 22176 25780 22188
rect 25832 22176 25838 22228
rect 24268 22120 24716 22148
rect 24268 22108 24274 22120
rect 24762 22108 24768 22160
rect 24820 22108 24826 22160
rect 20625 22083 20683 22089
rect 19260 22052 19748 22080
rect 7892 21984 8331 22012
rect 7892 21972 7898 21984
rect 8570 21972 8576 22024
rect 8628 21972 8634 22024
rect 8665 22015 8723 22021
rect 8665 21981 8677 22015
rect 8711 22012 8723 22015
rect 9125 22015 9183 22021
rect 9125 22012 9137 22015
rect 8711 21984 9137 22012
rect 8711 21981 8723 21984
rect 8665 21975 8723 21981
rect 2590 21904 2596 21956
rect 2648 21944 2654 21956
rect 2685 21947 2743 21953
rect 2685 21944 2697 21947
rect 2648 21916 2697 21944
rect 2648 21904 2654 21916
rect 2685 21913 2697 21916
rect 2731 21913 2743 21947
rect 2685 21907 2743 21913
rect 3510 21904 3516 21956
rect 3568 21944 3574 21956
rect 3694 21944 3700 21956
rect 3568 21916 3700 21944
rect 3568 21904 3574 21916
rect 3694 21904 3700 21916
rect 3752 21904 3758 21956
rect 4154 21944 4160 21956
rect 3896 21916 4160 21944
rect 1578 21876 1584 21888
rect 1539 21848 1584 21876
rect 1578 21836 1584 21848
rect 1636 21836 1642 21888
rect 2406 21876 2412 21888
rect 2367 21848 2412 21876
rect 2406 21836 2412 21848
rect 2464 21836 2470 21888
rect 3050 21876 3056 21888
rect 3011 21848 3056 21876
rect 3050 21836 3056 21848
rect 3108 21836 3114 21888
rect 3605 21879 3663 21885
rect 3605 21845 3617 21879
rect 3651 21876 3663 21879
rect 3896 21876 3924 21916
rect 4154 21904 4160 21916
rect 4212 21904 4218 21956
rect 4982 21944 4988 21956
rect 4943 21916 4988 21944
rect 4982 21904 4988 21916
rect 5040 21904 5046 21956
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 6362 21944 6368 21956
rect 5684 21916 6368 21944
rect 5684 21904 5690 21916
rect 6362 21904 6368 21916
rect 6420 21904 6426 21956
rect 4246 21876 4252 21888
rect 3651 21848 3924 21876
rect 4207 21848 4252 21876
rect 3651 21845 3663 21848
rect 3605 21839 3663 21845
rect 4246 21836 4252 21848
rect 4304 21836 4310 21888
rect 4430 21836 4436 21888
rect 4488 21876 4494 21888
rect 4617 21879 4675 21885
rect 4617 21876 4629 21879
rect 4488 21848 4629 21876
rect 4488 21836 4494 21848
rect 4617 21845 4629 21848
rect 4663 21845 4675 21879
rect 5994 21876 6000 21888
rect 5955 21848 6000 21876
rect 4617 21839 4675 21845
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 6178 21836 6184 21888
rect 6236 21876 6242 21888
rect 8113 21879 8171 21885
rect 8113 21876 8125 21879
rect 6236 21848 8125 21876
rect 6236 21836 6242 21848
rect 8113 21845 8125 21848
rect 8159 21845 8171 21879
rect 8113 21839 8171 21845
rect 8386 21836 8392 21888
rect 8444 21876 8450 21888
rect 8772 21876 8800 21984
rect 9125 21981 9137 21984
rect 9171 22012 9183 22015
rect 9398 22012 9404 22024
rect 9171 21984 9404 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 9398 21972 9404 21984
rect 9456 21972 9462 22024
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 22012 10287 22015
rect 10502 22012 10508 22024
rect 10275 21984 10508 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 10502 21972 10508 21984
rect 10560 21972 10566 22024
rect 10888 22012 10916 22040
rect 11790 22012 11796 22024
rect 10888 21984 11796 22012
rect 11790 21972 11796 21984
rect 11848 21972 11854 22024
rect 12250 22012 12256 22024
rect 12211 21984 12256 22012
rect 12250 21972 12256 21984
rect 12308 21972 12314 22024
rect 13081 22015 13139 22021
rect 13081 21981 13093 22015
rect 13127 22012 13139 22015
rect 13722 22012 13728 22024
rect 13127 21984 13728 22012
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 13722 21972 13728 21984
rect 13780 21972 13786 22024
rect 13817 22015 13875 22021
rect 13817 21981 13829 22015
rect 13863 22012 13875 22015
rect 13998 22012 14004 22024
rect 13863 21984 14004 22012
rect 13863 21981 13875 21984
rect 13817 21975 13875 21981
rect 13998 21972 14004 21984
rect 14056 21972 14062 22024
rect 15102 22012 15108 22024
rect 15063 21984 15108 22012
rect 15102 21972 15108 21984
rect 15160 21972 15166 22024
rect 16577 22015 16635 22021
rect 16577 21981 16589 22015
rect 16623 21981 16635 22015
rect 16577 21975 16635 21981
rect 9769 21947 9827 21953
rect 9769 21913 9781 21947
rect 9815 21944 9827 21947
rect 9858 21944 9864 21956
rect 9815 21916 9864 21944
rect 9815 21913 9827 21916
rect 9769 21907 9827 21913
rect 9858 21904 9864 21916
rect 9916 21904 9922 21956
rect 11330 21904 11336 21956
rect 11388 21944 11394 21956
rect 13265 21947 13323 21953
rect 13265 21944 13277 21947
rect 11388 21916 13277 21944
rect 11388 21904 11394 21916
rect 13265 21913 13277 21916
rect 13311 21913 13323 21947
rect 13265 21907 13323 21913
rect 14737 21947 14795 21953
rect 14737 21913 14749 21947
rect 14783 21944 14795 21947
rect 16482 21944 16488 21956
rect 14783 21916 16488 21944
rect 14783 21913 14795 21916
rect 14737 21907 14795 21913
rect 16482 21904 16488 21916
rect 16540 21904 16546 21956
rect 8444 21848 8800 21876
rect 8444 21836 8450 21848
rect 9214 21836 9220 21888
rect 9272 21876 9278 21888
rect 9401 21879 9459 21885
rect 9401 21876 9413 21879
rect 9272 21848 9413 21876
rect 9272 21836 9278 21848
rect 9401 21845 9413 21848
rect 9447 21845 9459 21879
rect 10778 21876 10784 21888
rect 10739 21848 10784 21876
rect 9401 21839 9459 21845
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 11054 21836 11060 21888
rect 11112 21876 11118 21888
rect 11701 21879 11759 21885
rect 11701 21876 11713 21879
rect 11112 21848 11713 21876
rect 11112 21836 11118 21848
rect 11701 21845 11713 21848
rect 11747 21845 11759 21879
rect 12710 21876 12716 21888
rect 12671 21848 12716 21876
rect 11701 21839 11759 21845
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 14274 21876 14280 21888
rect 14235 21848 14280 21876
rect 14274 21836 14280 21848
rect 14332 21836 14338 21888
rect 15562 21836 15568 21888
rect 15620 21876 15626 21888
rect 15930 21876 15936 21888
rect 15620 21848 15936 21876
rect 15620 21836 15626 21848
rect 15930 21836 15936 21848
rect 15988 21876 15994 21888
rect 16025 21879 16083 21885
rect 16025 21876 16037 21879
rect 15988 21848 16037 21876
rect 15988 21836 15994 21848
rect 16025 21845 16037 21848
rect 16071 21845 16083 21879
rect 16592 21876 16620 21975
rect 17678 21972 17684 22024
rect 17736 22012 17742 22024
rect 18782 22012 18788 22024
rect 17736 21984 18788 22012
rect 17736 21972 17742 21984
rect 18782 21972 18788 21984
rect 18840 21972 18846 22024
rect 19518 22012 19524 22024
rect 19479 21984 19524 22012
rect 19518 21972 19524 21984
rect 19576 21972 19582 22024
rect 19720 22021 19748 22052
rect 20625 22049 20637 22083
rect 20671 22080 20683 22083
rect 20714 22080 20720 22092
rect 20671 22052 20720 22080
rect 20671 22049 20683 22052
rect 20625 22043 20683 22049
rect 20714 22040 20720 22052
rect 20772 22040 20778 22092
rect 21082 22080 21088 22092
rect 20916 22052 21088 22080
rect 20916 22024 20944 22052
rect 21082 22040 21088 22052
rect 21140 22040 21146 22092
rect 22646 22040 22652 22092
rect 22704 22080 22710 22092
rect 22704 22052 23152 22080
rect 22704 22040 22710 22052
rect 19705 22015 19763 22021
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 19889 22015 19947 22021
rect 19889 22012 19901 22015
rect 19751 21984 19901 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 19889 21981 19901 21984
rect 19935 21981 19947 22015
rect 19889 21975 19947 21981
rect 20898 21972 20904 22024
rect 20956 21972 20962 22024
rect 21545 22015 21603 22021
rect 21545 21981 21557 22015
rect 21591 21981 21603 22015
rect 21545 21975 21603 21981
rect 19153 21947 19211 21953
rect 19153 21944 19165 21947
rect 17512 21916 19165 21944
rect 17218 21876 17224 21888
rect 16592 21848 17224 21876
rect 16025 21839 16083 21845
rect 17218 21836 17224 21848
rect 17276 21836 17282 21888
rect 17310 21836 17316 21888
rect 17368 21876 17374 21888
rect 17512 21876 17540 21916
rect 19153 21913 19165 21916
rect 19199 21913 19211 21947
rect 19153 21907 19211 21913
rect 21082 21904 21088 21956
rect 21140 21944 21146 21956
rect 21560 21944 21588 21975
rect 22738 21972 22744 22024
rect 22796 22012 22802 22024
rect 23124 22021 23152 22052
rect 24118 22040 24124 22092
rect 24176 22080 24182 22092
rect 24397 22083 24455 22089
rect 24397 22080 24409 22083
rect 24176 22052 24409 22080
rect 24176 22040 24182 22052
rect 24397 22049 24409 22052
rect 24443 22049 24455 22083
rect 24780 22080 24808 22108
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 24780 22052 25053 22080
rect 24397 22043 24455 22049
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 25041 22043 25099 22049
rect 23017 22015 23075 22021
rect 23017 22012 23029 22015
rect 22796 21984 23029 22012
rect 22796 21972 22802 21984
rect 23017 21981 23029 21984
rect 23063 21981 23075 22015
rect 23017 21975 23075 21981
rect 23109 22015 23167 22021
rect 23109 21981 23121 22015
rect 23155 22012 23167 22015
rect 23474 22012 23480 22024
rect 23155 21984 23480 22012
rect 23155 21981 23167 21984
rect 23109 21975 23167 21981
rect 22554 21944 22560 21956
rect 21140 21916 21588 21944
rect 22515 21916 22560 21944
rect 21140 21904 21146 21916
rect 22554 21904 22560 21916
rect 22612 21904 22618 21956
rect 23032 21888 23060 21975
rect 23474 21972 23480 21984
rect 23532 22012 23538 22024
rect 24673 22015 24731 22021
rect 24673 22012 24685 22015
rect 23532 21984 24685 22012
rect 23532 21972 23538 21984
rect 24673 21981 24685 21984
rect 24719 22012 24731 22015
rect 24719 21984 24900 22012
rect 24719 21981 24731 21984
rect 24673 21975 24731 21981
rect 23566 21904 23572 21956
rect 23624 21944 23630 21956
rect 24121 21947 24179 21953
rect 24121 21944 24133 21947
rect 23624 21916 24133 21944
rect 23624 21904 23630 21916
rect 24121 21913 24133 21916
rect 24167 21944 24179 21947
rect 24762 21944 24768 21956
rect 24167 21916 24768 21944
rect 24167 21913 24179 21916
rect 24121 21907 24179 21913
rect 24762 21904 24768 21916
rect 24820 21904 24826 21956
rect 24872 21944 24900 21984
rect 24946 21972 24952 22024
rect 25004 22012 25010 22024
rect 25409 22015 25467 22021
rect 25409 22012 25421 22015
rect 25004 21984 25421 22012
rect 25004 21972 25010 21984
rect 25409 21981 25421 21984
rect 25455 21981 25467 22015
rect 25409 21975 25467 21981
rect 25314 21944 25320 21956
rect 24872 21916 25320 21944
rect 25314 21904 25320 21916
rect 25372 21904 25378 21956
rect 17368 21848 17540 21876
rect 19889 21879 19947 21885
rect 17368 21836 17374 21848
rect 19889 21845 19901 21879
rect 19935 21876 19947 21879
rect 20165 21879 20223 21885
rect 20165 21876 20177 21879
rect 19935 21848 20177 21876
rect 19935 21845 19947 21848
rect 19889 21839 19947 21845
rect 20165 21845 20177 21848
rect 20211 21876 20223 21879
rect 20346 21876 20352 21888
rect 20211 21848 20352 21876
rect 20211 21845 20223 21848
rect 20165 21839 20223 21845
rect 20346 21836 20352 21848
rect 20404 21836 20410 21888
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 21913 21879 21971 21885
rect 21913 21876 21925 21879
rect 21600 21848 21925 21876
rect 21600 21836 21606 21848
rect 21913 21845 21925 21848
rect 21959 21845 21971 21879
rect 21913 21839 21971 21845
rect 22278 21836 22284 21888
rect 22336 21876 22342 21888
rect 22830 21876 22836 21888
rect 22336 21848 22836 21876
rect 22336 21836 22342 21848
rect 22830 21836 22836 21848
rect 22888 21836 22894 21888
rect 23014 21836 23020 21888
rect 23072 21836 23078 21888
rect 23658 21876 23664 21888
rect 23619 21848 23664 21876
rect 23658 21836 23664 21848
rect 23716 21836 23722 21888
rect 25222 21836 25228 21888
rect 25280 21876 25286 21888
rect 25777 21879 25835 21885
rect 25777 21876 25789 21879
rect 25280 21848 25789 21876
rect 25280 21836 25286 21848
rect 25777 21845 25789 21848
rect 25823 21845 25835 21879
rect 25777 21839 25835 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1302 21632 1308 21684
rect 1360 21672 1366 21684
rect 1670 21672 1676 21684
rect 1360 21644 1676 21672
rect 1360 21632 1366 21644
rect 1670 21632 1676 21644
rect 1728 21632 1734 21684
rect 2682 21632 2688 21684
rect 2740 21672 2746 21684
rect 2961 21675 3019 21681
rect 2961 21672 2973 21675
rect 2740 21644 2973 21672
rect 2740 21632 2746 21644
rect 2961 21641 2973 21644
rect 3007 21672 3019 21675
rect 4062 21672 4068 21684
rect 3007 21644 4068 21672
rect 3007 21641 3019 21644
rect 2961 21635 3019 21641
rect 4062 21632 4068 21644
rect 4120 21632 4126 21684
rect 5261 21675 5319 21681
rect 5261 21641 5273 21675
rect 5307 21672 5319 21675
rect 5442 21672 5448 21684
rect 5307 21644 5448 21672
rect 5307 21641 5319 21644
rect 5261 21635 5319 21641
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 7742 21632 7748 21684
rect 7800 21672 7806 21684
rect 10873 21675 10931 21681
rect 7800 21644 10456 21672
rect 7800 21632 7806 21644
rect 1210 21564 1216 21616
rect 1268 21604 1274 21616
rect 1486 21604 1492 21616
rect 1268 21576 1492 21604
rect 1268 21564 1274 21576
rect 1486 21564 1492 21576
rect 1544 21564 1550 21616
rect 3694 21604 3700 21616
rect 3655 21576 3700 21604
rect 3694 21564 3700 21576
rect 3752 21564 3758 21616
rect 4985 21607 5043 21613
rect 4985 21573 4997 21607
rect 5031 21604 5043 21607
rect 5534 21604 5540 21616
rect 5031 21576 5540 21604
rect 5031 21573 5043 21576
rect 4985 21567 5043 21573
rect 5534 21564 5540 21576
rect 5592 21604 5598 21616
rect 8018 21604 8024 21616
rect 5592 21576 8024 21604
rect 5592 21564 5598 21576
rect 8018 21564 8024 21576
rect 8076 21564 8082 21616
rect 10428 21604 10456 21644
rect 10873 21641 10885 21675
rect 10919 21672 10931 21675
rect 10962 21672 10968 21684
rect 10919 21644 10968 21672
rect 10919 21641 10931 21644
rect 10873 21635 10931 21641
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 11609 21675 11667 21681
rect 11609 21641 11621 21675
rect 11655 21672 11667 21675
rect 12710 21672 12716 21684
rect 11655 21644 12716 21672
rect 11655 21641 11667 21644
rect 11609 21635 11667 21641
rect 12710 21632 12716 21644
rect 12768 21632 12774 21684
rect 13354 21632 13360 21684
rect 13412 21672 13418 21684
rect 13630 21672 13636 21684
rect 13412 21644 13636 21672
rect 13412 21632 13418 21644
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 13814 21672 13820 21684
rect 13775 21644 13820 21672
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 15197 21675 15255 21681
rect 15197 21641 15209 21675
rect 15243 21672 15255 21675
rect 15378 21672 15384 21684
rect 15243 21644 15384 21672
rect 15243 21641 15255 21644
rect 15197 21635 15255 21641
rect 15378 21632 15384 21644
rect 15436 21632 15442 21684
rect 15473 21675 15531 21681
rect 15473 21641 15485 21675
rect 15519 21672 15531 21675
rect 15654 21672 15660 21684
rect 15519 21644 15660 21672
rect 15519 21641 15531 21644
rect 15473 21635 15531 21641
rect 15654 21632 15660 21644
rect 15712 21632 15718 21684
rect 16482 21672 16488 21684
rect 16443 21644 16488 21672
rect 16482 21632 16488 21644
rect 16540 21632 16546 21684
rect 16942 21632 16948 21684
rect 17000 21672 17006 21684
rect 17126 21672 17132 21684
rect 17000 21644 17132 21672
rect 17000 21632 17006 21644
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 17218 21632 17224 21684
rect 17276 21672 17282 21684
rect 17494 21672 17500 21684
rect 17276 21644 17500 21672
rect 17276 21632 17282 21644
rect 17494 21632 17500 21644
rect 17552 21672 17558 21684
rect 17589 21675 17647 21681
rect 17589 21672 17601 21675
rect 17552 21644 17601 21672
rect 17552 21632 17558 21644
rect 17589 21641 17601 21644
rect 17635 21641 17647 21675
rect 17589 21635 17647 21641
rect 17862 21632 17868 21684
rect 17920 21672 17926 21684
rect 18233 21675 18291 21681
rect 18233 21672 18245 21675
rect 17920 21644 18245 21672
rect 17920 21632 17926 21644
rect 18233 21641 18245 21644
rect 18279 21641 18291 21675
rect 18233 21635 18291 21641
rect 11422 21604 11428 21616
rect 10428 21576 11428 21604
rect 11422 21564 11428 21576
rect 11480 21564 11486 21616
rect 15930 21564 15936 21616
rect 15988 21604 15994 21616
rect 16114 21604 16120 21616
rect 15988 21576 16120 21604
rect 15988 21564 15994 21576
rect 16114 21564 16120 21576
rect 16172 21564 16178 21616
rect 2038 21536 2044 21548
rect 1999 21508 2044 21536
rect 2038 21496 2044 21508
rect 2096 21496 2102 21548
rect 2222 21496 2228 21548
rect 2280 21536 2286 21548
rect 5626 21536 5632 21548
rect 2280 21508 5632 21536
rect 2280 21496 2286 21508
rect 5626 21496 5632 21508
rect 5684 21496 5690 21548
rect 8036 21536 8064 21564
rect 8036 21508 8340 21536
rect 1765 21471 1823 21477
rect 1765 21437 1777 21471
rect 1811 21468 1823 21471
rect 2406 21468 2412 21480
rect 1811 21440 2412 21468
rect 1811 21437 1823 21440
rect 1765 21431 1823 21437
rect 2406 21428 2412 21440
rect 2464 21428 2470 21480
rect 3513 21471 3571 21477
rect 3513 21437 3525 21471
rect 3559 21468 3571 21471
rect 6914 21468 6920 21480
rect 3559 21440 4292 21468
rect 6875 21440 6920 21468
rect 3559 21437 3571 21440
rect 3513 21431 3571 21437
rect 3973 21403 4031 21409
rect 3973 21369 3985 21403
rect 4019 21400 4031 21403
rect 4062 21400 4068 21412
rect 4019 21372 4068 21400
rect 4019 21369 4031 21372
rect 3973 21363 4031 21369
rect 4062 21360 4068 21372
rect 4120 21360 4126 21412
rect 4264 21409 4292 21440
rect 6914 21428 6920 21440
rect 6972 21428 6978 21480
rect 8202 21468 8208 21480
rect 8036 21440 8208 21468
rect 4249 21403 4307 21409
rect 4249 21369 4261 21403
rect 4295 21400 4307 21403
rect 4522 21400 4528 21412
rect 4295 21372 4528 21400
rect 4295 21369 4307 21372
rect 4249 21363 4307 21369
rect 4522 21360 4528 21372
rect 4580 21360 4586 21412
rect 5166 21360 5172 21412
rect 5224 21400 5230 21412
rect 5534 21400 5540 21412
rect 5224 21372 5540 21400
rect 5224 21360 5230 21372
rect 5534 21360 5540 21372
rect 5592 21360 5598 21412
rect 5810 21400 5816 21412
rect 5771 21372 5816 21400
rect 5810 21360 5816 21372
rect 5868 21360 5874 21412
rect 5994 21360 6000 21412
rect 6052 21400 6058 21412
rect 6457 21403 6515 21409
rect 6457 21400 6469 21403
rect 6052 21372 6469 21400
rect 6052 21360 6058 21372
rect 6457 21369 6469 21372
rect 6503 21400 6515 21403
rect 7006 21400 7012 21412
rect 6503 21372 7012 21400
rect 6503 21369 6515 21372
rect 6457 21363 6515 21369
rect 7006 21360 7012 21372
rect 7064 21360 7070 21412
rect 7190 21400 7196 21412
rect 7151 21372 7196 21400
rect 7190 21360 7196 21372
rect 7248 21360 7254 21412
rect 7745 21403 7803 21409
rect 7745 21369 7757 21403
rect 7791 21400 7803 21403
rect 7834 21400 7840 21412
rect 7791 21372 7840 21400
rect 7791 21369 7803 21372
rect 7745 21363 7803 21369
rect 7834 21360 7840 21372
rect 7892 21360 7898 21412
rect 1673 21335 1731 21341
rect 1673 21301 1685 21335
rect 1719 21332 1731 21335
rect 1854 21332 1860 21344
rect 1719 21304 1860 21332
rect 1719 21301 1731 21304
rect 1673 21295 1731 21301
rect 1854 21292 1860 21304
rect 1912 21292 1918 21344
rect 2590 21332 2596 21344
rect 2551 21304 2596 21332
rect 2590 21292 2596 21304
rect 2648 21292 2654 21344
rect 4154 21332 4160 21344
rect 4115 21304 4160 21332
rect 4154 21292 4160 21304
rect 4212 21292 4218 21344
rect 5350 21292 5356 21344
rect 5408 21332 5414 21344
rect 5721 21335 5779 21341
rect 5721 21332 5733 21335
rect 5408 21304 5733 21332
rect 5408 21292 5414 21304
rect 5721 21301 5733 21304
rect 5767 21301 5779 21335
rect 5721 21295 5779 21301
rect 6638 21292 6644 21344
rect 6696 21332 6702 21344
rect 8036 21341 8064 21440
rect 8202 21428 8208 21440
rect 8260 21428 8266 21480
rect 8312 21468 8340 21508
rect 10962 21496 10968 21548
rect 11020 21536 11026 21548
rect 11333 21539 11391 21545
rect 11333 21536 11345 21539
rect 11020 21508 11345 21536
rect 11020 21496 11026 21508
rect 11333 21505 11345 21508
rect 11379 21536 11391 21539
rect 11974 21536 11980 21548
rect 11379 21508 11980 21536
rect 11379 21505 11391 21508
rect 11333 21499 11391 21505
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 14461 21539 14519 21545
rect 14461 21505 14473 21539
rect 14507 21536 14519 21539
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 14507 21508 16865 21536
rect 14507 21505 14519 21508
rect 14461 21499 14519 21505
rect 16853 21505 16865 21508
rect 16899 21536 16911 21539
rect 18138 21536 18144 21548
rect 16899 21508 18144 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 18138 21496 18144 21508
rect 18196 21496 18202 21548
rect 18248 21536 18276 21635
rect 21818 21632 21824 21684
rect 21876 21672 21882 21684
rect 22094 21672 22100 21684
rect 21876 21644 22100 21672
rect 21876 21632 21882 21644
rect 22094 21632 22100 21644
rect 22152 21632 22158 21684
rect 22557 21675 22615 21681
rect 22557 21641 22569 21675
rect 22603 21672 22615 21675
rect 22646 21672 22652 21684
rect 22603 21644 22652 21672
rect 22603 21641 22615 21644
rect 22557 21635 22615 21641
rect 22646 21632 22652 21644
rect 22704 21632 22710 21684
rect 23753 21675 23811 21681
rect 23753 21641 23765 21675
rect 23799 21672 23811 21675
rect 24762 21672 24768 21684
rect 23799 21644 24768 21672
rect 23799 21641 23811 21644
rect 23753 21635 23811 21641
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 26326 21672 26332 21684
rect 26287 21644 26332 21672
rect 26326 21632 26332 21644
rect 26384 21632 26390 21684
rect 21361 21607 21419 21613
rect 21361 21573 21373 21607
rect 21407 21604 21419 21607
rect 22830 21604 22836 21616
rect 21407 21576 22836 21604
rect 21407 21573 21419 21576
rect 21361 21567 21419 21573
rect 22830 21564 22836 21576
rect 22888 21564 22894 21616
rect 21818 21536 21824 21548
rect 18248 21508 18920 21536
rect 21779 21508 21824 21536
rect 8461 21471 8519 21477
rect 8461 21468 8473 21471
rect 8312 21440 8473 21468
rect 8461 21437 8473 21440
rect 8507 21437 8519 21471
rect 8461 21431 8519 21437
rect 10045 21471 10103 21477
rect 10045 21437 10057 21471
rect 10091 21468 10103 21471
rect 10226 21468 10232 21480
rect 10091 21440 10232 21468
rect 10091 21437 10103 21440
rect 10045 21431 10103 21437
rect 10226 21428 10232 21440
rect 10284 21428 10290 21480
rect 12161 21471 12219 21477
rect 12161 21437 12173 21471
rect 12207 21468 12219 21471
rect 12342 21468 12348 21480
rect 12207 21440 12348 21468
rect 12207 21437 12219 21440
rect 12161 21431 12219 21437
rect 12342 21428 12348 21440
rect 12400 21468 12406 21480
rect 12710 21477 12716 21480
rect 12437 21471 12495 21477
rect 12437 21468 12449 21471
rect 12400 21440 12449 21468
rect 12400 21428 12406 21440
rect 12437 21437 12449 21440
rect 12483 21437 12495 21471
rect 12704 21468 12716 21477
rect 12623 21440 12716 21468
rect 12437 21431 12495 21437
rect 12704 21431 12716 21440
rect 12768 21468 12774 21480
rect 13446 21468 13452 21480
rect 12768 21440 13452 21468
rect 12710 21428 12716 21431
rect 12768 21428 12774 21440
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 14826 21468 14832 21480
rect 14787 21440 14832 21468
rect 14826 21428 14832 21440
rect 14884 21428 14890 21480
rect 15289 21471 15347 21477
rect 15289 21437 15301 21471
rect 15335 21468 15347 21471
rect 16301 21471 16359 21477
rect 15335 21440 15976 21468
rect 15335 21437 15347 21440
rect 15289 21431 15347 21437
rect 9858 21360 9864 21412
rect 9916 21400 9922 21412
rect 10502 21400 10508 21412
rect 9916 21372 10508 21400
rect 9916 21360 9922 21372
rect 10502 21360 10508 21372
rect 10560 21360 10566 21412
rect 11330 21400 11336 21412
rect 11291 21372 11336 21400
rect 11330 21360 11336 21372
rect 11388 21360 11394 21412
rect 11425 21403 11483 21409
rect 11425 21369 11437 21403
rect 11471 21400 11483 21403
rect 11609 21403 11667 21409
rect 11609 21400 11621 21403
rect 11471 21372 11621 21400
rect 11471 21369 11483 21372
rect 11425 21363 11483 21369
rect 11609 21369 11621 21372
rect 11655 21369 11667 21403
rect 11609 21363 11667 21369
rect 8021 21335 8079 21341
rect 8021 21332 8033 21335
rect 6696 21304 8033 21332
rect 6696 21292 6702 21304
rect 8021 21301 8033 21304
rect 8067 21301 8079 21335
rect 8021 21295 8079 21301
rect 9490 21292 9496 21344
rect 9548 21332 9554 21344
rect 9585 21335 9643 21341
rect 9585 21332 9597 21335
rect 9548 21304 9597 21332
rect 9548 21292 9554 21304
rect 9585 21301 9597 21304
rect 9631 21301 9643 21335
rect 10042 21332 10048 21344
rect 9955 21304 10048 21332
rect 9585 21295 9643 21301
rect 10042 21292 10048 21304
rect 10100 21332 10106 21344
rect 10137 21335 10195 21341
rect 10137 21332 10149 21335
rect 10100 21304 10149 21332
rect 10100 21292 10106 21304
rect 10137 21301 10149 21304
rect 10183 21301 10195 21335
rect 10137 21295 10195 21301
rect 10778 21292 10784 21344
rect 10836 21332 10842 21344
rect 11440 21332 11468 21363
rect 10836 21304 11468 21332
rect 11885 21335 11943 21341
rect 10836 21292 10842 21304
rect 11885 21301 11897 21335
rect 11931 21332 11943 21335
rect 11974 21332 11980 21344
rect 11931 21304 11980 21332
rect 11931 21301 11943 21304
rect 11885 21295 11943 21301
rect 11974 21292 11980 21304
rect 12032 21292 12038 21344
rect 15948 21341 15976 21440
rect 16301 21437 16313 21471
rect 16347 21468 16359 21471
rect 16574 21468 16580 21480
rect 16347 21440 16580 21468
rect 16347 21437 16359 21440
rect 16301 21431 16359 21437
rect 16574 21428 16580 21440
rect 16632 21468 16638 21480
rect 16942 21468 16948 21480
rect 16632 21440 16948 21468
rect 16632 21428 16638 21440
rect 16942 21428 16948 21440
rect 17000 21428 17006 21480
rect 17037 21471 17095 21477
rect 17037 21437 17049 21471
rect 17083 21468 17095 21471
rect 17494 21468 17500 21480
rect 17083 21440 17500 21468
rect 17083 21437 17095 21440
rect 17037 21431 17095 21437
rect 17494 21428 17500 21440
rect 17552 21468 17558 21480
rect 17865 21471 17923 21477
rect 17865 21468 17877 21471
rect 17552 21440 17877 21468
rect 17552 21428 17558 21440
rect 17865 21437 17877 21440
rect 17911 21468 17923 21471
rect 18230 21468 18236 21480
rect 17911 21440 18236 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 18230 21428 18236 21440
rect 18288 21428 18294 21480
rect 18785 21471 18843 21477
rect 18785 21437 18797 21471
rect 18831 21437 18843 21471
rect 18892 21468 18920 21508
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 22152 21508 23397 21536
rect 22152 21496 22158 21508
rect 23385 21505 23397 21508
rect 23431 21536 23443 21539
rect 23750 21536 23756 21548
rect 23431 21508 23756 21536
rect 23431 21505 23443 21508
rect 23385 21499 23443 21505
rect 23750 21496 23756 21508
rect 23808 21496 23814 21548
rect 24026 21496 24032 21548
rect 24084 21536 24090 21548
rect 24213 21539 24271 21545
rect 24213 21536 24225 21539
rect 24084 21508 24225 21536
rect 24084 21496 24090 21508
rect 24213 21505 24225 21508
rect 24259 21536 24271 21539
rect 25038 21536 25044 21548
rect 24259 21508 25044 21536
rect 24259 21505 24271 21508
rect 24213 21499 24271 21505
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 19041 21471 19099 21477
rect 19041 21468 19053 21471
rect 18892 21440 19053 21468
rect 18785 21431 18843 21437
rect 19041 21437 19053 21440
rect 19087 21468 19099 21471
rect 19334 21468 19340 21480
rect 19087 21440 19340 21468
rect 19087 21437 19099 21440
rect 19041 21431 19099 21437
rect 16758 21360 16764 21412
rect 16816 21400 16822 21412
rect 17126 21400 17132 21412
rect 16816 21372 17132 21400
rect 16816 21360 16822 21372
rect 17126 21360 17132 21372
rect 17184 21360 17190 21412
rect 17405 21403 17463 21409
rect 17405 21369 17417 21403
rect 17451 21400 17463 21403
rect 17589 21403 17647 21409
rect 17589 21400 17601 21403
rect 17451 21372 17601 21400
rect 17451 21369 17463 21372
rect 17405 21363 17463 21369
rect 17589 21369 17601 21372
rect 17635 21400 17647 21403
rect 18693 21403 18751 21409
rect 18693 21400 18705 21403
rect 17635 21372 18705 21400
rect 17635 21369 17647 21372
rect 17589 21363 17647 21369
rect 18693 21369 18705 21372
rect 18739 21400 18751 21403
rect 18800 21400 18828 21431
rect 19334 21428 19340 21440
rect 19392 21428 19398 21480
rect 21542 21428 21548 21480
rect 21600 21468 21606 21480
rect 21913 21471 21971 21477
rect 21913 21468 21925 21471
rect 21600 21440 21925 21468
rect 21600 21428 21606 21440
rect 21913 21437 21925 21440
rect 21959 21437 21971 21471
rect 21913 21431 21971 21437
rect 22370 21428 22376 21480
rect 22428 21468 22434 21480
rect 24118 21468 24124 21480
rect 22428 21440 24124 21468
rect 22428 21428 22434 21440
rect 24118 21428 24124 21440
rect 24176 21468 24182 21480
rect 24673 21471 24731 21477
rect 24673 21468 24685 21471
rect 24176 21440 24685 21468
rect 24176 21428 24182 21440
rect 24673 21437 24685 21440
rect 24719 21437 24731 21471
rect 25222 21468 25228 21480
rect 25183 21440 25228 21468
rect 24673 21431 24731 21437
rect 20898 21400 20904 21412
rect 18739 21372 20904 21400
rect 18739 21369 18751 21372
rect 18693 21363 18751 21369
rect 20898 21360 20904 21372
rect 20956 21360 20962 21412
rect 22922 21360 22928 21412
rect 22980 21400 22986 21412
rect 24026 21400 24032 21412
rect 22980 21372 24032 21400
rect 22980 21360 22986 21372
rect 24026 21360 24032 21372
rect 24084 21400 24090 21412
rect 24305 21403 24363 21409
rect 24305 21400 24317 21403
rect 24084 21372 24317 21400
rect 24084 21360 24090 21372
rect 24305 21369 24317 21372
rect 24351 21369 24363 21403
rect 24688 21400 24716 21431
rect 25222 21428 25228 21440
rect 25280 21428 25286 21480
rect 26142 21468 26148 21480
rect 25332 21440 26148 21468
rect 25332 21400 25360 21440
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 25498 21400 25504 21412
rect 24688 21372 25360 21400
rect 25459 21372 25504 21400
rect 24305 21363 24363 21369
rect 25498 21360 25504 21372
rect 25556 21360 25562 21412
rect 15933 21335 15991 21341
rect 15933 21301 15945 21335
rect 15979 21332 15991 21335
rect 16114 21332 16120 21344
rect 15979 21304 16120 21332
rect 15979 21301 15991 21304
rect 15933 21295 15991 21301
rect 16114 21292 16120 21304
rect 16172 21292 16178 21344
rect 16945 21335 17003 21341
rect 16945 21301 16957 21335
rect 16991 21332 17003 21335
rect 17034 21332 17040 21344
rect 16991 21304 17040 21332
rect 16991 21301 17003 21304
rect 16945 21295 17003 21301
rect 17034 21292 17040 21304
rect 17092 21292 17098 21344
rect 19978 21292 19984 21344
rect 20036 21332 20042 21344
rect 20165 21335 20223 21341
rect 20165 21332 20177 21335
rect 20036 21304 20177 21332
rect 20036 21292 20042 21304
rect 20165 21301 20177 21304
rect 20211 21301 20223 21335
rect 20165 21295 20223 21301
rect 20346 21292 20352 21344
rect 20404 21332 20410 21344
rect 20993 21335 21051 21341
rect 20993 21332 21005 21335
rect 20404 21304 21005 21332
rect 20404 21292 20410 21304
rect 20993 21301 21005 21304
rect 21039 21332 21051 21335
rect 21542 21332 21548 21344
rect 21039 21304 21548 21332
rect 21039 21301 21051 21304
rect 20993 21295 21051 21301
rect 21542 21292 21548 21304
rect 21600 21292 21606 21344
rect 21821 21335 21879 21341
rect 21821 21301 21833 21335
rect 21867 21332 21879 21335
rect 22094 21332 22100 21344
rect 21867 21304 22100 21332
rect 21867 21301 21879 21304
rect 21821 21295 21879 21301
rect 22094 21292 22100 21304
rect 22152 21292 22158 21344
rect 22646 21292 22652 21344
rect 22704 21332 22710 21344
rect 23109 21335 23167 21341
rect 23109 21332 23121 21335
rect 22704 21304 23121 21332
rect 22704 21292 22710 21304
rect 23109 21301 23121 21304
rect 23155 21332 23167 21335
rect 24213 21335 24271 21341
rect 24213 21332 24225 21335
rect 23155 21304 24225 21332
rect 23155 21301 23167 21304
rect 23109 21295 23167 21301
rect 24213 21301 24225 21304
rect 24259 21301 24271 21335
rect 24213 21295 24271 21301
rect 25133 21335 25191 21341
rect 25133 21301 25145 21335
rect 25179 21332 25191 21335
rect 25314 21332 25320 21344
rect 25179 21304 25320 21332
rect 25179 21301 25191 21304
rect 25133 21295 25191 21301
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 25958 21332 25964 21344
rect 25919 21304 25964 21332
rect 25958 21292 25964 21304
rect 26016 21292 26022 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1762 21088 1768 21140
rect 1820 21128 1826 21140
rect 2038 21128 2044 21140
rect 1820 21100 2044 21128
rect 1820 21088 1826 21100
rect 2038 21088 2044 21100
rect 2096 21088 2102 21140
rect 2961 21131 3019 21137
rect 2961 21097 2973 21131
rect 3007 21128 3019 21131
rect 3007 21100 3464 21128
rect 3007 21097 3019 21100
rect 2961 21091 3019 21097
rect 2774 21020 2780 21072
rect 2832 21060 2838 21072
rect 3053 21063 3111 21069
rect 2832 21032 2877 21060
rect 2832 21020 2838 21032
rect 3053 21029 3065 21063
rect 3099 21060 3111 21063
rect 3326 21060 3332 21072
rect 3099 21032 3332 21060
rect 3099 21029 3111 21032
rect 3053 21023 3111 21029
rect 1946 20952 1952 21004
rect 2004 20992 2010 21004
rect 2222 20992 2228 21004
rect 2004 20964 2228 20992
rect 2004 20952 2010 20964
rect 2222 20952 2228 20964
rect 2280 20952 2286 21004
rect 3068 20924 3096 21023
rect 3326 21020 3332 21032
rect 3384 21020 3390 21072
rect 2056 20896 3096 20924
rect 1762 20788 1768 20800
rect 1723 20760 1768 20788
rect 1762 20748 1768 20760
rect 1820 20748 1826 20800
rect 1946 20748 1952 20800
rect 2004 20788 2010 20800
rect 2056 20797 2084 20896
rect 3326 20884 3332 20936
rect 3384 20924 3390 20936
rect 3436 20924 3464 21100
rect 4982 21088 4988 21140
rect 5040 21128 5046 21140
rect 5629 21131 5687 21137
rect 5629 21128 5641 21131
rect 5040 21100 5641 21128
rect 5040 21088 5046 21100
rect 5629 21097 5641 21100
rect 5675 21128 5687 21131
rect 6454 21128 6460 21140
rect 5675 21100 6460 21128
rect 5675 21097 5687 21100
rect 5629 21091 5687 21097
rect 6454 21088 6460 21100
rect 6512 21088 6518 21140
rect 6549 21131 6607 21137
rect 6549 21097 6561 21131
rect 6595 21128 6607 21131
rect 7098 21128 7104 21140
rect 6595 21100 7104 21128
rect 6595 21097 6607 21100
rect 6549 21091 6607 21097
rect 7098 21088 7104 21100
rect 7156 21128 7162 21140
rect 7742 21128 7748 21140
rect 7156 21100 7748 21128
rect 7156 21088 7162 21100
rect 7742 21088 7748 21100
rect 7800 21088 7806 21140
rect 8018 21128 8024 21140
rect 7979 21100 8024 21128
rect 8018 21088 8024 21100
rect 8076 21128 8082 21140
rect 8941 21131 8999 21137
rect 8941 21128 8953 21131
rect 8076 21100 8953 21128
rect 8076 21088 8082 21100
rect 8941 21097 8953 21100
rect 8987 21097 8999 21131
rect 8941 21091 8999 21097
rect 9493 21131 9551 21137
rect 9493 21097 9505 21131
rect 9539 21128 9551 21131
rect 9766 21128 9772 21140
rect 9539 21100 9772 21128
rect 9539 21097 9551 21100
rect 9493 21091 9551 21097
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 11054 21128 11060 21140
rect 11015 21100 11060 21128
rect 11054 21088 11060 21100
rect 11112 21088 11118 21140
rect 12069 21131 12127 21137
rect 12069 21097 12081 21131
rect 12115 21128 12127 21131
rect 12250 21128 12256 21140
rect 12115 21100 12256 21128
rect 12115 21097 12127 21100
rect 12069 21091 12127 21097
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 13906 21128 13912 21140
rect 13867 21100 13912 21128
rect 13906 21088 13912 21100
rect 13964 21088 13970 21140
rect 14277 21131 14335 21137
rect 14277 21097 14289 21131
rect 14323 21128 14335 21131
rect 14366 21128 14372 21140
rect 14323 21100 14372 21128
rect 14323 21097 14335 21100
rect 14277 21091 14335 21097
rect 14366 21088 14372 21100
rect 14424 21088 14430 21140
rect 15010 21128 15016 21140
rect 14971 21100 15016 21128
rect 15010 21088 15016 21100
rect 15068 21088 15074 21140
rect 15838 21128 15844 21140
rect 15799 21100 15844 21128
rect 15838 21088 15844 21100
rect 15896 21088 15902 21140
rect 16485 21131 16543 21137
rect 16485 21097 16497 21131
rect 16531 21128 16543 21131
rect 16758 21128 16764 21140
rect 16531 21100 16764 21128
rect 16531 21097 16543 21100
rect 16485 21091 16543 21097
rect 16758 21088 16764 21100
rect 16816 21128 16822 21140
rect 19521 21131 19579 21137
rect 16816 21100 17540 21128
rect 16816 21088 16822 21100
rect 17512 21072 17540 21100
rect 19521 21097 19533 21131
rect 19567 21128 19579 21131
rect 20346 21128 20352 21140
rect 19567 21100 20352 21128
rect 19567 21097 19579 21100
rect 19521 21091 19579 21097
rect 20346 21088 20352 21100
rect 20404 21088 20410 21140
rect 21358 21088 21364 21140
rect 21416 21128 21422 21140
rect 21453 21131 21511 21137
rect 21453 21128 21465 21131
rect 21416 21100 21465 21128
rect 21416 21088 21422 21100
rect 21453 21097 21465 21100
rect 21499 21097 21511 21131
rect 21453 21091 21511 21097
rect 22922 21088 22928 21140
rect 22980 21128 22986 21140
rect 23198 21128 23204 21140
rect 22980 21100 23204 21128
rect 22980 21088 22986 21100
rect 23198 21088 23204 21100
rect 23256 21088 23262 21140
rect 24854 21088 24860 21140
rect 24912 21128 24918 21140
rect 25409 21131 25467 21137
rect 25409 21128 25421 21131
rect 24912 21100 25421 21128
rect 24912 21088 24918 21100
rect 25409 21097 25421 21100
rect 25455 21097 25467 21131
rect 25409 21091 25467 21097
rect 25774 21088 25780 21140
rect 25832 21128 25838 21140
rect 26145 21131 26203 21137
rect 26145 21128 26157 21131
rect 25832 21100 26157 21128
rect 25832 21088 25838 21100
rect 26145 21097 26157 21100
rect 26191 21097 26203 21131
rect 26145 21091 26203 21097
rect 5258 21020 5264 21072
rect 5316 21060 5322 21072
rect 5442 21060 5448 21072
rect 5316 21032 5448 21060
rect 5316 21020 5322 21032
rect 5442 21020 5448 21032
rect 5500 21020 5506 21072
rect 8570 21060 8576 21072
rect 8531 21032 8576 21060
rect 8570 21020 8576 21032
rect 8628 21020 8634 21072
rect 9674 21020 9680 21072
rect 9732 21060 9738 21072
rect 9922 21063 9980 21069
rect 9922 21060 9934 21063
rect 9732 21032 9934 21060
rect 9732 21020 9738 21032
rect 9922 21029 9934 21032
rect 9968 21029 9980 21063
rect 9922 21023 9980 21029
rect 13081 21063 13139 21069
rect 13081 21029 13093 21063
rect 13127 21060 13139 21063
rect 13127 21032 14320 21060
rect 13127 21029 13139 21032
rect 13081 21023 13139 21029
rect 14292 21004 14320 21032
rect 14826 21020 14832 21072
rect 14884 21060 14890 21072
rect 15657 21063 15715 21069
rect 15657 21060 15669 21063
rect 14884 21032 15669 21060
rect 14884 21020 14890 21032
rect 15657 21029 15669 21032
rect 15703 21060 15715 21063
rect 15746 21060 15752 21072
rect 15703 21032 15752 21060
rect 15703 21029 15715 21032
rect 15657 21023 15715 21029
rect 15746 21020 15752 21032
rect 15804 21020 15810 21072
rect 16298 21020 16304 21072
rect 16356 21060 16362 21072
rect 17221 21063 17279 21069
rect 17221 21060 17233 21063
rect 16356 21032 17233 21060
rect 16356 21020 16362 21032
rect 17221 21029 17233 21032
rect 17267 21029 17279 21063
rect 17221 21023 17279 21029
rect 17310 21020 17316 21072
rect 17368 21069 17374 21072
rect 17368 21063 17417 21069
rect 17368 21029 17371 21063
rect 17405 21029 17417 21063
rect 17494 21060 17500 21072
rect 17455 21032 17500 21060
rect 17368 21023 17417 21029
rect 17368 21020 17374 21023
rect 17494 21020 17500 21032
rect 17552 21020 17558 21072
rect 18966 21060 18972 21072
rect 18927 21032 18972 21060
rect 18966 21020 18972 21032
rect 19024 21020 19030 21072
rect 20073 21063 20131 21069
rect 20073 21029 20085 21063
rect 20119 21060 20131 21063
rect 20530 21060 20536 21072
rect 20119 21032 20536 21060
rect 20119 21029 20131 21032
rect 20073 21023 20131 21029
rect 20530 21020 20536 21032
rect 20588 21060 20594 21072
rect 21082 21060 21088 21072
rect 20588 21032 21088 21060
rect 20588 21020 20594 21032
rect 21082 21020 21088 21032
rect 21140 21020 21146 21072
rect 21542 21060 21548 21072
rect 21503 21032 21548 21060
rect 21542 21020 21548 21032
rect 21600 21020 21606 21072
rect 23017 21063 23075 21069
rect 23017 21029 23029 21063
rect 23063 21060 23075 21063
rect 23750 21060 23756 21072
rect 23063 21032 23756 21060
rect 23063 21029 23075 21032
rect 23017 21023 23075 21029
rect 23750 21020 23756 21032
rect 23808 21020 23814 21072
rect 24581 21063 24639 21069
rect 24581 21029 24593 21063
rect 24627 21060 24639 21063
rect 24670 21060 24676 21072
rect 24627 21032 24676 21060
rect 24627 21029 24639 21032
rect 24581 21023 24639 21029
rect 24670 21020 24676 21032
rect 24728 21020 24734 21072
rect 25038 21060 25044 21072
rect 24999 21032 25044 21060
rect 25038 21020 25044 21032
rect 25096 21020 25102 21072
rect 3697 20995 3755 21001
rect 3697 20961 3709 20995
rect 3743 20992 3755 20995
rect 4246 20992 4252 21004
rect 3743 20964 4252 20992
rect 3743 20961 3755 20964
rect 3697 20955 3755 20961
rect 4246 20952 4252 20964
rect 4304 20992 4310 21004
rect 5810 20992 5816 21004
rect 4304 20964 5816 20992
rect 4304 20952 4310 20964
rect 5810 20952 5816 20964
rect 5868 20992 5874 21004
rect 6181 20995 6239 21001
rect 6181 20992 6193 20995
rect 5868 20964 6193 20992
rect 5868 20952 5874 20964
rect 6181 20961 6193 20964
rect 6227 20992 6239 20995
rect 6908 20995 6966 21001
rect 6908 20992 6920 20995
rect 6227 20964 6920 20992
rect 6227 20961 6239 20964
rect 6181 20955 6239 20961
rect 6908 20961 6920 20964
rect 6954 20992 6966 20995
rect 7282 20992 7288 21004
rect 6954 20964 7288 20992
rect 6954 20961 6966 20964
rect 6908 20955 6966 20961
rect 7282 20952 7288 20964
rect 7340 20952 7346 21004
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 12897 20995 12955 21001
rect 12897 20992 12909 20995
rect 12492 20964 12909 20992
rect 12492 20952 12498 20964
rect 12897 20961 12909 20964
rect 12943 20992 12955 20995
rect 13538 20992 13544 21004
rect 12943 20964 13544 20992
rect 12943 20961 12955 20964
rect 12897 20955 12955 20961
rect 13538 20952 13544 20964
rect 13596 20952 13602 21004
rect 14093 20995 14151 21001
rect 14093 20961 14105 20995
rect 14139 20961 14151 20995
rect 14093 20955 14151 20961
rect 4062 20924 4068 20936
rect 3384 20896 3464 20924
rect 4023 20896 4068 20924
rect 3384 20884 3390 20896
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 5442 20884 5448 20936
rect 5500 20924 5506 20936
rect 5537 20927 5595 20933
rect 5537 20924 5549 20927
rect 5500 20896 5549 20924
rect 5500 20884 5506 20896
rect 5537 20893 5549 20896
rect 5583 20893 5595 20927
rect 5537 20887 5595 20893
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20924 5779 20927
rect 5994 20924 6000 20936
rect 5767 20896 6000 20924
rect 5767 20893 5779 20896
rect 5721 20887 5779 20893
rect 5169 20859 5227 20865
rect 5169 20856 5181 20859
rect 4172 20828 5181 20856
rect 2041 20791 2099 20797
rect 2041 20788 2053 20791
rect 2004 20760 2053 20788
rect 2004 20748 2010 20760
rect 2041 20757 2053 20760
rect 2087 20757 2099 20791
rect 2041 20751 2099 20757
rect 2501 20791 2559 20797
rect 2501 20757 2513 20791
rect 2547 20788 2559 20791
rect 2682 20788 2688 20800
rect 2547 20760 2688 20788
rect 2547 20757 2559 20760
rect 2501 20751 2559 20757
rect 2682 20748 2688 20760
rect 2740 20748 2746 20800
rect 3050 20748 3056 20800
rect 3108 20788 3114 20800
rect 3326 20788 3332 20800
rect 3108 20760 3332 20788
rect 3108 20748 3114 20760
rect 3326 20748 3332 20760
rect 3384 20748 3390 20800
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 4172 20788 4200 20828
rect 5169 20825 5181 20828
rect 5215 20825 5227 20859
rect 5169 20819 5227 20825
rect 4120 20760 4200 20788
rect 4120 20748 4126 20760
rect 4430 20748 4436 20800
rect 4488 20788 4494 20800
rect 4525 20791 4583 20797
rect 4525 20788 4537 20791
rect 4488 20760 4537 20788
rect 4488 20748 4494 20760
rect 4525 20757 4537 20760
rect 4571 20757 4583 20791
rect 4525 20751 4583 20757
rect 4985 20791 5043 20797
rect 4985 20757 4997 20791
rect 5031 20788 5043 20791
rect 5736 20788 5764 20887
rect 5994 20884 6000 20896
rect 6052 20884 6058 20936
rect 6638 20924 6644 20936
rect 6599 20896 6644 20924
rect 6638 20884 6644 20896
rect 6696 20884 6702 20936
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 11698 20924 11704 20936
rect 9732 20896 9777 20924
rect 11659 20896 11704 20924
rect 9732 20884 9738 20896
rect 11698 20884 11704 20896
rect 11756 20884 11762 20936
rect 12526 20924 12532 20936
rect 12439 20896 12532 20924
rect 12250 20816 12256 20868
rect 12308 20856 12314 20868
rect 12452 20865 12480 20896
rect 12526 20884 12532 20896
rect 12584 20924 12590 20936
rect 13173 20927 13231 20933
rect 13173 20924 13185 20927
rect 12584 20896 13185 20924
rect 12584 20884 12590 20896
rect 13173 20893 13185 20896
rect 13219 20924 13231 20927
rect 14108 20924 14136 20955
rect 14274 20952 14280 21004
rect 14332 20952 14338 21004
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20992 18843 20995
rect 19242 20992 19248 21004
rect 18831 20964 19248 20992
rect 18831 20961 18843 20964
rect 18785 20955 18843 20961
rect 19242 20952 19248 20964
rect 19300 20952 19306 21004
rect 22830 20992 22836 21004
rect 22743 20964 22836 20992
rect 22830 20952 22836 20964
rect 22888 20992 22894 21004
rect 23290 20992 23296 21004
rect 22888 20964 23296 20992
rect 22888 20952 22894 20964
rect 23290 20952 23296 20964
rect 23348 20952 23354 21004
rect 24118 20952 24124 21004
rect 24176 20992 24182 21004
rect 24176 20964 24716 20992
rect 24176 20952 24182 20964
rect 14642 20924 14648 20936
rect 13219 20896 13676 20924
rect 14108 20896 14648 20924
rect 13219 20893 13231 20896
rect 13173 20887 13231 20893
rect 12437 20859 12495 20865
rect 12437 20856 12449 20859
rect 12308 20828 12449 20856
rect 12308 20816 12314 20828
rect 12437 20825 12449 20828
rect 12483 20825 12495 20859
rect 12437 20819 12495 20825
rect 5031 20760 5764 20788
rect 5031 20757 5043 20760
rect 4985 20751 5043 20757
rect 6362 20748 6368 20800
rect 6420 20788 6426 20800
rect 8938 20788 8944 20800
rect 6420 20760 8944 20788
rect 6420 20748 6426 20760
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 11238 20788 11244 20800
rect 11112 20760 11244 20788
rect 11112 20748 11118 20760
rect 11238 20748 11244 20760
rect 11296 20748 11302 20800
rect 12618 20788 12624 20800
rect 12579 20760 12624 20788
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 13648 20797 13676 20896
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 15746 20884 15752 20936
rect 15804 20924 15810 20936
rect 15933 20927 15991 20933
rect 15933 20924 15945 20927
rect 15804 20896 15945 20924
rect 15804 20884 15810 20896
rect 15933 20893 15945 20896
rect 15979 20893 15991 20927
rect 19058 20924 19064 20936
rect 19019 20896 19064 20924
rect 15933 20887 15991 20893
rect 19058 20884 19064 20896
rect 19116 20884 19122 20936
rect 21082 20884 21088 20936
rect 21140 20924 21146 20936
rect 21361 20927 21419 20933
rect 21361 20924 21373 20927
rect 21140 20896 21373 20924
rect 21140 20884 21146 20896
rect 21361 20893 21373 20896
rect 21407 20893 21419 20927
rect 23106 20924 23112 20936
rect 23067 20896 23112 20924
rect 21361 20887 21419 20893
rect 23106 20884 23112 20896
rect 23164 20884 23170 20936
rect 24688 20933 24716 20964
rect 24581 20927 24639 20933
rect 24581 20893 24593 20927
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24673 20927 24731 20933
rect 24673 20893 24685 20927
rect 24719 20893 24731 20927
rect 25774 20924 25780 20936
rect 25735 20896 25780 20924
rect 24673 20887 24731 20893
rect 13906 20816 13912 20868
rect 13964 20856 13970 20868
rect 15381 20859 15439 20865
rect 15381 20856 15393 20859
rect 13964 20828 15393 20856
rect 13964 20816 13970 20828
rect 15381 20825 15393 20828
rect 15427 20825 15439 20859
rect 15381 20819 15439 20825
rect 16850 20816 16856 20868
rect 16908 20856 16914 20868
rect 16945 20859 17003 20865
rect 16945 20856 16957 20859
rect 16908 20828 16957 20856
rect 16908 20816 16914 20828
rect 16945 20825 16957 20828
rect 16991 20825 17003 20859
rect 16945 20819 17003 20825
rect 18141 20859 18199 20865
rect 18141 20825 18153 20859
rect 18187 20856 18199 20859
rect 18782 20856 18788 20868
rect 18187 20828 18788 20856
rect 18187 20825 18199 20828
rect 18141 20819 18199 20825
rect 18782 20816 18788 20828
rect 18840 20816 18846 20868
rect 20990 20856 20996 20868
rect 20951 20828 20996 20856
rect 20990 20816 20996 20828
rect 21048 20816 21054 20868
rect 22554 20856 22560 20868
rect 22515 20828 22560 20856
rect 22554 20816 22560 20828
rect 22612 20816 22618 20868
rect 23014 20816 23020 20868
rect 23072 20856 23078 20868
rect 24121 20859 24179 20865
rect 24121 20856 24133 20859
rect 23072 20828 24133 20856
rect 23072 20816 23078 20828
rect 24121 20825 24133 20828
rect 24167 20825 24179 20859
rect 24596 20856 24624 20887
rect 25774 20884 25780 20896
rect 25832 20884 25838 20936
rect 25038 20856 25044 20868
rect 24596 20828 25044 20856
rect 24121 20819 24179 20825
rect 25038 20816 25044 20828
rect 25096 20816 25102 20868
rect 25314 20816 25320 20868
rect 25372 20856 25378 20868
rect 25958 20856 25964 20868
rect 25372 20828 25964 20856
rect 25372 20816 25378 20828
rect 25958 20816 25964 20828
rect 26016 20816 26022 20868
rect 13633 20791 13691 20797
rect 13633 20757 13645 20791
rect 13679 20788 13691 20791
rect 13998 20788 14004 20800
rect 13679 20760 14004 20788
rect 13679 20757 13691 20760
rect 13633 20751 13691 20757
rect 13998 20748 14004 20760
rect 14056 20748 14062 20800
rect 18506 20788 18512 20800
rect 18467 20760 18512 20788
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 20346 20788 20352 20800
rect 20307 20760 20352 20788
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 22002 20788 22008 20800
rect 21963 20760 22008 20788
rect 22002 20748 22008 20760
rect 22060 20748 22066 20800
rect 22370 20788 22376 20800
rect 22331 20760 22376 20788
rect 22370 20748 22376 20760
rect 22428 20748 22434 20800
rect 22830 20748 22836 20800
rect 22888 20788 22894 20800
rect 23661 20791 23719 20797
rect 23661 20788 23673 20791
rect 22888 20760 23673 20788
rect 22888 20748 22894 20760
rect 23661 20757 23673 20760
rect 23707 20788 23719 20791
rect 24026 20788 24032 20800
rect 23707 20760 24032 20788
rect 23707 20757 23719 20760
rect 23661 20751 23719 20757
rect 24026 20748 24032 20760
rect 24084 20748 24090 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 2869 20587 2927 20593
rect 2869 20584 2881 20587
rect 2832 20556 2881 20584
rect 2832 20544 2838 20556
rect 2869 20553 2881 20556
rect 2915 20553 2927 20587
rect 2869 20547 2927 20553
rect 3050 20544 3056 20596
rect 3108 20584 3114 20596
rect 3421 20587 3479 20593
rect 3421 20584 3433 20587
rect 3108 20556 3433 20584
rect 3108 20544 3114 20556
rect 3421 20553 3433 20556
rect 3467 20553 3479 20587
rect 3421 20547 3479 20553
rect 3697 20587 3755 20593
rect 3697 20553 3709 20587
rect 3743 20584 3755 20587
rect 3878 20584 3884 20596
rect 3743 20556 3884 20584
rect 3743 20553 3755 20556
rect 3697 20547 3755 20553
rect 3878 20544 3884 20556
rect 3936 20544 3942 20596
rect 4154 20544 4160 20596
rect 4212 20584 4218 20596
rect 4709 20587 4767 20593
rect 4709 20584 4721 20587
rect 4212 20556 4721 20584
rect 4212 20544 4218 20556
rect 4709 20553 4721 20556
rect 4755 20584 4767 20587
rect 5442 20584 5448 20596
rect 4755 20556 5448 20584
rect 4755 20553 4767 20556
rect 4709 20547 4767 20553
rect 5442 20544 5448 20556
rect 5500 20544 5506 20596
rect 7561 20587 7619 20593
rect 7561 20553 7573 20587
rect 7607 20584 7619 20587
rect 7650 20584 7656 20596
rect 7607 20556 7656 20584
rect 7607 20553 7619 20556
rect 7561 20547 7619 20553
rect 7650 20544 7656 20556
rect 7708 20544 7714 20596
rect 9306 20584 9312 20596
rect 9267 20556 9312 20584
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 10873 20587 10931 20593
rect 10873 20553 10885 20587
rect 10919 20584 10931 20587
rect 10962 20584 10968 20596
rect 10919 20556 10968 20584
rect 10919 20553 10931 20556
rect 10873 20547 10931 20553
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 12066 20544 12072 20596
rect 12124 20584 12130 20596
rect 12253 20587 12311 20593
rect 12253 20584 12265 20587
rect 12124 20556 12265 20584
rect 12124 20544 12130 20556
rect 12253 20553 12265 20556
rect 12299 20584 12311 20587
rect 12434 20584 12440 20596
rect 12299 20556 12440 20584
rect 12299 20553 12311 20556
rect 12253 20547 12311 20553
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 14826 20584 14832 20596
rect 14787 20556 14832 20584
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15896 20556 15945 20584
rect 15896 20544 15902 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 16758 20584 16764 20596
rect 16719 20556 16764 20584
rect 15933 20547 15991 20553
rect 16758 20544 16764 20556
rect 16816 20544 16822 20596
rect 17037 20587 17095 20593
rect 17037 20553 17049 20587
rect 17083 20584 17095 20587
rect 17678 20584 17684 20596
rect 17083 20556 17684 20584
rect 17083 20553 17095 20556
rect 17037 20547 17095 20553
rect 17678 20544 17684 20556
rect 17736 20544 17742 20596
rect 17862 20544 17868 20596
rect 17920 20584 17926 20596
rect 17920 20556 17965 20584
rect 17920 20544 17926 20556
rect 18138 20544 18144 20596
rect 18196 20584 18202 20596
rect 18509 20587 18567 20593
rect 18509 20584 18521 20587
rect 18196 20556 18521 20584
rect 18196 20544 18202 20556
rect 18509 20553 18521 20556
rect 18555 20584 18567 20587
rect 19058 20584 19064 20596
rect 18555 20556 19064 20584
rect 18555 20553 18567 20556
rect 18509 20547 18567 20553
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19518 20544 19524 20596
rect 19576 20584 19582 20596
rect 20441 20587 20499 20593
rect 20441 20584 20453 20587
rect 19576 20556 20453 20584
rect 19576 20544 19582 20556
rect 20441 20553 20453 20556
rect 20487 20553 20499 20587
rect 20441 20547 20499 20553
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21542 20584 21548 20596
rect 20956 20556 21548 20584
rect 20956 20544 20962 20556
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 21818 20544 21824 20596
rect 21876 20584 21882 20596
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 21876 20556 22017 20584
rect 21876 20544 21882 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 22005 20547 22063 20553
rect 22094 20544 22100 20596
rect 22152 20584 22158 20596
rect 22152 20556 23428 20584
rect 22152 20544 22158 20556
rect 1762 20476 1768 20528
rect 1820 20516 1826 20528
rect 2133 20519 2191 20525
rect 2133 20516 2145 20519
rect 1820 20488 2145 20516
rect 1820 20476 1826 20488
rect 2133 20485 2145 20488
rect 2179 20516 2191 20519
rect 2590 20516 2596 20528
rect 2179 20488 2596 20516
rect 2179 20485 2191 20488
rect 2133 20479 2191 20485
rect 2590 20476 2596 20488
rect 2648 20476 2654 20528
rect 4062 20516 4068 20528
rect 3988 20488 4068 20516
rect 1946 20408 1952 20460
rect 2004 20448 2010 20460
rect 2685 20451 2743 20457
rect 2685 20448 2697 20451
rect 2004 20420 2697 20448
rect 2004 20408 2010 20420
rect 2685 20417 2697 20420
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 1118 20340 1124 20392
rect 1176 20380 1182 20392
rect 1176 20352 3188 20380
rect 1176 20340 1182 20352
rect 1854 20272 1860 20324
rect 1912 20312 1918 20324
rect 1949 20315 2007 20321
rect 1949 20312 1961 20315
rect 1912 20284 1961 20312
rect 1912 20272 1918 20284
rect 1949 20281 1961 20284
rect 1995 20312 2007 20315
rect 2409 20315 2467 20321
rect 2409 20312 2421 20315
rect 1995 20284 2421 20312
rect 1995 20281 2007 20284
rect 1949 20275 2007 20281
rect 2409 20281 2421 20284
rect 2455 20281 2467 20315
rect 3160 20312 3188 20352
rect 3234 20340 3240 20392
rect 3292 20380 3298 20392
rect 3988 20389 4016 20488
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 5261 20519 5319 20525
rect 5261 20485 5273 20519
rect 5307 20516 5319 20519
rect 5350 20516 5356 20528
rect 5307 20488 5356 20516
rect 5307 20485 5319 20488
rect 5261 20479 5319 20485
rect 5350 20476 5356 20488
rect 5408 20476 5414 20528
rect 4246 20448 4252 20460
rect 4207 20420 4252 20448
rect 4246 20408 4252 20420
rect 4304 20408 4310 20460
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20448 5871 20451
rect 5994 20448 6000 20460
rect 5859 20420 6000 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 5994 20408 6000 20420
rect 6052 20448 6058 20460
rect 6454 20448 6460 20460
rect 6052 20420 6460 20448
rect 6052 20408 6058 20420
rect 6454 20408 6460 20420
rect 6512 20408 6518 20460
rect 7668 20448 7696 20544
rect 9674 20476 9680 20528
rect 9732 20516 9738 20528
rect 10321 20519 10379 20525
rect 10321 20516 10333 20519
rect 9732 20488 10333 20516
rect 9732 20476 9738 20488
rect 10321 20485 10333 20488
rect 10367 20516 10379 20519
rect 12342 20516 12348 20528
rect 10367 20488 12348 20516
rect 10367 20485 10379 20488
rect 10321 20479 10379 20485
rect 12342 20476 12348 20488
rect 12400 20476 12406 20528
rect 13814 20476 13820 20528
rect 13872 20516 13878 20528
rect 15013 20519 15071 20525
rect 15013 20516 15025 20519
rect 13872 20488 15025 20516
rect 13872 20476 13878 20488
rect 15013 20485 15025 20488
rect 15059 20485 15071 20519
rect 16850 20516 16856 20528
rect 15013 20479 15071 20485
rect 15212 20488 16856 20516
rect 8113 20451 8171 20457
rect 8113 20448 8125 20451
rect 7668 20420 8125 20448
rect 8113 20417 8125 20420
rect 8159 20417 8171 20451
rect 8113 20411 8171 20417
rect 8297 20451 8355 20457
rect 8297 20417 8309 20451
rect 8343 20448 8355 20451
rect 8386 20448 8392 20460
rect 8343 20420 8392 20448
rect 8343 20417 8355 20420
rect 8297 20411 8355 20417
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 9769 20451 9827 20457
rect 9769 20417 9781 20451
rect 9815 20448 9827 20451
rect 9950 20448 9956 20460
rect 9815 20420 9956 20448
rect 9815 20417 9827 20420
rect 9769 20411 9827 20417
rect 9950 20408 9956 20420
rect 10008 20408 10014 20460
rect 10778 20448 10784 20460
rect 10612 20420 10784 20448
rect 3973 20383 4031 20389
rect 3973 20380 3985 20383
rect 3292 20352 3985 20380
rect 3292 20340 3298 20352
rect 3973 20349 3985 20352
rect 4019 20349 4031 20383
rect 3973 20343 4031 20349
rect 5258 20340 5264 20392
rect 5316 20380 5322 20392
rect 5537 20383 5595 20389
rect 5537 20380 5549 20383
rect 5316 20352 5549 20380
rect 5316 20340 5322 20352
rect 5537 20349 5549 20352
rect 5583 20380 5595 20383
rect 7727 20383 7785 20389
rect 7727 20380 7739 20383
rect 5583 20352 7739 20380
rect 5583 20349 5595 20352
rect 5537 20343 5595 20349
rect 7727 20349 7739 20352
rect 7773 20349 7785 20383
rect 7727 20343 7785 20349
rect 9125 20383 9183 20389
rect 9125 20349 9137 20383
rect 9171 20380 9183 20383
rect 9861 20383 9919 20389
rect 9861 20380 9873 20383
rect 9171 20352 9873 20380
rect 9171 20349 9183 20352
rect 9125 20343 9183 20349
rect 9861 20349 9873 20352
rect 9907 20380 9919 20383
rect 10612 20380 10640 20420
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 11330 20448 11336 20460
rect 11291 20420 11336 20448
rect 11330 20408 11336 20420
rect 11388 20408 11394 20460
rect 11808 20420 12572 20448
rect 11808 20389 11836 20420
rect 12544 20392 12572 20420
rect 14734 20408 14740 20460
rect 14792 20448 14798 20460
rect 15212 20448 15240 20488
rect 16850 20476 16856 20488
rect 16908 20516 16914 20528
rect 17405 20519 17463 20525
rect 17405 20516 17417 20519
rect 16908 20488 17417 20516
rect 16908 20476 16914 20488
rect 17405 20485 17417 20488
rect 17451 20516 17463 20519
rect 18598 20516 18604 20528
rect 17451 20488 18604 20516
rect 17451 20485 17463 20488
rect 17405 20479 17463 20485
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 18874 20516 18880 20528
rect 18835 20488 18880 20516
rect 18874 20476 18880 20488
rect 18932 20476 18938 20528
rect 21729 20519 21787 20525
rect 21729 20485 21741 20519
rect 21775 20516 21787 20519
rect 22462 20516 22468 20528
rect 21775 20488 22468 20516
rect 21775 20485 21787 20488
rect 21729 20479 21787 20485
rect 22462 20476 22468 20488
rect 22520 20516 22526 20528
rect 22520 20488 22692 20516
rect 22520 20476 22526 20488
rect 15378 20448 15384 20460
rect 14792 20420 15240 20448
rect 15339 20420 15384 20448
rect 14792 20408 14798 20420
rect 15378 20408 15384 20420
rect 15436 20408 15442 20460
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 16206 20448 16212 20460
rect 15620 20420 16212 20448
rect 15620 20408 15626 20420
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 19242 20448 19248 20460
rect 19203 20420 19248 20448
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 20070 20408 20076 20460
rect 20128 20448 20134 20460
rect 20257 20451 20315 20457
rect 20257 20448 20269 20451
rect 20128 20420 20269 20448
rect 20128 20408 20134 20420
rect 20257 20417 20269 20420
rect 20303 20448 20315 20451
rect 20898 20448 20904 20460
rect 20303 20420 20904 20448
rect 20303 20417 20315 20420
rect 20257 20411 20315 20417
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 22370 20408 22376 20460
rect 22428 20448 22434 20460
rect 22557 20451 22615 20457
rect 22557 20448 22569 20451
rect 22428 20420 22569 20448
rect 22428 20408 22434 20420
rect 22557 20417 22569 20420
rect 22603 20417 22615 20451
rect 22557 20411 22615 20417
rect 9907 20352 10640 20380
rect 10689 20383 10747 20389
rect 9907 20349 9919 20352
rect 9861 20343 9919 20349
rect 10689 20349 10701 20383
rect 10735 20380 10747 20383
rect 11425 20383 11483 20389
rect 11425 20380 11437 20383
rect 10735 20352 11437 20380
rect 10735 20349 10747 20352
rect 10689 20343 10747 20349
rect 11425 20349 11437 20352
rect 11471 20380 11483 20383
rect 11793 20383 11851 20389
rect 11793 20380 11805 20383
rect 11471 20352 11805 20380
rect 11471 20349 11483 20352
rect 11425 20343 11483 20349
rect 11793 20349 11805 20352
rect 11839 20349 11851 20383
rect 12434 20380 12440 20392
rect 12395 20352 12440 20380
rect 11793 20343 11851 20349
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 12526 20340 12532 20392
rect 12584 20380 12590 20392
rect 12693 20383 12751 20389
rect 12693 20380 12705 20383
rect 12584 20352 12705 20380
rect 12584 20340 12590 20352
rect 12693 20349 12705 20352
rect 12739 20349 12751 20383
rect 12693 20343 12751 20349
rect 16850 20340 16856 20392
rect 16908 20389 16914 20392
rect 16908 20380 16917 20389
rect 16908 20352 16953 20380
rect 16908 20343 16917 20352
rect 16908 20340 16914 20343
rect 20346 20340 20352 20392
rect 20404 20380 20410 20392
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20404 20352 21005 20380
rect 20404 20340 20410 20352
rect 20993 20349 21005 20352
rect 21039 20349 21051 20383
rect 22664 20380 22692 20488
rect 23400 20392 23428 20556
rect 23474 20544 23480 20596
rect 23532 20584 23538 20596
rect 23753 20587 23811 20593
rect 23753 20584 23765 20587
rect 23532 20556 23765 20584
rect 23532 20544 23538 20556
rect 23753 20553 23765 20556
rect 23799 20553 23811 20587
rect 23753 20547 23811 20553
rect 20993 20343 21051 20349
rect 22480 20352 22692 20380
rect 5350 20312 5356 20324
rect 3160 20284 5356 20312
rect 2409 20275 2467 20281
rect 5350 20272 5356 20284
rect 5408 20272 5414 20324
rect 5902 20272 5908 20324
rect 5960 20312 5966 20324
rect 6549 20315 6607 20321
rect 6549 20312 6561 20315
rect 5960 20284 6561 20312
rect 5960 20272 5966 20284
rect 6549 20281 6561 20284
rect 6595 20312 6607 20315
rect 6638 20312 6644 20324
rect 6595 20284 6644 20312
rect 6595 20281 6607 20284
rect 6549 20275 6607 20281
rect 6638 20272 6644 20284
rect 6696 20272 6702 20324
rect 9766 20312 9772 20324
rect 9727 20284 9772 20312
rect 9766 20272 9772 20284
rect 9824 20272 9830 20324
rect 11238 20272 11244 20324
rect 11296 20312 11302 20324
rect 11333 20315 11391 20321
rect 11333 20312 11345 20315
rect 11296 20284 11345 20312
rect 11296 20272 11302 20284
rect 11333 20281 11345 20284
rect 11379 20281 11391 20315
rect 15470 20312 15476 20324
rect 15431 20284 15476 20312
rect 11333 20275 11391 20281
rect 15470 20272 15476 20284
rect 15528 20272 15534 20324
rect 15565 20315 15623 20321
rect 15565 20281 15577 20315
rect 15611 20281 15623 20315
rect 19426 20312 19432 20324
rect 19387 20284 19432 20312
rect 15565 20275 15623 20281
rect 1302 20204 1308 20256
rect 1360 20244 1366 20256
rect 1578 20244 1584 20256
rect 1360 20216 1584 20244
rect 1360 20204 1366 20216
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 2130 20204 2136 20256
rect 2188 20244 2194 20256
rect 2593 20247 2651 20253
rect 2593 20244 2605 20247
rect 2188 20216 2605 20244
rect 2188 20204 2194 20216
rect 2593 20213 2605 20216
rect 2639 20213 2651 20247
rect 2593 20207 2651 20213
rect 2869 20247 2927 20253
rect 2869 20213 2881 20247
rect 2915 20244 2927 20247
rect 3145 20247 3203 20253
rect 3145 20244 3157 20247
rect 2915 20216 3157 20244
rect 2915 20213 2927 20216
rect 2869 20207 2927 20213
rect 3145 20213 3157 20216
rect 3191 20244 3203 20247
rect 3234 20244 3240 20256
rect 3191 20216 3240 20244
rect 3191 20213 3203 20216
rect 3145 20207 3203 20213
rect 3234 20204 3240 20216
rect 3292 20204 3298 20256
rect 3970 20204 3976 20256
rect 4028 20244 4034 20256
rect 4157 20247 4215 20253
rect 4157 20244 4169 20247
rect 4028 20216 4169 20244
rect 4028 20204 4034 20216
rect 4157 20213 4169 20216
rect 4203 20213 4215 20247
rect 4157 20207 4215 20213
rect 4246 20204 4252 20256
rect 4304 20244 4310 20256
rect 4982 20244 4988 20256
rect 4304 20216 4988 20244
rect 4304 20204 4310 20216
rect 4982 20204 4988 20216
rect 5040 20204 5046 20256
rect 5721 20247 5779 20253
rect 5721 20213 5733 20247
rect 5767 20244 5779 20247
rect 6178 20244 6184 20256
rect 5767 20216 6184 20244
rect 5767 20213 5779 20216
rect 5721 20207 5779 20213
rect 6178 20204 6184 20216
rect 6236 20204 6242 20256
rect 6273 20247 6331 20253
rect 6273 20213 6285 20247
rect 6319 20244 6331 20247
rect 6454 20244 6460 20256
rect 6319 20216 6460 20244
rect 6319 20213 6331 20216
rect 6273 20207 6331 20213
rect 6454 20204 6460 20216
rect 6512 20204 6518 20256
rect 7193 20247 7251 20253
rect 7193 20213 7205 20247
rect 7239 20244 7251 20247
rect 8018 20244 8024 20256
rect 7239 20216 8024 20244
rect 7239 20213 7251 20216
rect 7193 20207 7251 20213
rect 8018 20204 8024 20216
rect 8076 20244 8082 20256
rect 8205 20247 8263 20253
rect 8205 20244 8217 20247
rect 8076 20216 8217 20244
rect 8076 20204 8082 20216
rect 8205 20213 8217 20216
rect 8251 20213 8263 20247
rect 8205 20207 8263 20213
rect 8386 20204 8392 20256
rect 8444 20244 8450 20256
rect 8665 20247 8723 20253
rect 8665 20244 8677 20247
rect 8444 20216 8677 20244
rect 8444 20204 8450 20216
rect 8665 20213 8677 20216
rect 8711 20213 8723 20247
rect 8665 20207 8723 20213
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 12342 20244 12348 20256
rect 9732 20216 12348 20244
rect 9732 20204 9738 20216
rect 12342 20204 12348 20216
rect 12400 20204 12406 20256
rect 13446 20204 13452 20256
rect 13504 20244 13510 20256
rect 13817 20247 13875 20253
rect 13817 20244 13829 20247
rect 13504 20216 13829 20244
rect 13504 20204 13510 20216
rect 13817 20213 13829 20216
rect 13863 20213 13875 20247
rect 14366 20244 14372 20256
rect 14327 20216 14372 20244
rect 13817 20207 13875 20213
rect 14366 20204 14372 20216
rect 14424 20244 14430 20256
rect 15580 20244 15608 20275
rect 19426 20272 19432 20284
rect 19484 20272 19490 20324
rect 22094 20272 22100 20324
rect 22152 20312 22158 20324
rect 22480 20321 22508 20352
rect 22281 20315 22339 20321
rect 22281 20312 22293 20315
rect 22152 20284 22293 20312
rect 22152 20272 22158 20284
rect 22281 20281 22293 20284
rect 22327 20281 22339 20315
rect 22281 20275 22339 20281
rect 22465 20315 22523 20321
rect 22465 20281 22477 20315
rect 22511 20281 22523 20315
rect 22465 20275 22523 20281
rect 22572 20256 22600 20352
rect 23382 20340 23388 20392
rect 23440 20340 23446 20392
rect 25222 20380 25228 20392
rect 23860 20352 24164 20380
rect 25183 20352 25228 20380
rect 23109 20315 23167 20321
rect 23109 20281 23121 20315
rect 23155 20312 23167 20315
rect 23860 20312 23888 20352
rect 24136 20324 24164 20352
rect 25222 20340 25228 20352
rect 25280 20380 25286 20392
rect 25961 20383 26019 20389
rect 25961 20380 25973 20383
rect 25280 20352 25973 20380
rect 25280 20340 25286 20352
rect 25961 20349 25973 20352
rect 26007 20349 26019 20383
rect 25961 20343 26019 20349
rect 24026 20312 24032 20324
rect 23155 20284 23888 20312
rect 23987 20284 24032 20312
rect 23155 20281 23167 20284
rect 23109 20275 23167 20281
rect 24026 20272 24032 20284
rect 24084 20272 24090 20324
rect 24118 20272 24124 20324
rect 24176 20312 24182 20324
rect 24302 20312 24308 20324
rect 24176 20284 24308 20312
rect 24176 20272 24182 20284
rect 24302 20272 24308 20284
rect 24360 20272 24366 20324
rect 25501 20315 25559 20321
rect 25501 20281 25513 20315
rect 25547 20312 25559 20315
rect 25774 20312 25780 20324
rect 25547 20284 25780 20312
rect 25547 20281 25559 20284
rect 25501 20275 25559 20281
rect 25774 20272 25780 20284
rect 25832 20272 25838 20324
rect 15746 20244 15752 20256
rect 14424 20216 15752 20244
rect 14424 20204 14430 20216
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 16393 20247 16451 20253
rect 16393 20213 16405 20247
rect 16439 20244 16451 20247
rect 16666 20244 16672 20256
rect 16439 20216 16672 20244
rect 16439 20213 16451 20216
rect 16393 20207 16451 20213
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 19334 20244 19340 20256
rect 19295 20216 19340 20244
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19797 20247 19855 20253
rect 19797 20244 19809 20247
rect 19576 20216 19809 20244
rect 19576 20204 19582 20216
rect 19797 20213 19809 20216
rect 19843 20213 19855 20247
rect 20898 20244 20904 20256
rect 20859 20216 20904 20244
rect 19797 20207 19855 20213
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 21358 20244 21364 20256
rect 21319 20216 21364 20244
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 22554 20204 22560 20256
rect 22612 20204 22618 20256
rect 23474 20244 23480 20256
rect 23435 20216 23480 20244
rect 23474 20204 23480 20216
rect 23532 20244 23538 20256
rect 24213 20247 24271 20253
rect 24213 20244 24225 20247
rect 23532 20216 24225 20244
rect 23532 20204 23538 20216
rect 24213 20213 24225 20216
rect 24259 20213 24271 20247
rect 24670 20244 24676 20256
rect 24631 20216 24676 20244
rect 24213 20207 24271 20213
rect 24670 20204 24676 20216
rect 24728 20204 24734 20256
rect 25038 20244 25044 20256
rect 24999 20216 25044 20244
rect 25038 20204 25044 20216
rect 25096 20204 25102 20256
rect 26326 20244 26332 20256
rect 26287 20216 26332 20244
rect 26326 20204 26332 20216
rect 26384 20204 26390 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1765 20043 1823 20049
rect 1765 20009 1777 20043
rect 1811 20040 1823 20043
rect 1946 20040 1952 20052
rect 1811 20012 1952 20040
rect 1811 20009 1823 20012
rect 1765 20003 1823 20009
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 2130 20040 2136 20052
rect 2091 20012 2136 20040
rect 2130 20000 2136 20012
rect 2188 20000 2194 20052
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 2961 20043 3019 20049
rect 2961 20040 2973 20043
rect 2924 20012 2973 20040
rect 2924 20000 2930 20012
rect 2961 20009 2973 20012
rect 3007 20040 3019 20043
rect 3510 20040 3516 20052
rect 3007 20012 3516 20040
rect 3007 20009 3019 20012
rect 2961 20003 3019 20009
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 3786 20000 3792 20052
rect 3844 20040 3850 20052
rect 4893 20043 4951 20049
rect 4893 20040 4905 20043
rect 3844 20012 4905 20040
rect 3844 20000 3850 20012
rect 4893 20009 4905 20012
rect 4939 20040 4951 20043
rect 5258 20040 5264 20052
rect 4939 20012 5264 20040
rect 4939 20009 4951 20012
rect 4893 20003 4951 20009
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 7282 20040 7288 20052
rect 7243 20012 7288 20040
rect 7282 20000 7288 20012
rect 7340 20000 7346 20052
rect 7929 20043 7987 20049
rect 7929 20009 7941 20043
rect 7975 20040 7987 20043
rect 8294 20040 8300 20052
rect 7975 20012 8300 20040
rect 7975 20009 7987 20012
rect 7929 20003 7987 20009
rect 4709 19975 4767 19981
rect 4709 19941 4721 19975
rect 4755 19972 4767 19975
rect 5166 19972 5172 19984
rect 4755 19944 5172 19972
rect 4755 19941 4767 19944
rect 4709 19935 4767 19941
rect 5166 19932 5172 19944
rect 5224 19932 5230 19984
rect 5813 19975 5871 19981
rect 5813 19941 5825 19975
rect 5859 19972 5871 19975
rect 6086 19972 6092 19984
rect 5859 19944 6092 19972
rect 5859 19941 5871 19944
rect 5813 19935 5871 19941
rect 6086 19932 6092 19944
rect 6144 19972 6150 19984
rect 7944 19972 7972 20003
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 9493 20043 9551 20049
rect 9493 20009 9505 20043
rect 9539 20040 9551 20043
rect 9582 20040 9588 20052
rect 9539 20012 9588 20040
rect 9539 20009 9551 20012
rect 9493 20003 9551 20009
rect 9582 20000 9588 20012
rect 9640 20000 9646 20052
rect 12894 20000 12900 20052
rect 12952 20040 12958 20052
rect 13446 20040 13452 20052
rect 12952 20012 13452 20040
rect 12952 20000 12958 20012
rect 13446 20000 13452 20012
rect 13504 20040 13510 20052
rect 13633 20043 13691 20049
rect 13633 20040 13645 20043
rect 13504 20012 13645 20040
rect 13504 20000 13510 20012
rect 13633 20009 13645 20012
rect 13679 20009 13691 20043
rect 13633 20003 13691 20009
rect 14185 20043 14243 20049
rect 14185 20009 14197 20043
rect 14231 20040 14243 20043
rect 14366 20040 14372 20052
rect 14231 20012 14372 20040
rect 14231 20009 14243 20012
rect 14185 20003 14243 20009
rect 14366 20000 14372 20012
rect 14424 20000 14430 20052
rect 14642 20040 14648 20052
rect 14603 20012 14648 20040
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 15013 20043 15071 20049
rect 15013 20009 15025 20043
rect 15059 20040 15071 20043
rect 15470 20040 15476 20052
rect 15059 20012 15476 20040
rect 15059 20009 15071 20012
rect 15013 20003 15071 20009
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 15746 20040 15752 20052
rect 15707 20012 15752 20040
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 16942 20000 16948 20052
rect 17000 20040 17006 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 17000 20012 17693 20040
rect 17000 20000 17006 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 17681 20003 17739 20009
rect 18877 20043 18935 20049
rect 18877 20009 18889 20043
rect 18923 20040 18935 20043
rect 19426 20040 19432 20052
rect 18923 20012 19432 20040
rect 18923 20009 18935 20012
rect 18877 20003 18935 20009
rect 19426 20000 19432 20012
rect 19484 20000 19490 20052
rect 19521 20043 19579 20049
rect 19521 20009 19533 20043
rect 19567 20040 19579 20043
rect 19889 20043 19947 20049
rect 19889 20040 19901 20043
rect 19567 20012 19901 20040
rect 19567 20009 19579 20012
rect 19521 20003 19579 20009
rect 19889 20009 19901 20012
rect 19935 20009 19947 20043
rect 19889 20003 19947 20009
rect 24118 20000 24124 20052
rect 24176 20040 24182 20052
rect 25409 20043 25467 20049
rect 25409 20040 25421 20043
rect 24176 20012 25421 20040
rect 24176 20000 24182 20012
rect 25409 20009 25421 20012
rect 25455 20009 25467 20043
rect 25409 20003 25467 20009
rect 6144 19944 7972 19972
rect 6144 19932 6150 19944
rect 9674 19932 9680 19984
rect 9732 19972 9738 19984
rect 10229 19975 10287 19981
rect 10229 19972 10241 19975
rect 9732 19944 10241 19972
rect 9732 19932 9738 19944
rect 10229 19941 10241 19944
rect 10275 19941 10287 19975
rect 10229 19935 10287 19941
rect 11330 19932 11336 19984
rect 11388 19972 11394 19984
rect 12069 19975 12127 19981
rect 12069 19972 12081 19975
rect 11388 19944 12081 19972
rect 11388 19932 11394 19944
rect 12069 19941 12081 19944
rect 12115 19941 12127 19975
rect 12069 19935 12127 19941
rect 12342 19932 12348 19984
rect 12400 19972 12406 19984
rect 15286 19972 15292 19984
rect 12400 19944 13860 19972
rect 15247 19944 15292 19972
rect 12400 19932 12406 19944
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 3697 19907 3755 19913
rect 2832 19876 2877 19904
rect 2832 19864 2838 19876
rect 3697 19873 3709 19907
rect 3743 19904 3755 19907
rect 5445 19907 5503 19913
rect 3743 19876 5028 19904
rect 3743 19873 3755 19876
rect 3697 19867 3755 19873
rect 5000 19848 5028 19876
rect 5445 19873 5457 19907
rect 5491 19904 5503 19907
rect 5534 19904 5540 19916
rect 5491 19876 5540 19904
rect 5491 19873 5503 19876
rect 5445 19867 5503 19873
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 5902 19904 5908 19916
rect 5863 19876 5908 19904
rect 5902 19864 5908 19876
rect 5960 19864 5966 19916
rect 6172 19907 6230 19913
rect 6172 19904 6184 19907
rect 6012 19876 6184 19904
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19836 3111 19839
rect 3234 19836 3240 19848
rect 3099 19808 3240 19836
rect 3099 19805 3111 19808
rect 3053 19799 3111 19805
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 4982 19836 4988 19848
rect 4895 19808 4988 19836
rect 4982 19796 4988 19808
rect 5040 19836 5046 19848
rect 6012 19836 6040 19876
rect 6172 19873 6184 19876
rect 6218 19904 6230 19907
rect 6454 19904 6460 19916
rect 6218 19876 6460 19904
rect 6218 19873 6230 19876
rect 6172 19867 6230 19873
rect 6454 19864 6460 19876
rect 6512 19904 6518 19916
rect 6638 19904 6644 19916
rect 6512 19876 6644 19904
rect 6512 19864 6518 19876
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19904 9183 19907
rect 10045 19907 10103 19913
rect 10045 19904 10057 19907
rect 9171 19876 10057 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 10045 19873 10057 19876
rect 10091 19904 10103 19907
rect 10594 19904 10600 19916
rect 10091 19876 10600 19904
rect 10091 19873 10103 19876
rect 10045 19867 10103 19873
rect 10594 19864 10600 19876
rect 10652 19864 10658 19916
rect 11425 19907 11483 19913
rect 11425 19873 11437 19907
rect 11471 19904 11483 19907
rect 12161 19907 12219 19913
rect 12161 19904 12173 19907
rect 11471 19876 12173 19904
rect 11471 19873 11483 19876
rect 11425 19867 11483 19873
rect 12161 19873 12173 19876
rect 12207 19904 12219 19907
rect 12894 19904 12900 19916
rect 12207 19876 12900 19904
rect 12207 19873 12219 19876
rect 12161 19867 12219 19873
rect 12894 19864 12900 19876
rect 12952 19904 12958 19916
rect 12989 19907 13047 19913
rect 12989 19904 13001 19907
rect 12952 19876 13001 19904
rect 12952 19864 12958 19876
rect 12989 19873 13001 19876
rect 13035 19904 13047 19907
rect 13725 19907 13783 19913
rect 13725 19904 13737 19907
rect 13035 19876 13737 19904
rect 13035 19873 13047 19876
rect 12989 19867 13047 19873
rect 13725 19873 13737 19876
rect 13771 19873 13783 19907
rect 13832 19904 13860 19944
rect 15286 19932 15292 19944
rect 15344 19932 15350 19984
rect 16482 19932 16488 19984
rect 16540 19981 16546 19984
rect 16540 19975 16604 19981
rect 16540 19941 16558 19975
rect 16592 19941 16604 19975
rect 16540 19935 16604 19941
rect 19613 19975 19671 19981
rect 19613 19941 19625 19975
rect 19659 19972 19671 19975
rect 19978 19972 19984 19984
rect 19659 19944 19984 19972
rect 19659 19941 19671 19944
rect 19613 19935 19671 19941
rect 16540 19932 16546 19935
rect 19978 19932 19984 19944
rect 20036 19932 20042 19984
rect 20073 19975 20131 19981
rect 20073 19941 20085 19975
rect 20119 19972 20131 19975
rect 21450 19972 21456 19984
rect 20119 19944 21456 19972
rect 20119 19941 20131 19944
rect 20073 19935 20131 19941
rect 21450 19932 21456 19944
rect 21508 19932 21514 19984
rect 21542 19932 21548 19984
rect 21600 19932 21606 19984
rect 23106 19972 23112 19984
rect 22480 19944 23112 19972
rect 16390 19904 16396 19916
rect 13832 19876 16396 19904
rect 13725 19867 13783 19873
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 19150 19864 19156 19916
rect 19208 19904 19214 19916
rect 20441 19907 20499 19913
rect 20441 19904 20453 19907
rect 19208 19876 20453 19904
rect 19208 19864 19214 19876
rect 20441 19873 20453 19876
rect 20487 19904 20499 19907
rect 20898 19904 20904 19916
rect 20487 19876 20904 19904
rect 20487 19873 20499 19876
rect 20441 19867 20499 19873
rect 20898 19864 20904 19876
rect 20956 19864 20962 19916
rect 21358 19904 21364 19916
rect 21271 19876 21364 19904
rect 21358 19864 21364 19876
rect 21416 19904 21422 19916
rect 21560 19904 21588 19932
rect 21416 19876 21588 19904
rect 21628 19907 21686 19913
rect 21416 19864 21422 19876
rect 21628 19873 21640 19907
rect 21674 19904 21686 19907
rect 22094 19904 22100 19916
rect 21674 19876 22100 19904
rect 21674 19873 21686 19876
rect 21628 19867 21686 19873
rect 22094 19864 22100 19876
rect 22152 19904 22158 19916
rect 22480 19904 22508 19944
rect 23106 19932 23112 19944
rect 23164 19972 23170 19984
rect 23385 19975 23443 19981
rect 23385 19972 23397 19975
rect 23164 19944 23397 19972
rect 23164 19932 23170 19944
rect 23385 19941 23397 19944
rect 23431 19941 23443 19975
rect 23385 19935 23443 19941
rect 23566 19932 23572 19984
rect 23624 19972 23630 19984
rect 24397 19975 24455 19981
rect 24397 19972 24409 19975
rect 23624 19944 24409 19972
rect 23624 19932 23630 19944
rect 24397 19941 24409 19944
rect 24443 19941 24455 19975
rect 24397 19935 24455 19941
rect 22152 19876 22508 19904
rect 22152 19864 22158 19876
rect 22830 19864 22836 19916
rect 22888 19864 22894 19916
rect 23290 19864 23296 19916
rect 23348 19904 23354 19916
rect 25869 19907 25927 19913
rect 25869 19904 25881 19907
rect 23348 19876 25881 19904
rect 23348 19864 23354 19876
rect 25869 19873 25881 19876
rect 25915 19873 25927 19907
rect 25869 19867 25927 19873
rect 5040 19808 6040 19836
rect 8573 19839 8631 19845
rect 5040 19796 5046 19808
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 9858 19836 9864 19848
rect 8619 19808 9864 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 10321 19839 10379 19845
rect 10321 19805 10333 19839
rect 10367 19836 10379 19839
rect 10778 19836 10784 19848
rect 10367 19808 10784 19836
rect 10367 19805 10379 19808
rect 10321 19799 10379 19805
rect 10778 19796 10784 19808
rect 10836 19796 10842 19848
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 11977 19839 12035 19845
rect 11977 19836 11989 19839
rect 11664 19808 11989 19836
rect 11664 19796 11670 19808
rect 11977 19805 11989 19808
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 12342 19796 12348 19848
rect 12400 19796 12406 19848
rect 13630 19836 13636 19848
rect 13591 19808 13636 19836
rect 13630 19796 13636 19808
rect 13688 19796 13694 19848
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16301 19839 16359 19845
rect 16301 19836 16313 19839
rect 15988 19808 16313 19836
rect 15988 19796 15994 19808
rect 16301 19805 16313 19808
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 17862 19796 17868 19848
rect 17920 19836 17926 19848
rect 18322 19836 18328 19848
rect 17920 19808 18328 19836
rect 17920 19796 17926 19808
rect 18322 19796 18328 19808
rect 18380 19836 18386 19848
rect 19521 19839 19579 19845
rect 18380 19808 19380 19836
rect 18380 19796 18386 19808
rect 2498 19768 2504 19780
rect 2459 19740 2504 19768
rect 2498 19728 2504 19740
rect 2556 19728 2562 19780
rect 4433 19771 4491 19777
rect 4433 19737 4445 19771
rect 4479 19768 4491 19771
rect 5442 19768 5448 19780
rect 4479 19740 5448 19768
rect 4479 19737 4491 19740
rect 4433 19731 4491 19737
rect 5442 19728 5448 19740
rect 5500 19728 5506 19780
rect 10870 19728 10876 19780
rect 10928 19768 10934 19780
rect 11698 19768 11704 19780
rect 10928 19740 11704 19768
rect 10928 19728 10934 19740
rect 11698 19728 11704 19740
rect 11756 19768 11762 19780
rect 12360 19768 12388 19796
rect 11756 19740 12388 19768
rect 11756 19728 11762 19740
rect 12434 19728 12440 19780
rect 12492 19768 12498 19780
rect 12621 19771 12679 19777
rect 12621 19768 12633 19771
rect 12492 19740 12633 19768
rect 12492 19728 12498 19740
rect 12621 19737 12633 19740
rect 12667 19768 12679 19771
rect 13722 19768 13728 19780
rect 12667 19740 13728 19768
rect 12667 19737 12679 19740
rect 12621 19731 12679 19737
rect 13722 19728 13728 19740
rect 13780 19728 13786 19780
rect 19061 19771 19119 19777
rect 19061 19737 19073 19771
rect 19107 19768 19119 19771
rect 19242 19768 19248 19780
rect 19107 19740 19248 19768
rect 19107 19737 19119 19740
rect 19061 19731 19119 19737
rect 19242 19728 19248 19740
rect 19300 19728 19306 19780
rect 19352 19768 19380 19808
rect 19521 19805 19533 19839
rect 19567 19836 19579 19839
rect 20346 19836 20352 19848
rect 19567 19808 20352 19836
rect 19567 19805 19579 19808
rect 19521 19799 19579 19805
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 22848 19768 22876 19864
rect 23474 19796 23480 19848
rect 23532 19836 23538 19848
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 23532 19808 23673 19836
rect 23532 19796 23538 19808
rect 23661 19805 23673 19808
rect 23707 19836 23719 19839
rect 24026 19836 24032 19848
rect 23707 19808 24032 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19805 24455 19839
rect 24397 19799 24455 19805
rect 24489 19839 24547 19845
rect 24489 19805 24501 19839
rect 24535 19836 24547 19839
rect 24762 19836 24768 19848
rect 24535 19808 24768 19836
rect 24535 19805 24547 19808
rect 24489 19799 24547 19805
rect 23290 19768 23296 19780
rect 19352 19740 21220 19768
rect 22848 19740 23296 19768
rect 3878 19660 3884 19712
rect 3936 19700 3942 19712
rect 7834 19700 7840 19712
rect 3936 19672 7840 19700
rect 3936 19660 3942 19672
rect 7834 19660 7840 19672
rect 7892 19660 7898 19712
rect 9766 19700 9772 19712
rect 9727 19672 9772 19700
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 10781 19703 10839 19709
rect 10781 19669 10793 19703
rect 10827 19700 10839 19703
rect 10962 19700 10968 19712
rect 10827 19672 10968 19700
rect 10827 19669 10839 19672
rect 10781 19663 10839 19669
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 11609 19703 11667 19709
rect 11609 19669 11621 19703
rect 11655 19700 11667 19703
rect 12250 19700 12256 19712
rect 11655 19672 12256 19700
rect 11655 19669 11667 19672
rect 11609 19663 11667 19669
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 13170 19700 13176 19712
rect 13131 19672 13176 19700
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 16114 19700 16120 19712
rect 16075 19672 16120 19700
rect 16114 19660 16120 19672
rect 16172 19660 16178 19712
rect 18322 19700 18328 19712
rect 18283 19672 18328 19700
rect 18322 19660 18328 19672
rect 18380 19660 18386 19712
rect 19889 19703 19947 19709
rect 19889 19669 19901 19703
rect 19935 19700 19947 19703
rect 20070 19700 20076 19712
rect 19935 19672 20076 19700
rect 19935 19669 19947 19672
rect 19889 19663 19947 19669
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20898 19660 20904 19712
rect 20956 19700 20962 19712
rect 21082 19700 21088 19712
rect 20956 19672 21088 19700
rect 20956 19660 20962 19672
rect 21082 19660 21088 19672
rect 21140 19660 21146 19712
rect 21192 19700 21220 19740
rect 23290 19728 23296 19740
rect 23348 19728 23354 19780
rect 24302 19728 24308 19780
rect 24360 19728 24366 19780
rect 24412 19768 24440 19799
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 24670 19768 24676 19780
rect 24412 19740 24676 19768
rect 24670 19728 24676 19740
rect 24728 19728 24734 19780
rect 25222 19768 25228 19780
rect 25183 19740 25228 19768
rect 25222 19728 25228 19740
rect 25280 19728 25286 19780
rect 22738 19700 22744 19712
rect 21192 19672 22744 19700
rect 22738 19660 22744 19672
rect 22796 19660 22802 19712
rect 23937 19703 23995 19709
rect 23937 19669 23949 19703
rect 23983 19700 23995 19703
rect 24118 19700 24124 19712
rect 23983 19672 24124 19700
rect 23983 19669 23995 19672
rect 23937 19663 23995 19669
rect 24118 19660 24124 19672
rect 24176 19660 24182 19712
rect 24320 19700 24348 19728
rect 24949 19703 25007 19709
rect 24949 19700 24961 19703
rect 24320 19672 24961 19700
rect 24949 19669 24961 19672
rect 24995 19700 25007 19703
rect 25958 19700 25964 19712
rect 24995 19672 25964 19700
rect 24995 19669 25007 19672
rect 24949 19663 25007 19669
rect 25958 19660 25964 19672
rect 26016 19660 26022 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 3697 19499 3755 19505
rect 3697 19465 3709 19499
rect 3743 19496 3755 19499
rect 4062 19496 4068 19508
rect 3743 19468 4068 19496
rect 3743 19465 3755 19468
rect 3697 19459 3755 19465
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 5258 19496 5264 19508
rect 5219 19468 5264 19496
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 5350 19456 5356 19508
rect 5408 19496 5414 19508
rect 6454 19496 6460 19508
rect 5408 19468 6460 19496
rect 5408 19456 5414 19468
rect 6454 19456 6460 19468
rect 6512 19456 6518 19508
rect 7006 19496 7012 19508
rect 6967 19468 7012 19496
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 10594 19496 10600 19508
rect 10555 19468 10600 19496
rect 10594 19456 10600 19468
rect 10652 19456 10658 19508
rect 13446 19496 13452 19508
rect 13407 19468 13452 19496
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 14550 19456 14556 19508
rect 14608 19496 14614 19508
rect 15930 19496 15936 19508
rect 14608 19468 15936 19496
rect 14608 19456 14614 19468
rect 15930 19456 15936 19468
rect 15988 19496 15994 19508
rect 16206 19496 16212 19508
rect 15988 19468 16068 19496
rect 16167 19468 16212 19496
rect 15988 19456 15994 19468
rect 3050 19388 3056 19440
rect 3108 19428 3114 19440
rect 3786 19428 3792 19440
rect 3108 19400 3792 19428
rect 3108 19388 3114 19400
rect 3786 19388 3792 19400
rect 3844 19388 3850 19440
rect 6914 19428 6920 19440
rect 5368 19400 6920 19428
rect 4249 19363 4307 19369
rect 4249 19329 4261 19363
rect 4295 19360 4307 19363
rect 4982 19360 4988 19372
rect 4295 19332 4988 19360
rect 4295 19329 4307 19332
rect 4249 19323 4307 19329
rect 4982 19320 4988 19332
rect 5040 19320 5046 19372
rect 2406 19292 2412 19304
rect 2367 19264 2412 19292
rect 2406 19252 2412 19264
rect 2464 19252 2470 19304
rect 3050 19252 3056 19304
rect 3108 19292 3114 19304
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 3108 19264 3433 19292
rect 3108 19252 3114 19264
rect 3421 19261 3433 19264
rect 3467 19292 3479 19295
rect 3973 19295 4031 19301
rect 3973 19292 3985 19295
rect 3467 19264 3985 19292
rect 3467 19261 3479 19264
rect 3421 19255 3479 19261
rect 3973 19261 3985 19264
rect 4019 19261 4031 19295
rect 3973 19255 4031 19261
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4525 19295 4583 19301
rect 4525 19292 4537 19295
rect 4212 19264 4537 19292
rect 4212 19252 4218 19264
rect 4525 19261 4537 19264
rect 4571 19261 4583 19295
rect 5368 19292 5396 19400
rect 6914 19388 6920 19400
rect 6972 19388 6978 19440
rect 9490 19388 9496 19440
rect 9548 19428 9554 19440
rect 11054 19428 11060 19440
rect 9548 19400 11060 19428
rect 9548 19388 9554 19400
rect 11054 19388 11060 19400
rect 11112 19428 11118 19440
rect 11698 19428 11704 19440
rect 11112 19400 11704 19428
rect 11112 19388 11118 19400
rect 11698 19388 11704 19400
rect 11756 19388 11762 19440
rect 11790 19388 11796 19440
rect 11848 19428 11854 19440
rect 11848 19400 11928 19428
rect 11848 19388 11854 19400
rect 5813 19363 5871 19369
rect 5813 19329 5825 19363
rect 5859 19360 5871 19363
rect 6086 19360 6092 19372
rect 5859 19332 6092 19360
rect 5859 19329 5871 19332
rect 5813 19323 5871 19329
rect 6086 19320 6092 19332
rect 6144 19320 6150 19372
rect 6178 19320 6184 19372
rect 6236 19360 6242 19372
rect 6273 19363 6331 19369
rect 6273 19360 6285 19363
rect 6236 19332 6285 19360
rect 6236 19320 6242 19332
rect 6273 19329 6285 19332
rect 6319 19360 6331 19363
rect 6319 19332 6960 19360
rect 6319 19329 6331 19332
rect 6273 19323 6331 19329
rect 5534 19292 5540 19304
rect 4525 19255 4583 19261
rect 4632 19264 5396 19292
rect 5495 19264 5540 19292
rect 1949 19227 2007 19233
rect 1949 19193 1961 19227
rect 1995 19224 2007 19227
rect 2590 19224 2596 19236
rect 1995 19196 2452 19224
rect 2551 19196 2596 19224
rect 1995 19193 2007 19196
rect 1949 19187 2007 19193
rect 2123 19159 2181 19165
rect 2123 19125 2135 19159
rect 2169 19156 2181 19159
rect 2222 19156 2228 19168
rect 2169 19128 2228 19156
rect 2169 19125 2181 19128
rect 2123 19119 2181 19125
rect 2222 19116 2228 19128
rect 2280 19116 2286 19168
rect 2424 19156 2452 19196
rect 2590 19184 2596 19196
rect 2648 19184 2654 19236
rect 2685 19227 2743 19233
rect 2685 19193 2697 19227
rect 2731 19224 2743 19227
rect 4632 19224 4660 19264
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6472 19264 6837 19292
rect 2731 19196 2765 19224
rect 4172 19196 4660 19224
rect 4709 19227 4767 19233
rect 2731 19193 2743 19196
rect 2685 19187 2743 19193
rect 2498 19156 2504 19168
rect 2424 19128 2504 19156
rect 2498 19116 2504 19128
rect 2556 19156 2562 19168
rect 2700 19156 2728 19187
rect 3053 19159 3111 19165
rect 3053 19156 3065 19159
rect 2556 19128 3065 19156
rect 2556 19116 2562 19128
rect 3053 19125 3065 19128
rect 3099 19156 3111 19159
rect 3234 19156 3240 19168
rect 3099 19128 3240 19156
rect 3099 19125 3111 19128
rect 3053 19119 3111 19125
rect 3234 19116 3240 19128
rect 3292 19116 3298 19168
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 4172 19165 4200 19196
rect 4709 19193 4721 19227
rect 4755 19224 4767 19227
rect 5166 19224 5172 19236
rect 4755 19196 5172 19224
rect 4755 19193 4767 19196
rect 4709 19187 4767 19193
rect 5166 19184 5172 19196
rect 5224 19224 5230 19236
rect 6362 19224 6368 19236
rect 5224 19196 6368 19224
rect 5224 19184 5230 19196
rect 6362 19184 6368 19196
rect 6420 19184 6426 19236
rect 4157 19159 4215 19165
rect 4157 19156 4169 19159
rect 4120 19128 4169 19156
rect 4120 19116 4126 19128
rect 4157 19125 4169 19128
rect 4203 19125 4215 19159
rect 4157 19119 4215 19125
rect 4525 19159 4583 19165
rect 4525 19125 4537 19159
rect 4571 19156 4583 19159
rect 4985 19159 5043 19165
rect 4985 19156 4997 19159
rect 4571 19128 4997 19156
rect 4571 19125 4583 19128
rect 4525 19119 4583 19125
rect 4985 19125 4997 19128
rect 5031 19156 5043 19159
rect 5721 19159 5779 19165
rect 5721 19156 5733 19159
rect 5031 19128 5733 19156
rect 5031 19125 5043 19128
rect 4985 19119 5043 19125
rect 5721 19125 5733 19128
rect 5767 19125 5779 19159
rect 5721 19119 5779 19125
rect 5902 19116 5908 19168
rect 5960 19156 5966 19168
rect 6472 19156 6500 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 6932 19292 6960 19332
rect 7837 19295 7895 19301
rect 7837 19292 7849 19295
rect 6932 19264 7849 19292
rect 6825 19255 6883 19261
rect 7837 19261 7849 19264
rect 7883 19292 7895 19295
rect 8021 19295 8079 19301
rect 8021 19292 8033 19295
rect 7883 19264 8033 19292
rect 7883 19261 7895 19264
rect 7837 19255 7895 19261
rect 8021 19261 8033 19264
rect 8067 19261 8079 19295
rect 8021 19255 8079 19261
rect 9950 19252 9956 19304
rect 10008 19292 10014 19304
rect 10321 19295 10379 19301
rect 10321 19292 10333 19295
rect 10008 19264 10333 19292
rect 10008 19252 10014 19264
rect 10321 19261 10333 19264
rect 10367 19292 10379 19295
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 10367 19264 11161 19292
rect 10367 19261 10379 19264
rect 10321 19255 10379 19261
rect 11149 19261 11161 19264
rect 11195 19292 11207 19295
rect 11790 19292 11796 19304
rect 11195 19264 11796 19292
rect 11195 19261 11207 19264
rect 11149 19255 11207 19261
rect 11790 19252 11796 19264
rect 11848 19252 11854 19304
rect 6638 19224 6644 19236
rect 6551 19196 6644 19224
rect 6638 19184 6644 19196
rect 6696 19224 6702 19236
rect 8288 19227 8346 19233
rect 6696 19196 8248 19224
rect 6696 19184 6702 19196
rect 7469 19159 7527 19165
rect 7469 19156 7481 19159
rect 5960 19128 7481 19156
rect 5960 19116 5966 19128
rect 7469 19125 7481 19128
rect 7515 19156 7527 19159
rect 7650 19156 7656 19168
rect 7515 19128 7656 19156
rect 7515 19125 7527 19128
rect 7469 19119 7527 19125
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 8220 19156 8248 19196
rect 8288 19193 8300 19227
rect 8334 19224 8346 19227
rect 8386 19224 8392 19236
rect 8334 19196 8392 19224
rect 8334 19193 8346 19196
rect 8288 19187 8346 19193
rect 8386 19184 8392 19196
rect 8444 19184 8450 19236
rect 10870 19224 10876 19236
rect 10831 19196 10876 19224
rect 10870 19184 10876 19196
rect 10928 19184 10934 19236
rect 11900 19224 11928 19400
rect 12894 19388 12900 19440
rect 12952 19388 12958 19440
rect 14642 19388 14648 19440
rect 14700 19428 14706 19440
rect 15378 19428 15384 19440
rect 14700 19400 15384 19428
rect 14700 19388 14706 19400
rect 15378 19388 15384 19400
rect 15436 19388 15442 19440
rect 16040 19428 16068 19468
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 19426 19456 19432 19508
rect 19484 19496 19490 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19484 19468 19625 19496
rect 19484 19456 19490 19468
rect 19613 19465 19625 19468
rect 19659 19465 19671 19499
rect 19613 19459 19671 19465
rect 20625 19499 20683 19505
rect 20625 19465 20637 19499
rect 20671 19496 20683 19499
rect 21358 19496 21364 19508
rect 20671 19468 21364 19496
rect 20671 19465 20683 19468
rect 20625 19459 20683 19465
rect 16040 19400 17264 19428
rect 12250 19320 12256 19372
rect 12308 19360 12314 19372
rect 12912 19360 12940 19388
rect 12308 19332 12940 19360
rect 12308 19320 12314 19332
rect 16114 19320 16120 19372
rect 16172 19360 16178 19372
rect 16577 19363 16635 19369
rect 16577 19360 16589 19363
rect 16172 19332 16589 19360
rect 16172 19320 16178 19332
rect 16577 19329 16589 19332
rect 16623 19329 16635 19363
rect 16577 19323 16635 19329
rect 17236 19304 17264 19400
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 19610 19360 19616 19372
rect 19392 19332 19616 19360
rect 19392 19320 19398 19332
rect 19610 19320 19616 19332
rect 19668 19320 19674 19372
rect 20732 19369 20760 19468
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 22094 19496 22100 19508
rect 22055 19468 22100 19496
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 23750 19496 23756 19508
rect 23711 19468 23756 19496
rect 23750 19456 23756 19468
rect 23808 19456 23814 19508
rect 24762 19456 24768 19508
rect 24820 19456 24826 19508
rect 22738 19388 22744 19440
rect 22796 19428 22802 19440
rect 23109 19431 23167 19437
rect 23109 19428 23121 19431
rect 22796 19400 23121 19428
rect 22796 19388 22802 19400
rect 23109 19397 23121 19400
rect 23155 19428 23167 19431
rect 24780 19428 24808 19456
rect 25038 19428 25044 19440
rect 23155 19400 24808 19428
rect 24964 19400 25044 19428
rect 23155 19397 23167 19400
rect 23109 19391 23167 19397
rect 20717 19363 20775 19369
rect 20717 19329 20729 19363
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19292 12587 19295
rect 12710 19292 12716 19304
rect 12575 19264 12716 19292
rect 12575 19261 12587 19264
rect 12529 19255 12587 19261
rect 12710 19252 12716 19264
rect 12768 19292 12774 19304
rect 12894 19292 12900 19304
rect 12768 19264 12900 19292
rect 12768 19252 12774 19264
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19261 13691 19295
rect 13633 19255 13691 19261
rect 13900 19295 13958 19301
rect 13900 19261 13912 19295
rect 13946 19292 13958 19295
rect 14366 19292 14372 19304
rect 13946 19264 14372 19292
rect 13946 19261 13958 19264
rect 13900 19255 13958 19261
rect 11256 19196 11928 19224
rect 13648 19224 13676 19255
rect 14366 19252 14372 19264
rect 14424 19292 14430 19304
rect 15565 19295 15623 19301
rect 15565 19292 15577 19295
rect 14424 19264 15577 19292
rect 14424 19252 14430 19264
rect 15565 19261 15577 19264
rect 15611 19292 15623 19295
rect 15930 19292 15936 19304
rect 15611 19264 15936 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 15930 19252 15936 19264
rect 15988 19292 15994 19304
rect 16761 19295 16819 19301
rect 16761 19292 16773 19295
rect 15988 19264 16773 19292
rect 15988 19252 15994 19264
rect 16761 19261 16773 19264
rect 16807 19261 16819 19295
rect 17218 19292 17224 19304
rect 17131 19264 17224 19292
rect 16761 19255 16819 19261
rect 17218 19252 17224 19264
rect 17276 19292 17282 19304
rect 17865 19295 17923 19301
rect 17865 19292 17877 19295
rect 17276 19264 17877 19292
rect 17276 19252 17282 19264
rect 17865 19261 17877 19264
rect 17911 19292 17923 19295
rect 18233 19295 18291 19301
rect 18233 19292 18245 19295
rect 17911 19264 18245 19292
rect 17911 19261 17923 19264
rect 17865 19255 17923 19261
rect 18233 19261 18245 19264
rect 18279 19292 18291 19295
rect 20732 19292 20760 19323
rect 23566 19320 23572 19372
rect 23624 19360 23630 19372
rect 23842 19360 23848 19372
rect 23624 19332 23848 19360
rect 23624 19320 23630 19332
rect 23842 19320 23848 19332
rect 23900 19320 23906 19372
rect 24026 19320 24032 19372
rect 24084 19360 24090 19372
rect 24302 19360 24308 19372
rect 24084 19332 24308 19360
rect 24084 19320 24090 19332
rect 24302 19320 24308 19332
rect 24360 19320 24366 19372
rect 24486 19320 24492 19372
rect 24544 19360 24550 19372
rect 24964 19360 24992 19400
rect 25038 19388 25044 19400
rect 25096 19388 25102 19440
rect 24544 19332 24992 19360
rect 24544 19320 24550 19332
rect 18279 19264 20760 19292
rect 20984 19295 21042 19301
rect 18279 19261 18291 19264
rect 18233 19255 18291 19261
rect 20984 19261 20996 19295
rect 21030 19292 21042 19295
rect 21450 19292 21456 19304
rect 21030 19264 21456 19292
rect 21030 19261 21042 19264
rect 20984 19255 21042 19261
rect 21450 19252 21456 19264
rect 21508 19252 21514 19304
rect 23014 19252 23020 19304
rect 23072 19292 23078 19304
rect 25041 19295 25099 19301
rect 25041 19292 25053 19295
rect 23072 19264 23888 19292
rect 23072 19252 23078 19264
rect 23860 19236 23888 19264
rect 24228 19264 25053 19292
rect 24228 19236 24256 19264
rect 25041 19261 25053 19264
rect 25087 19261 25099 19295
rect 25222 19292 25228 19304
rect 25183 19264 25228 19292
rect 25041 19255 25099 19261
rect 25222 19252 25228 19264
rect 25280 19292 25286 19304
rect 25777 19295 25835 19301
rect 25777 19292 25789 19295
rect 25280 19264 25789 19292
rect 25280 19252 25286 19264
rect 25777 19261 25789 19264
rect 25823 19261 25835 19295
rect 25777 19255 25835 19261
rect 13722 19224 13728 19236
rect 13648 19196 13728 19224
rect 11256 19168 11284 19196
rect 13722 19184 13728 19196
rect 13780 19224 13786 19236
rect 14550 19224 14556 19236
rect 13780 19196 14556 19224
rect 13780 19184 13786 19196
rect 14550 19184 14556 19196
rect 14608 19184 14614 19236
rect 18322 19184 18328 19236
rect 18380 19224 18386 19236
rect 18500 19227 18558 19233
rect 18500 19224 18512 19227
rect 18380 19196 18512 19224
rect 18380 19184 18386 19196
rect 18500 19193 18512 19196
rect 18546 19224 18558 19227
rect 19426 19224 19432 19236
rect 18546 19196 19432 19224
rect 18546 19193 18558 19196
rect 18500 19187 18558 19193
rect 19426 19184 19432 19196
rect 19484 19184 19490 19236
rect 22741 19227 22799 19233
rect 22741 19193 22753 19227
rect 22787 19224 22799 19227
rect 23106 19224 23112 19236
rect 22787 19196 23112 19224
rect 22787 19193 22799 19196
rect 22741 19187 22799 19193
rect 23106 19184 23112 19196
rect 23164 19184 23170 19236
rect 23842 19184 23848 19236
rect 23900 19184 23906 19236
rect 24026 19224 24032 19236
rect 23987 19196 24032 19224
rect 24026 19184 24032 19196
rect 24084 19184 24090 19236
rect 24210 19224 24216 19236
rect 24171 19196 24216 19224
rect 24210 19184 24216 19196
rect 24268 19184 24274 19236
rect 24305 19227 24363 19233
rect 24305 19193 24317 19227
rect 24351 19193 24363 19227
rect 24670 19224 24676 19236
rect 24631 19196 24676 19224
rect 24305 19187 24363 19193
rect 9401 19159 9459 19165
rect 9401 19156 9413 19159
rect 8220 19128 9413 19156
rect 9401 19125 9413 19128
rect 9447 19125 9459 19159
rect 9401 19119 9459 19125
rect 10045 19159 10103 19165
rect 10045 19125 10057 19159
rect 10091 19156 10103 19159
rect 10778 19156 10784 19168
rect 10091 19128 10784 19156
rect 10091 19125 10103 19128
rect 10045 19119 10103 19125
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11054 19156 11060 19168
rect 11015 19128 11060 19156
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 11238 19116 11244 19168
rect 11296 19116 11302 19168
rect 11330 19116 11336 19168
rect 11388 19156 11394 19168
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 11388 19128 11529 19156
rect 11388 19116 11394 19128
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 11517 19119 11575 19125
rect 11606 19116 11612 19168
rect 11664 19156 11670 19168
rect 11885 19159 11943 19165
rect 11885 19156 11897 19159
rect 11664 19128 11897 19156
rect 11664 19116 11670 19128
rect 11885 19125 11897 19128
rect 11931 19125 11943 19159
rect 11885 19119 11943 19125
rect 12713 19159 12771 19165
rect 12713 19125 12725 19159
rect 12759 19156 12771 19159
rect 12802 19156 12808 19168
rect 12759 19128 12808 19156
rect 12759 19125 12771 19128
rect 12713 19119 12771 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13173 19159 13231 19165
rect 13173 19125 13185 19159
rect 13219 19156 13231 19159
rect 13630 19156 13636 19168
rect 13219 19128 13636 19156
rect 13219 19125 13231 19128
rect 13173 19119 13231 19125
rect 13630 19116 13636 19128
rect 13688 19116 13694 19168
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 15013 19159 15071 19165
rect 15013 19156 15025 19159
rect 14056 19128 15025 19156
rect 14056 19116 14062 19128
rect 15013 19125 15025 19128
rect 15059 19125 15071 19159
rect 15013 19119 15071 19125
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15252 19128 16037 19156
rect 15252 19116 15258 19128
rect 16025 19125 16037 19128
rect 16071 19156 16083 19159
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 16071 19128 16681 19156
rect 16071 19125 16083 19128
rect 16025 19119 16083 19125
rect 16669 19125 16681 19128
rect 16715 19156 16727 19159
rect 16850 19156 16856 19168
rect 16715 19128 16856 19156
rect 16715 19125 16727 19128
rect 16669 19119 16727 19125
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 20070 19116 20076 19168
rect 20128 19156 20134 19168
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 20128 19128 20177 19156
rect 20128 19116 20134 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 23474 19156 23480 19168
rect 23435 19128 23480 19156
rect 20165 19119 20223 19125
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 23658 19116 23664 19168
rect 23716 19156 23722 19168
rect 24320 19156 24348 19187
rect 24670 19184 24676 19196
rect 24728 19184 24734 19236
rect 25406 19156 25412 19168
rect 23716 19128 24348 19156
rect 25367 19128 25412 19156
rect 23716 19116 23722 19128
rect 25406 19116 25412 19128
rect 25464 19116 25470 19168
rect 26237 19159 26295 19165
rect 26237 19125 26249 19159
rect 26283 19156 26295 19159
rect 26326 19156 26332 19168
rect 26283 19128 26332 19156
rect 26283 19125 26295 19128
rect 26237 19119 26295 19125
rect 26326 19116 26332 19128
rect 26384 19116 26390 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1394 18912 1400 18964
rect 1452 18952 1458 18964
rect 2483 18955 2541 18961
rect 2483 18952 2495 18955
rect 1452 18924 2495 18952
rect 1452 18912 1458 18924
rect 2483 18921 2495 18924
rect 2529 18921 2541 18955
rect 2483 18915 2541 18921
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 3878 18952 3884 18964
rect 3007 18924 3884 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 3068 18896 3096 18924
rect 3878 18912 3884 18924
rect 3936 18912 3942 18964
rect 4709 18955 4767 18961
rect 4709 18921 4721 18955
rect 4755 18952 4767 18955
rect 4982 18952 4988 18964
rect 4755 18924 4988 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 4982 18912 4988 18924
rect 5040 18912 5046 18964
rect 5994 18952 6000 18964
rect 5955 18924 6000 18952
rect 5994 18912 6000 18924
rect 6052 18912 6058 18964
rect 6089 18955 6147 18961
rect 6089 18921 6101 18955
rect 6135 18952 6147 18955
rect 9125 18955 9183 18961
rect 6135 18924 8708 18952
rect 6135 18921 6147 18924
rect 6089 18915 6147 18921
rect 1949 18887 2007 18893
rect 1949 18853 1961 18887
rect 1995 18884 2007 18887
rect 2866 18884 2872 18896
rect 1995 18856 2872 18884
rect 1995 18853 2007 18856
rect 1949 18847 2007 18853
rect 2866 18844 2872 18856
rect 2924 18844 2930 18896
rect 3050 18844 3056 18896
rect 3108 18844 3114 18896
rect 3697 18887 3755 18893
rect 3697 18853 3709 18887
rect 3743 18884 3755 18887
rect 4062 18884 4068 18896
rect 3743 18856 4068 18884
rect 3743 18853 3755 18856
rect 3697 18847 3755 18853
rect 4062 18844 4068 18856
rect 4120 18844 4126 18896
rect 5258 18884 5264 18896
rect 5219 18856 5264 18884
rect 5258 18844 5264 18856
rect 5316 18844 5322 18896
rect 5442 18884 5448 18896
rect 5403 18856 5448 18884
rect 5442 18844 5448 18856
rect 5500 18884 5506 18896
rect 6270 18884 6276 18896
rect 5500 18856 6276 18884
rect 5500 18844 5506 18856
rect 6270 18844 6276 18856
rect 6328 18844 6334 18896
rect 6454 18844 6460 18896
rect 6512 18884 6518 18896
rect 7009 18887 7067 18893
rect 7009 18884 7021 18887
rect 6512 18856 7021 18884
rect 6512 18844 6518 18856
rect 7009 18853 7021 18856
rect 7055 18884 7067 18887
rect 7282 18884 7288 18896
rect 7055 18856 7288 18884
rect 7055 18853 7067 18856
rect 7009 18847 7067 18853
rect 7282 18844 7288 18856
rect 7340 18844 7346 18896
rect 8110 18844 8116 18896
rect 8168 18884 8174 18896
rect 8570 18884 8576 18896
rect 8168 18856 8576 18884
rect 8168 18844 8174 18856
rect 8570 18844 8576 18856
rect 8628 18844 8634 18896
rect 4430 18776 4436 18828
rect 4488 18816 4494 18828
rect 4982 18816 4988 18828
rect 4488 18788 4988 18816
rect 4488 18776 4494 18788
rect 4982 18776 4988 18788
rect 5040 18776 5046 18828
rect 5902 18816 5908 18828
rect 5092 18788 5908 18816
rect 1397 18751 1455 18757
rect 1397 18717 1409 18751
rect 1443 18748 1455 18751
rect 2038 18748 2044 18760
rect 1443 18720 2044 18748
rect 1443 18717 1455 18720
rect 1397 18711 1455 18717
rect 2038 18708 2044 18720
rect 2096 18708 2102 18760
rect 2866 18748 2872 18760
rect 2827 18720 2872 18748
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18717 3111 18751
rect 3053 18711 3111 18717
rect 2317 18683 2375 18689
rect 2317 18649 2329 18683
rect 2363 18680 2375 18683
rect 3068 18680 3096 18711
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 5092 18748 5120 18788
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 7190 18816 7196 18828
rect 7024 18788 7196 18816
rect 5534 18748 5540 18760
rect 3476 18720 5120 18748
rect 5495 18720 5540 18748
rect 3476 18708 3482 18720
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 7024 18757 7052 18788
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18717 7067 18751
rect 7009 18711 7067 18717
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 2363 18652 4559 18680
rect 2363 18649 2375 18652
rect 2317 18643 2375 18649
rect 4341 18615 4399 18621
rect 4341 18581 4353 18615
rect 4387 18612 4399 18615
rect 4430 18612 4436 18624
rect 4387 18584 4436 18612
rect 4387 18581 4399 18584
rect 4341 18575 4399 18581
rect 4430 18572 4436 18584
rect 4488 18572 4494 18624
rect 4531 18612 4559 18652
rect 4798 18640 4804 18692
rect 4856 18680 4862 18692
rect 4985 18683 5043 18689
rect 4985 18680 4997 18683
rect 4856 18652 4997 18680
rect 4856 18640 4862 18652
rect 4985 18649 4997 18652
rect 5031 18649 5043 18683
rect 4985 18643 5043 18649
rect 6270 18640 6276 18692
rect 6328 18680 6334 18692
rect 6365 18683 6423 18689
rect 6365 18680 6377 18683
rect 6328 18652 6377 18680
rect 6328 18640 6334 18652
rect 6365 18649 6377 18652
rect 6411 18680 6423 18683
rect 7116 18680 7144 18711
rect 7466 18708 7472 18760
rect 7524 18748 7530 18760
rect 8478 18748 8484 18760
rect 7524 18720 8156 18748
rect 8439 18720 8484 18748
rect 7524 18708 7530 18720
rect 8128 18689 8156 18720
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 8680 18757 8708 18924
rect 9125 18921 9137 18955
rect 9171 18952 9183 18955
rect 9582 18952 9588 18964
rect 9171 18924 9588 18952
rect 9171 18921 9183 18924
rect 9125 18915 9183 18921
rect 9582 18912 9588 18924
rect 9640 18912 9646 18964
rect 11790 18952 11796 18964
rect 11751 18924 11796 18952
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 13722 18912 13728 18964
rect 13780 18952 13786 18964
rect 13909 18955 13967 18961
rect 13909 18952 13921 18955
rect 13780 18924 13921 18952
rect 13780 18912 13786 18924
rect 13909 18921 13921 18924
rect 13955 18921 13967 18955
rect 13909 18915 13967 18921
rect 16393 18955 16451 18961
rect 16393 18921 16405 18955
rect 16439 18952 16451 18955
rect 16482 18952 16488 18964
rect 16439 18924 16488 18952
rect 16439 18921 16451 18924
rect 16393 18915 16451 18921
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 18138 18952 18144 18964
rect 18099 18924 18144 18952
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 19426 18952 19432 18964
rect 19076 18924 19432 18952
rect 9493 18887 9551 18893
rect 9493 18853 9505 18887
rect 9539 18884 9551 18887
rect 10870 18884 10876 18896
rect 9539 18856 10876 18884
rect 9539 18853 9551 18856
rect 9493 18847 9551 18853
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 13446 18884 13452 18896
rect 13407 18856 13452 18884
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 15841 18887 15899 18893
rect 15841 18853 15853 18887
rect 15887 18884 15899 18887
rect 16206 18884 16212 18896
rect 15887 18856 16212 18884
rect 15887 18853 15899 18856
rect 15841 18847 15899 18853
rect 16206 18844 16212 18856
rect 16264 18844 16270 18896
rect 17402 18884 17408 18896
rect 17363 18856 17408 18884
rect 17402 18844 17408 18856
rect 17460 18844 17466 18896
rect 18966 18884 18972 18896
rect 18927 18856 18972 18884
rect 18966 18844 18972 18856
rect 19024 18844 19030 18896
rect 19076 18893 19104 18924
rect 19426 18912 19432 18924
rect 19484 18952 19490 18964
rect 19889 18955 19947 18961
rect 19889 18952 19901 18955
rect 19484 18924 19901 18952
rect 19484 18912 19490 18924
rect 19889 18921 19901 18924
rect 19935 18952 19947 18955
rect 19978 18952 19984 18964
rect 19935 18924 19984 18952
rect 19935 18921 19947 18924
rect 19889 18915 19947 18921
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20717 18955 20775 18961
rect 20717 18921 20729 18955
rect 20763 18952 20775 18955
rect 21542 18952 21548 18964
rect 20763 18924 21548 18952
rect 20763 18921 20775 18924
rect 20717 18915 20775 18921
rect 21542 18912 21548 18924
rect 21600 18912 21606 18964
rect 22005 18955 22063 18961
rect 22005 18921 22017 18955
rect 22051 18952 22063 18955
rect 22094 18952 22100 18964
rect 22051 18924 22100 18952
rect 22051 18921 22063 18924
rect 22005 18915 22063 18921
rect 22094 18912 22100 18924
rect 22152 18912 22158 18964
rect 24026 18912 24032 18964
rect 24084 18952 24090 18964
rect 25409 18955 25467 18961
rect 25409 18952 25421 18955
rect 24084 18924 25421 18952
rect 24084 18912 24090 18924
rect 25409 18921 25421 18924
rect 25455 18921 25467 18955
rect 25409 18915 25467 18921
rect 19061 18887 19119 18893
rect 19061 18853 19073 18887
rect 19107 18853 19119 18887
rect 19061 18847 19119 18853
rect 19518 18844 19524 18896
rect 19576 18884 19582 18896
rect 20070 18884 20076 18896
rect 19576 18856 20076 18884
rect 19576 18844 19582 18856
rect 20070 18844 20076 18856
rect 20128 18884 20134 18896
rect 20165 18887 20223 18893
rect 20165 18884 20177 18887
rect 20128 18856 20177 18884
rect 20128 18844 20134 18856
rect 20165 18853 20177 18856
rect 20211 18853 20223 18887
rect 20165 18847 20223 18853
rect 10680 18819 10738 18825
rect 10680 18785 10692 18819
rect 10726 18816 10738 18819
rect 11790 18816 11796 18828
rect 10726 18788 11796 18816
rect 10726 18785 10738 18788
rect 10680 18779 10738 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 12308 18788 13553 18816
rect 12308 18776 12314 18788
rect 13541 18785 13553 18788
rect 13587 18785 13599 18819
rect 15102 18816 15108 18828
rect 15063 18788 15108 18816
rect 13541 18779 13599 18785
rect 15102 18776 15108 18788
rect 15160 18776 15166 18828
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 15930 18816 15936 18828
rect 15891 18788 15936 18816
rect 15930 18776 15936 18788
rect 15988 18816 15994 18828
rect 16669 18819 16727 18825
rect 16669 18816 16681 18819
rect 15988 18788 16681 18816
rect 15988 18776 15994 18788
rect 16669 18785 16681 18788
rect 16715 18816 16727 18819
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 16715 18788 17509 18816
rect 16715 18785 16727 18788
rect 16669 18779 16727 18785
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 18506 18776 18512 18828
rect 18564 18816 18570 18828
rect 18785 18819 18843 18825
rect 18785 18816 18797 18819
rect 18564 18788 18797 18816
rect 18564 18776 18570 18788
rect 18785 18785 18797 18788
rect 18831 18785 18843 18819
rect 20180 18816 20208 18847
rect 20530 18844 20536 18896
rect 20588 18884 20594 18896
rect 21450 18884 21456 18896
rect 20588 18856 21456 18884
rect 20588 18844 20594 18856
rect 21450 18844 21456 18856
rect 21508 18844 21514 18896
rect 22278 18844 22284 18896
rect 22336 18884 22342 18896
rect 22738 18884 22744 18896
rect 22336 18856 22744 18884
rect 22336 18844 22342 18856
rect 22738 18844 22744 18856
rect 22796 18844 22802 18896
rect 23014 18884 23020 18896
rect 22975 18856 23020 18884
rect 23014 18844 23020 18856
rect 23072 18844 23078 18896
rect 24581 18887 24639 18893
rect 24581 18853 24593 18887
rect 24627 18884 24639 18887
rect 24670 18884 24676 18896
rect 24627 18856 24676 18884
rect 24627 18853 24639 18856
rect 24581 18847 24639 18853
rect 24670 18844 24676 18856
rect 24728 18844 24734 18896
rect 25038 18884 25044 18896
rect 24999 18856 25044 18884
rect 25038 18844 25044 18856
rect 25096 18844 25102 18896
rect 21545 18819 21603 18825
rect 21545 18816 21557 18819
rect 20180 18788 21557 18816
rect 18785 18779 18843 18785
rect 21545 18785 21557 18788
rect 21591 18816 21603 18819
rect 22370 18816 22376 18828
rect 21591 18788 22376 18816
rect 21591 18785 21603 18788
rect 21545 18779 21603 18785
rect 22370 18776 22376 18788
rect 22428 18816 22434 18828
rect 23109 18819 23167 18825
rect 23109 18816 23121 18819
rect 22428 18788 23121 18816
rect 22428 18776 22434 18788
rect 23109 18785 23121 18788
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 8665 18751 8723 18757
rect 8665 18717 8677 18751
rect 8711 18748 8723 18751
rect 9490 18748 9496 18760
rect 8711 18720 9496 18748
rect 8711 18717 8723 18720
rect 8665 18711 8723 18717
rect 9490 18708 9496 18720
rect 9548 18708 9554 18760
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 10134 18748 10140 18760
rect 9824 18720 10140 18748
rect 9824 18708 9830 18720
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10226 18708 10232 18760
rect 10284 18748 10290 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 10284 18720 10425 18748
rect 10284 18708 10290 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 10413 18711 10471 18717
rect 12728 18720 13369 18748
rect 6411 18652 7144 18680
rect 8113 18683 8171 18689
rect 6411 18649 6423 18652
rect 6365 18643 6423 18649
rect 8113 18649 8125 18683
rect 8159 18649 8171 18683
rect 8113 18643 8171 18649
rect 12728 18624 12756 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13906 18708 13912 18760
rect 13964 18748 13970 18760
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 13964 18720 14657 18748
rect 13964 18708 13970 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 17310 18748 17316 18760
rect 17271 18720 17316 18748
rect 14645 18711 14703 18717
rect 17310 18708 17316 18720
rect 17368 18708 17374 18760
rect 17770 18708 17776 18760
rect 17828 18748 17834 18760
rect 20898 18748 20904 18760
rect 17828 18720 20904 18748
rect 17828 18708 17834 18720
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 21450 18748 21456 18760
rect 21411 18720 21456 18748
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22060 18720 22937 18748
rect 22060 18708 22066 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 22925 18711 22983 18717
rect 24210 18708 24216 18760
rect 24268 18748 24274 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24268 18720 24593 18748
rect 24268 18708 24274 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18748 24731 18751
rect 24854 18748 24860 18760
rect 24719 18720 24860 18748
rect 24719 18717 24731 18720
rect 24673 18711 24731 18717
rect 12894 18640 12900 18692
rect 12952 18680 12958 18692
rect 15378 18680 15384 18692
rect 12952 18652 14412 18680
rect 15339 18652 15384 18680
rect 12952 18640 12958 18652
rect 6089 18615 6147 18621
rect 6089 18612 6101 18615
rect 4531 18584 6101 18612
rect 6089 18581 6101 18584
rect 6135 18581 6147 18615
rect 6089 18575 6147 18581
rect 6549 18615 6607 18621
rect 6549 18581 6561 18615
rect 6595 18612 6607 18615
rect 6638 18612 6644 18624
rect 6595 18584 6644 18612
rect 6595 18581 6607 18584
rect 6549 18575 6607 18581
rect 6638 18572 6644 18584
rect 6696 18572 6702 18624
rect 7466 18612 7472 18624
rect 7427 18584 7472 18612
rect 7466 18572 7472 18584
rect 7524 18572 7530 18624
rect 7834 18612 7840 18624
rect 7795 18584 7840 18612
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 9950 18612 9956 18624
rect 9911 18584 9956 18612
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10134 18572 10140 18624
rect 10192 18612 10198 18624
rect 10229 18615 10287 18621
rect 10229 18612 10241 18615
rect 10192 18584 10241 18612
rect 10192 18572 10198 18584
rect 10229 18581 10241 18584
rect 10275 18581 10287 18615
rect 10229 18575 10287 18581
rect 12250 18572 12256 18624
rect 12308 18612 12314 18624
rect 12434 18612 12440 18624
rect 12308 18584 12440 18612
rect 12308 18572 12314 18584
rect 12434 18572 12440 18584
rect 12492 18572 12498 18624
rect 12710 18612 12716 18624
rect 12671 18584 12716 18612
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 12989 18615 13047 18621
rect 12989 18581 13001 18615
rect 13035 18612 13047 18615
rect 13722 18612 13728 18624
rect 13035 18584 13728 18612
rect 13035 18581 13047 18584
rect 12989 18575 13047 18581
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 13998 18572 14004 18624
rect 14056 18612 14062 18624
rect 14277 18615 14335 18621
rect 14277 18612 14289 18615
rect 14056 18584 14289 18612
rect 14056 18572 14062 18584
rect 14277 18581 14289 18584
rect 14323 18581 14335 18615
rect 14384 18612 14412 18652
rect 15378 18640 15384 18652
rect 15436 18640 15442 18692
rect 16942 18680 16948 18692
rect 16903 18652 16948 18680
rect 16942 18640 16948 18652
rect 17000 18640 17006 18692
rect 18509 18683 18567 18689
rect 18509 18649 18521 18683
rect 18555 18680 18567 18683
rect 19242 18680 19248 18692
rect 18555 18652 19248 18680
rect 18555 18649 18567 18652
rect 18509 18643 18567 18649
rect 19242 18640 19248 18652
rect 19300 18640 19306 18692
rect 20990 18680 20996 18692
rect 20951 18652 20996 18680
rect 20990 18640 20996 18652
rect 21048 18640 21054 18692
rect 22557 18683 22615 18689
rect 22557 18649 22569 18683
rect 22603 18680 22615 18683
rect 22830 18680 22836 18692
rect 22603 18652 22836 18680
rect 22603 18649 22615 18652
rect 22557 18643 22615 18649
rect 22830 18640 22836 18652
rect 22888 18640 22894 18692
rect 24026 18640 24032 18692
rect 24084 18680 24090 18692
rect 24302 18680 24308 18692
rect 24084 18652 24308 18680
rect 24084 18640 24090 18652
rect 24302 18640 24308 18652
rect 24360 18640 24366 18692
rect 24394 18640 24400 18692
rect 24452 18640 24458 18692
rect 24596 18680 24624 18711
rect 24854 18708 24860 18720
rect 24912 18748 24918 18760
rect 25038 18748 25044 18760
rect 24912 18720 25044 18748
rect 24912 18708 24918 18720
rect 25038 18708 25044 18720
rect 25096 18708 25102 18760
rect 26418 18680 26424 18692
rect 24596 18652 26424 18680
rect 26418 18640 26424 18652
rect 26476 18640 26482 18692
rect 15470 18612 15476 18624
rect 14384 18584 15476 18612
rect 14277 18575 14335 18581
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 19521 18615 19579 18621
rect 19521 18581 19533 18615
rect 19567 18612 19579 18615
rect 19978 18612 19984 18624
rect 19567 18584 19984 18612
rect 19567 18581 19579 18584
rect 19521 18575 19579 18581
rect 19978 18572 19984 18584
rect 20036 18612 20042 18624
rect 20346 18612 20352 18624
rect 20036 18584 20352 18612
rect 20036 18572 20042 18584
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 22370 18612 22376 18624
rect 22331 18584 22376 18612
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 23658 18612 23664 18624
rect 23619 18584 23664 18612
rect 23658 18572 23664 18584
rect 23716 18572 23722 18624
rect 24121 18615 24179 18621
rect 24121 18581 24133 18615
rect 24167 18612 24179 18615
rect 24412 18612 24440 18640
rect 24167 18584 24440 18612
rect 24167 18581 24179 18584
rect 24121 18575 24179 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2225 18411 2283 18417
rect 2225 18377 2237 18411
rect 2271 18408 2283 18411
rect 3050 18408 3056 18420
rect 2271 18380 3056 18408
rect 2271 18377 2283 18380
rect 2225 18371 2283 18377
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 3786 18408 3792 18420
rect 3747 18380 3792 18408
rect 3786 18368 3792 18380
rect 3844 18368 3850 18420
rect 4157 18411 4215 18417
rect 4157 18377 4169 18411
rect 4203 18408 4215 18411
rect 5166 18408 5172 18420
rect 4203 18380 5172 18408
rect 4203 18377 4215 18380
rect 4157 18371 4215 18377
rect 2774 18300 2780 18352
rect 2832 18340 2838 18352
rect 2832 18312 2877 18340
rect 2832 18300 2838 18312
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 2593 18275 2651 18281
rect 2593 18272 2605 18275
rect 1636 18244 2605 18272
rect 1636 18232 1642 18244
rect 2593 18241 2605 18244
rect 2639 18272 2651 18275
rect 3234 18272 3240 18284
rect 2639 18244 3240 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 4264 18281 4292 18380
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 6273 18411 6331 18417
rect 6273 18377 6285 18411
rect 6319 18408 6331 18411
rect 6454 18408 6460 18420
rect 6319 18380 6460 18408
rect 6319 18377 6331 18380
rect 6273 18371 6331 18377
rect 6454 18368 6460 18380
rect 6512 18368 6518 18420
rect 8110 18408 8116 18420
rect 8071 18380 8116 18408
rect 8110 18368 8116 18380
rect 8168 18368 8174 18420
rect 8294 18368 8300 18420
rect 8352 18408 8358 18420
rect 8573 18411 8631 18417
rect 8573 18408 8585 18411
rect 8352 18380 8585 18408
rect 8352 18368 8358 18380
rect 8573 18377 8585 18380
rect 8619 18377 8631 18411
rect 8573 18371 8631 18377
rect 9769 18411 9827 18417
rect 9769 18377 9781 18411
rect 9815 18408 9827 18411
rect 10226 18408 10232 18420
rect 9815 18380 10232 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 5442 18300 5448 18352
rect 5500 18340 5506 18352
rect 6917 18343 6975 18349
rect 6917 18340 6929 18343
rect 5500 18312 6929 18340
rect 5500 18300 5506 18312
rect 6917 18309 6929 18312
rect 6963 18309 6975 18343
rect 7650 18340 7656 18352
rect 6917 18303 6975 18309
rect 7024 18312 7656 18340
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18241 4307 18275
rect 4249 18235 4307 18241
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 7024 18272 7052 18312
rect 7650 18300 7656 18312
rect 7708 18300 7714 18352
rect 7466 18272 7472 18284
rect 5316 18244 7052 18272
rect 7427 18244 7472 18272
rect 5316 18232 5322 18244
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 9876 18281 9904 18380
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 11054 18368 11060 18420
rect 11112 18408 11118 18420
rect 12529 18411 12587 18417
rect 12529 18408 12541 18411
rect 11112 18380 12541 18408
rect 11112 18368 11118 18380
rect 12529 18377 12541 18380
rect 12575 18377 12587 18411
rect 13446 18408 13452 18420
rect 13407 18380 13452 18408
rect 12529 18371 12587 18377
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 14185 18411 14243 18417
rect 14185 18377 14197 18411
rect 14231 18408 14243 18411
rect 14550 18408 14556 18420
rect 14231 18380 14556 18408
rect 14231 18377 14243 18380
rect 14185 18371 14243 18377
rect 10870 18300 10876 18352
rect 10928 18300 10934 18352
rect 12618 18300 12624 18352
rect 12676 18340 12682 18352
rect 13078 18340 13084 18352
rect 12676 18312 13084 18340
rect 12676 18300 12682 18312
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18241 9919 18275
rect 10888 18272 10916 18300
rect 14292 18284 14320 18380
rect 14550 18368 14556 18380
rect 14608 18368 14614 18420
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 15344 18380 15669 18408
rect 15344 18368 15350 18380
rect 15657 18377 15669 18380
rect 15703 18408 15715 18411
rect 15930 18408 15936 18420
rect 15703 18380 15936 18408
rect 15703 18377 15715 18380
rect 15657 18371 15715 18377
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 17034 18408 17040 18420
rect 16995 18380 17040 18408
rect 17034 18368 17040 18380
rect 17092 18368 17098 18420
rect 18966 18368 18972 18420
rect 19024 18408 19030 18420
rect 19061 18411 19119 18417
rect 19061 18408 19073 18411
rect 19024 18380 19073 18408
rect 19024 18368 19030 18380
rect 19061 18377 19073 18380
rect 19107 18377 19119 18411
rect 19426 18408 19432 18420
rect 19387 18380 19432 18408
rect 19061 18371 19119 18377
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 21358 18408 21364 18420
rect 19536 18380 21036 18408
rect 21319 18380 21364 18408
rect 18138 18340 18144 18352
rect 18099 18312 18144 18340
rect 18138 18300 18144 18312
rect 18196 18300 18202 18352
rect 18690 18300 18696 18352
rect 18748 18340 18754 18352
rect 19536 18340 19564 18380
rect 18748 18312 19564 18340
rect 21008 18340 21036 18380
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 21450 18368 21456 18420
rect 21508 18408 21514 18420
rect 21913 18411 21971 18417
rect 21913 18408 21925 18411
rect 21508 18380 21925 18408
rect 21508 18368 21514 18380
rect 21913 18377 21925 18380
rect 21959 18377 21971 18411
rect 21913 18371 21971 18377
rect 22002 18368 22008 18420
rect 22060 18408 22066 18420
rect 22189 18411 22247 18417
rect 22189 18408 22201 18411
rect 22060 18380 22201 18408
rect 22060 18368 22066 18380
rect 22189 18377 22201 18380
rect 22235 18377 22247 18411
rect 22646 18408 22652 18420
rect 22607 18380 22652 18408
rect 22189 18371 22247 18377
rect 22646 18368 22652 18380
rect 22704 18368 22710 18420
rect 23477 18411 23535 18417
rect 23477 18377 23489 18411
rect 23523 18408 23535 18411
rect 23658 18408 23664 18420
rect 23523 18380 23664 18408
rect 23523 18377 23535 18380
rect 23477 18371 23535 18377
rect 23658 18368 23664 18380
rect 23716 18408 23722 18420
rect 24210 18408 24216 18420
rect 23716 18380 24216 18408
rect 23716 18368 23722 18380
rect 24210 18368 24216 18380
rect 24268 18368 24274 18420
rect 25038 18408 25044 18420
rect 24999 18380 25044 18408
rect 25038 18368 25044 18380
rect 25096 18368 25102 18420
rect 25409 18411 25467 18417
rect 25409 18377 25421 18411
rect 25455 18408 25467 18411
rect 25590 18408 25596 18420
rect 25455 18380 25596 18408
rect 25455 18377 25467 18380
rect 25409 18371 25467 18377
rect 25590 18368 25596 18380
rect 25648 18368 25654 18420
rect 25774 18408 25780 18420
rect 25735 18380 25780 18408
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 23753 18343 23811 18349
rect 23753 18340 23765 18343
rect 21008 18312 23765 18340
rect 18748 18300 18754 18312
rect 23753 18309 23765 18312
rect 23799 18309 23811 18343
rect 26234 18340 26240 18352
rect 26195 18312 26240 18340
rect 23753 18303 23811 18309
rect 26234 18300 26240 18312
rect 26292 18300 26298 18352
rect 11054 18272 11060 18284
rect 10888 18244 11060 18272
rect 9861 18235 9919 18241
rect 1394 18204 1400 18216
rect 1355 18176 1400 18204
rect 1394 18164 1400 18176
rect 1452 18164 1458 18216
rect 6362 18164 6368 18216
rect 6420 18204 6426 18216
rect 6641 18207 6699 18213
rect 6641 18204 6653 18207
rect 6420 18176 6653 18204
rect 6420 18164 6426 18176
rect 6641 18173 6653 18176
rect 6687 18204 6699 18207
rect 8389 18207 8447 18213
rect 6687 18176 7420 18204
rect 6687 18173 6699 18176
rect 6641 18167 6699 18173
rect 7392 18148 7420 18176
rect 8389 18173 8401 18207
rect 8435 18204 8447 18207
rect 8435 18176 9076 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 1578 18096 1584 18148
rect 1636 18136 1642 18148
rect 1673 18139 1731 18145
rect 1673 18136 1685 18139
rect 1636 18108 1685 18136
rect 1636 18096 1642 18108
rect 1673 18105 1685 18108
rect 1719 18105 1731 18139
rect 1673 18099 1731 18105
rect 3050 18096 3056 18148
rect 3108 18136 3114 18148
rect 3329 18139 3387 18145
rect 3329 18136 3341 18139
rect 3108 18108 3341 18136
rect 3108 18096 3114 18108
rect 3329 18105 3341 18108
rect 3375 18105 3387 18139
rect 3329 18099 3387 18105
rect 4516 18139 4574 18145
rect 4516 18105 4528 18139
rect 4562 18136 4574 18139
rect 5442 18136 5448 18148
rect 4562 18108 5448 18136
rect 4562 18105 4574 18108
rect 4516 18099 4574 18105
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 3602 18068 3608 18080
rect 3283 18040 3608 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 3602 18028 3608 18040
rect 3660 18028 3666 18080
rect 4430 18028 4436 18080
rect 4488 18068 4494 18080
rect 4531 18068 4559 18099
rect 5442 18096 5448 18108
rect 5500 18096 5506 18148
rect 6822 18096 6828 18148
rect 6880 18136 6886 18148
rect 7193 18139 7251 18145
rect 7193 18136 7205 18139
rect 6880 18108 7205 18136
rect 6880 18096 6886 18108
rect 7193 18105 7205 18108
rect 7239 18105 7251 18139
rect 7374 18136 7380 18148
rect 7335 18108 7380 18136
rect 7193 18099 7251 18105
rect 7374 18096 7380 18108
rect 7432 18096 7438 18148
rect 4488 18040 4559 18068
rect 4488 18028 4494 18040
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 9048 18077 9076 18176
rect 5629 18071 5687 18077
rect 5629 18068 5641 18071
rect 5592 18040 5641 18068
rect 5592 18028 5598 18040
rect 5629 18037 5641 18040
rect 5675 18037 5687 18071
rect 5629 18031 5687 18037
rect 9033 18071 9091 18077
rect 9033 18037 9045 18071
rect 9079 18068 9091 18071
rect 9306 18068 9312 18080
rect 9079 18040 9312 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18068 9459 18071
rect 9490 18068 9496 18080
rect 9447 18040 9496 18068
rect 9447 18037 9459 18040
rect 9401 18031 9459 18037
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 9582 18028 9588 18080
rect 9640 18068 9646 18080
rect 9876 18068 9904 18235
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11422 18232 11428 18284
rect 11480 18272 11486 18284
rect 11977 18275 12035 18281
rect 11977 18272 11989 18275
rect 11480 18244 11989 18272
rect 11480 18232 11486 18244
rect 11977 18241 11989 18244
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18272 13047 18275
rect 13354 18272 13360 18284
rect 13035 18244 13360 18272
rect 13035 18241 13047 18244
rect 12989 18235 13047 18241
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 14274 18272 14280 18284
rect 14187 18244 14280 18272
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 16114 18232 16120 18284
rect 16172 18272 16178 18284
rect 16298 18272 16304 18284
rect 16172 18244 16304 18272
rect 16172 18232 16178 18244
rect 16298 18232 16304 18244
rect 16356 18272 16362 18284
rect 17402 18272 17408 18284
rect 16356 18244 17408 18272
rect 16356 18232 16362 18244
rect 17402 18232 17408 18244
rect 17460 18272 17466 18284
rect 17773 18275 17831 18281
rect 17773 18272 17785 18275
rect 17460 18244 17785 18272
rect 17460 18232 17466 18244
rect 17773 18241 17785 18244
rect 17819 18241 17831 18275
rect 18598 18272 18604 18284
rect 18559 18244 18604 18272
rect 17773 18235 17831 18241
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 23842 18232 23848 18284
rect 23900 18272 23906 18284
rect 24305 18275 24363 18281
rect 24305 18272 24317 18275
rect 23900 18244 24317 18272
rect 23900 18232 23906 18244
rect 24305 18241 24317 18244
rect 24351 18272 24363 18275
rect 24854 18272 24860 18284
rect 24351 18244 24860 18272
rect 24351 18241 24363 18244
rect 24305 18235 24363 18241
rect 24854 18232 24860 18244
rect 24912 18232 24918 18284
rect 10594 18164 10600 18216
rect 10652 18204 10658 18216
rect 10870 18204 10876 18216
rect 10652 18176 10876 18204
rect 10652 18164 10658 18176
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 13081 18207 13139 18213
rect 13081 18204 13093 18207
rect 11808 18176 13093 18204
rect 9950 18096 9956 18148
rect 10008 18136 10014 18148
rect 10128 18139 10186 18145
rect 10128 18136 10140 18139
rect 10008 18108 10140 18136
rect 10008 18096 10014 18108
rect 10128 18105 10140 18108
rect 10174 18136 10186 18139
rect 10686 18136 10692 18148
rect 10174 18108 10692 18136
rect 10174 18105 10186 18108
rect 10128 18099 10186 18105
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 11808 18080 11836 18176
rect 13081 18173 13093 18176
rect 13127 18173 13139 18207
rect 13081 18167 13139 18173
rect 16853 18207 16911 18213
rect 16853 18173 16865 18207
rect 16899 18173 16911 18207
rect 16853 18167 16911 18173
rect 14550 18145 14556 18148
rect 14544 18136 14556 18145
rect 14511 18108 14556 18136
rect 14544 18099 14556 18108
rect 14550 18096 14556 18099
rect 14608 18096 14614 18148
rect 9640 18040 9904 18068
rect 9640 18028 9646 18040
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 11146 18068 11152 18080
rect 10836 18040 11152 18068
rect 10836 18028 10842 18040
rect 11146 18028 11152 18040
rect 11204 18068 11210 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 11204 18040 11253 18068
rect 11204 18028 11210 18040
rect 11241 18037 11253 18040
rect 11287 18037 11299 18071
rect 11790 18068 11796 18080
rect 11751 18040 11796 18068
rect 11241 18031 11299 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 11977 18071 12035 18077
rect 11977 18037 11989 18071
rect 12023 18068 12035 18071
rect 12253 18071 12311 18077
rect 12253 18068 12265 18071
rect 12023 18040 12265 18068
rect 12023 18037 12035 18040
rect 11977 18031 12035 18037
rect 12253 18037 12265 18040
rect 12299 18068 12311 18071
rect 12989 18071 13047 18077
rect 12989 18068 13001 18071
rect 12299 18040 13001 18068
rect 12299 18037 12311 18040
rect 12253 18031 12311 18037
rect 12989 18037 13001 18040
rect 13035 18068 13047 18071
rect 15378 18068 15384 18080
rect 13035 18040 15384 18068
rect 13035 18037 13047 18040
rect 12989 18031 13047 18037
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 16206 18068 16212 18080
rect 16167 18040 16212 18068
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16761 18071 16819 18077
rect 16761 18037 16773 18071
rect 16807 18068 16819 18071
rect 16868 18068 16896 18167
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 18693 18207 18751 18213
rect 18693 18204 18705 18207
rect 18288 18176 18705 18204
rect 18288 18164 18294 18176
rect 18693 18173 18705 18176
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 19981 18207 20039 18213
rect 19981 18173 19993 18207
rect 20027 18173 20039 18207
rect 19981 18167 20039 18173
rect 17402 18068 17408 18080
rect 16807 18040 17408 18068
rect 16807 18037 16819 18040
rect 16761 18031 16819 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 18601 18071 18659 18077
rect 18601 18037 18613 18071
rect 18647 18068 18659 18071
rect 18782 18068 18788 18080
rect 18647 18040 18788 18068
rect 18647 18037 18659 18040
rect 18601 18031 18659 18037
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 19889 18071 19947 18077
rect 19889 18037 19901 18071
rect 19935 18068 19947 18071
rect 19996 18068 20024 18167
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20237 18207 20295 18213
rect 20237 18204 20249 18207
rect 20128 18176 20249 18204
rect 20128 18164 20134 18176
rect 20237 18173 20249 18176
rect 20283 18204 20295 18207
rect 20283 18176 20944 18204
rect 20283 18173 20295 18176
rect 20237 18167 20295 18173
rect 20916 18148 20944 18176
rect 22370 18164 22376 18216
rect 22428 18204 22434 18216
rect 22465 18207 22523 18213
rect 22465 18204 22477 18207
rect 22428 18176 22477 18204
rect 22428 18164 22434 18176
rect 22465 18173 22477 18176
rect 22511 18173 22523 18207
rect 24026 18204 24032 18216
rect 23987 18176 24032 18204
rect 22465 18167 22523 18173
rect 24026 18164 24032 18176
rect 24084 18204 24090 18216
rect 25038 18204 25044 18216
rect 24084 18176 25044 18204
rect 24084 18164 24090 18176
rect 25038 18164 25044 18176
rect 25096 18164 25102 18216
rect 25225 18207 25283 18213
rect 25225 18173 25237 18207
rect 25271 18204 25283 18207
rect 25774 18204 25780 18216
rect 25271 18176 25780 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25774 18164 25780 18176
rect 25832 18164 25838 18216
rect 20898 18096 20904 18148
rect 20956 18096 20962 18148
rect 21542 18096 21548 18148
rect 21600 18096 21606 18148
rect 22094 18096 22100 18148
rect 22152 18136 22158 18148
rect 23014 18136 23020 18148
rect 22152 18108 23020 18136
rect 22152 18096 22158 18108
rect 23014 18096 23020 18108
rect 23072 18096 23078 18148
rect 24118 18096 24124 18148
rect 24176 18136 24182 18148
rect 24213 18139 24271 18145
rect 24213 18136 24225 18139
rect 24176 18108 24225 18136
rect 24176 18096 24182 18108
rect 24213 18105 24225 18108
rect 24259 18105 24271 18139
rect 24213 18099 24271 18105
rect 21560 18068 21588 18096
rect 22186 18068 22192 18080
rect 19935 18040 21588 18068
rect 22099 18040 22192 18068
rect 19935 18037 19947 18040
rect 19889 18031 19947 18037
rect 22186 18028 22192 18040
rect 22244 18068 22250 18080
rect 22281 18071 22339 18077
rect 22281 18068 22293 18071
rect 22244 18040 22293 18068
rect 22244 18028 22250 18040
rect 22281 18037 22293 18040
rect 22327 18037 22339 18071
rect 22281 18031 22339 18037
rect 23842 18028 23848 18080
rect 23900 18068 23906 18080
rect 24670 18068 24676 18080
rect 23900 18040 24676 18068
rect 23900 18028 23906 18040
rect 24670 18028 24676 18040
rect 24728 18028 24734 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1949 17867 2007 17873
rect 1949 17833 1961 17867
rect 1995 17864 2007 17867
rect 2682 17864 2688 17876
rect 1995 17836 2688 17864
rect 1995 17833 2007 17836
rect 1949 17827 2007 17833
rect 2682 17824 2688 17836
rect 2740 17824 2746 17876
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 3510 17864 3516 17876
rect 2832 17836 3516 17864
rect 2832 17824 2838 17836
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 3602 17824 3608 17876
rect 3660 17864 3666 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 3660 17836 3801 17864
rect 3660 17824 3666 17836
rect 3789 17833 3801 17836
rect 3835 17833 3847 17867
rect 6822 17864 6828 17876
rect 3789 17827 3847 17833
rect 4724 17836 6828 17864
rect 2317 17799 2375 17805
rect 2317 17765 2329 17799
rect 2363 17796 2375 17799
rect 2590 17796 2596 17808
rect 2363 17768 2596 17796
rect 2363 17765 2375 17768
rect 2317 17759 2375 17765
rect 2590 17756 2596 17768
rect 2648 17756 2654 17808
rect 2866 17756 2872 17808
rect 2924 17796 2930 17808
rect 2961 17799 3019 17805
rect 2961 17796 2973 17799
rect 2924 17768 2973 17796
rect 2924 17756 2930 17768
rect 2961 17765 2973 17768
rect 3007 17765 3019 17799
rect 2961 17759 3019 17765
rect 2682 17688 2688 17740
rect 2740 17728 2746 17740
rect 4724 17728 4752 17836
rect 6822 17824 6828 17836
rect 6880 17864 6886 17876
rect 6917 17867 6975 17873
rect 6917 17864 6929 17867
rect 6880 17836 6929 17864
rect 6880 17824 6886 17836
rect 6917 17833 6929 17836
rect 6963 17833 6975 17867
rect 6917 17827 6975 17833
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 7285 17867 7343 17873
rect 7285 17864 7297 17867
rect 7156 17836 7297 17864
rect 7156 17824 7162 17836
rect 7285 17833 7297 17836
rect 7331 17864 7343 17867
rect 7374 17864 7380 17876
rect 7331 17836 7380 17864
rect 7331 17833 7343 17836
rect 7285 17827 7343 17833
rect 7374 17824 7380 17836
rect 7432 17824 7438 17876
rect 8478 17864 8484 17876
rect 8439 17836 8484 17864
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 12529 17867 12587 17873
rect 8855 17836 12480 17864
rect 5166 17796 5172 17808
rect 2740 17700 4752 17728
rect 4816 17768 5172 17796
rect 2740 17688 2746 17700
rect 1394 17660 1400 17672
rect 1355 17632 1400 17660
rect 1394 17620 1400 17632
rect 1452 17620 1458 17672
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17660 3111 17663
rect 3602 17660 3608 17672
rect 3099 17632 3608 17660
rect 3099 17629 3111 17632
rect 3053 17623 3111 17629
rect 2976 17592 3004 17623
rect 3602 17620 3608 17632
rect 3660 17620 3666 17672
rect 4430 17620 4436 17672
rect 4488 17660 4494 17672
rect 4706 17660 4712 17672
rect 4488 17632 4712 17660
rect 4488 17620 4494 17632
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 4816 17660 4844 17768
rect 5166 17756 5172 17768
rect 5224 17796 5230 17808
rect 6178 17796 6184 17808
rect 5224 17768 6184 17796
rect 5224 17756 5230 17768
rect 6178 17756 6184 17768
rect 6236 17756 6242 17808
rect 8021 17799 8079 17805
rect 8021 17765 8033 17799
rect 8067 17796 8079 17799
rect 8297 17799 8355 17805
rect 8297 17796 8309 17799
rect 8067 17768 8309 17796
rect 8067 17765 8079 17768
rect 8021 17759 8079 17765
rect 8297 17765 8309 17768
rect 8343 17765 8355 17799
rect 8297 17759 8355 17765
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17728 4951 17731
rect 5252 17731 5310 17737
rect 5252 17728 5264 17731
rect 4939 17700 5264 17728
rect 4939 17697 4951 17700
rect 4893 17691 4951 17697
rect 5252 17697 5264 17700
rect 5298 17728 5310 17731
rect 5534 17728 5540 17740
rect 5298 17700 5540 17728
rect 5298 17697 5310 17700
rect 5252 17691 5310 17697
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 7006 17688 7012 17740
rect 7064 17688 7070 17740
rect 7558 17688 7564 17740
rect 7616 17728 7622 17740
rect 7742 17728 7748 17740
rect 7616 17700 7748 17728
rect 7616 17688 7622 17700
rect 7742 17688 7748 17700
rect 7800 17728 7806 17740
rect 8855 17728 8883 17836
rect 9493 17799 9551 17805
rect 9493 17765 9505 17799
rect 9539 17796 9551 17799
rect 10318 17796 10324 17808
rect 9539 17768 10324 17796
rect 9539 17765 9551 17768
rect 9493 17759 9551 17765
rect 10318 17756 10324 17768
rect 10376 17756 10382 17808
rect 11885 17799 11943 17805
rect 11885 17765 11897 17799
rect 11931 17796 11943 17799
rect 12066 17796 12072 17808
rect 11931 17768 12072 17796
rect 11931 17765 11943 17768
rect 11885 17759 11943 17765
rect 12066 17756 12072 17768
rect 12124 17756 12130 17808
rect 7800 17700 8883 17728
rect 7800 17688 7806 17700
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9858 17728 9864 17740
rect 9456 17700 9864 17728
rect 9456 17688 9462 17700
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 10134 17728 10140 17740
rect 10095 17700 10140 17728
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 11790 17728 11796 17740
rect 11532 17700 11796 17728
rect 4985 17663 5043 17669
rect 4985 17660 4997 17663
rect 4816 17632 4997 17660
rect 4985 17629 4997 17632
rect 5031 17629 5043 17663
rect 4985 17623 5043 17629
rect 3694 17592 3700 17604
rect 2976 17564 3700 17592
rect 3694 17552 3700 17564
rect 3752 17552 3758 17604
rect 5994 17552 6000 17604
rect 6052 17592 6058 17604
rect 7024 17592 7052 17688
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17629 7987 17663
rect 8110 17660 8116 17672
rect 8071 17632 8116 17660
rect 7929 17623 7987 17629
rect 7944 17592 7972 17623
rect 8110 17620 8116 17632
rect 8168 17620 8174 17672
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 9582 17660 9588 17672
rect 8996 17632 9588 17660
rect 8996 17620 9002 17632
rect 9582 17620 9588 17632
rect 9640 17660 9646 17672
rect 10413 17663 10471 17669
rect 9640 17632 9996 17660
rect 9640 17620 9646 17632
rect 8202 17592 8208 17604
rect 6052 17564 6500 17592
rect 7024 17564 7696 17592
rect 7944 17564 8208 17592
rect 6052 17552 6058 17564
rect 2130 17484 2136 17536
rect 2188 17524 2194 17536
rect 2501 17527 2559 17533
rect 2501 17524 2513 17527
rect 2188 17496 2513 17524
rect 2188 17484 2194 17496
rect 2501 17493 2513 17496
rect 2547 17493 2559 17527
rect 2501 17487 2559 17493
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 4706 17524 4712 17536
rect 4387 17496 4712 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 4706 17484 4712 17496
rect 4764 17524 4770 17536
rect 6178 17524 6184 17536
rect 4764 17496 6184 17524
rect 4764 17484 4770 17496
rect 6178 17484 6184 17496
rect 6236 17524 6242 17536
rect 6365 17527 6423 17533
rect 6365 17524 6377 17527
rect 6236 17496 6377 17524
rect 6236 17484 6242 17496
rect 6365 17493 6377 17496
rect 6411 17493 6423 17527
rect 6472 17524 6500 17564
rect 7668 17536 7696 17564
rect 8202 17552 8208 17564
rect 8260 17552 8266 17604
rect 8297 17595 8355 17601
rect 8297 17561 8309 17595
rect 8343 17592 8355 17595
rect 8343 17564 8984 17592
rect 8343 17561 8355 17564
rect 8297 17555 8355 17561
rect 7561 17527 7619 17533
rect 7561 17524 7573 17527
rect 6472 17496 7573 17524
rect 6365 17487 6423 17493
rect 7561 17493 7573 17496
rect 7607 17493 7619 17527
rect 7561 17487 7619 17493
rect 7650 17484 7656 17536
rect 7708 17484 7714 17536
rect 8956 17533 8984 17564
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 9861 17595 9919 17601
rect 9861 17592 9873 17595
rect 9732 17564 9873 17592
rect 9732 17552 9738 17564
rect 9861 17561 9873 17564
rect 9907 17561 9919 17595
rect 9861 17555 9919 17561
rect 8941 17527 8999 17533
rect 8941 17493 8953 17527
rect 8987 17524 8999 17527
rect 9582 17524 9588 17536
rect 8987 17496 9588 17524
rect 8987 17493 8999 17496
rect 8941 17487 8999 17493
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 9968 17524 9996 17632
rect 10413 17629 10425 17663
rect 10459 17660 10471 17663
rect 10686 17660 10692 17672
rect 10459 17632 10692 17660
rect 10459 17629 10471 17632
rect 10413 17623 10471 17629
rect 10686 17620 10692 17632
rect 10744 17620 10750 17672
rect 11054 17552 11060 17604
rect 11112 17592 11118 17604
rect 11425 17595 11483 17601
rect 11425 17592 11437 17595
rect 11112 17564 11437 17592
rect 11112 17552 11118 17564
rect 11425 17561 11437 17564
rect 11471 17561 11483 17595
rect 11425 17555 11483 17561
rect 10778 17524 10784 17536
rect 9968 17496 10784 17524
rect 10778 17484 10784 17496
rect 10836 17484 10842 17536
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11149 17527 11207 17533
rect 11149 17524 11161 17527
rect 11020 17496 11161 17524
rect 11020 17484 11026 17496
rect 11149 17493 11161 17496
rect 11195 17524 11207 17527
rect 11532 17524 11560 17700
rect 11790 17688 11796 17700
rect 11848 17728 11854 17740
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11848 17700 11989 17728
rect 11848 17688 11854 17700
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 12452 17728 12480 17836
rect 12529 17833 12541 17867
rect 12575 17864 12587 17867
rect 12894 17864 12900 17876
rect 12575 17836 12900 17864
rect 12575 17833 12587 17836
rect 12529 17827 12587 17833
rect 12894 17824 12900 17836
rect 12952 17864 12958 17876
rect 13354 17864 13360 17876
rect 12952 17836 13360 17864
rect 12952 17824 12958 17836
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 13449 17867 13507 17873
rect 13449 17833 13461 17867
rect 13495 17864 13507 17867
rect 13538 17864 13544 17876
rect 13495 17836 13544 17864
rect 13495 17833 13507 17836
rect 13449 17827 13507 17833
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 15102 17864 15108 17876
rect 15063 17836 15108 17864
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 15749 17867 15807 17873
rect 15749 17833 15761 17867
rect 15795 17864 15807 17867
rect 16022 17864 16028 17876
rect 15795 17836 16028 17864
rect 15795 17833 15807 17836
rect 15749 17827 15807 17833
rect 16022 17824 16028 17836
rect 16080 17824 16086 17876
rect 18046 17864 18052 17876
rect 18007 17836 18052 17864
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 18506 17824 18512 17876
rect 18564 17864 18570 17876
rect 18601 17867 18659 17873
rect 18601 17864 18613 17867
rect 18564 17836 18613 17864
rect 18564 17824 18570 17836
rect 18601 17833 18613 17836
rect 18647 17833 18659 17867
rect 18601 17827 18659 17833
rect 20717 17867 20775 17873
rect 20717 17833 20729 17867
rect 20763 17864 20775 17867
rect 20898 17864 20904 17876
rect 20763 17836 20904 17864
rect 20763 17833 20775 17836
rect 20717 17827 20775 17833
rect 20898 17824 20904 17836
rect 20956 17824 20962 17876
rect 21913 17867 21971 17873
rect 21913 17864 21925 17867
rect 21284 17836 21925 17864
rect 12802 17756 12808 17808
rect 12860 17796 12866 17808
rect 13262 17796 13268 17808
rect 12860 17768 13268 17796
rect 12860 17756 12866 17768
rect 13262 17756 13268 17768
rect 13320 17756 13326 17808
rect 16936 17799 16994 17805
rect 14200 17768 15608 17796
rect 14200 17728 14228 17768
rect 12452 17700 14228 17728
rect 11977 17691 12035 17697
rect 14274 17688 14280 17740
rect 14332 17688 14338 17740
rect 14550 17688 14556 17740
rect 14608 17688 14614 17740
rect 15580 17737 15608 17768
rect 16936 17765 16948 17799
rect 16982 17796 16994 17799
rect 17862 17796 17868 17808
rect 16982 17768 17868 17796
rect 16982 17765 16994 17768
rect 16936 17759 16994 17765
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 19794 17796 19800 17808
rect 19755 17768 19800 17796
rect 19794 17756 19800 17768
rect 19852 17756 19858 17808
rect 20806 17756 20812 17808
rect 20864 17796 20870 17808
rect 21284 17805 21312 17836
rect 21913 17833 21925 17836
rect 21959 17833 21971 17867
rect 22278 17864 22284 17876
rect 22239 17836 22284 17864
rect 21913 17827 21971 17833
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 23658 17864 23664 17876
rect 23619 17836 23664 17864
rect 23658 17824 23664 17836
rect 23716 17824 23722 17876
rect 23750 17824 23756 17876
rect 23808 17864 23814 17876
rect 24581 17867 24639 17873
rect 24581 17864 24593 17867
rect 23808 17836 24593 17864
rect 23808 17824 23814 17836
rect 24581 17833 24593 17836
rect 24627 17833 24639 17867
rect 24581 17827 24639 17833
rect 21269 17799 21327 17805
rect 21269 17796 21281 17799
rect 20864 17768 21281 17796
rect 20864 17756 20870 17768
rect 21269 17765 21281 17768
rect 21315 17765 21327 17799
rect 21269 17759 21327 17765
rect 21453 17799 21511 17805
rect 21453 17765 21465 17799
rect 21499 17765 21511 17799
rect 21453 17759 21511 17765
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17728 15623 17731
rect 16206 17728 16212 17740
rect 15611 17700 16212 17728
rect 15611 17697 15623 17700
rect 15565 17691 15623 17697
rect 16206 17688 16212 17700
rect 16264 17728 16270 17740
rect 16574 17728 16580 17740
rect 16264 17700 16580 17728
rect 16264 17688 16270 17700
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 16669 17731 16727 17737
rect 16669 17697 16681 17731
rect 16715 17728 16727 17731
rect 17218 17728 17224 17740
rect 16715 17700 17224 17728
rect 16715 17697 16727 17700
rect 16669 17691 16727 17697
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 19889 17731 19947 17737
rect 19889 17728 19901 17731
rect 19484 17700 19901 17728
rect 19484 17688 19490 17700
rect 19889 17697 19901 17700
rect 19935 17697 19947 17731
rect 19889 17691 19947 17697
rect 20438 17688 20444 17740
rect 20496 17728 20502 17740
rect 21468 17728 21496 17759
rect 21542 17756 21548 17808
rect 21600 17796 21606 17808
rect 22830 17796 22836 17808
rect 21600 17768 22836 17796
rect 21600 17756 21606 17768
rect 22830 17756 22836 17768
rect 22888 17756 22894 17808
rect 23017 17799 23075 17805
rect 23017 17765 23029 17799
rect 23063 17796 23075 17799
rect 23106 17796 23112 17808
rect 23063 17768 23112 17796
rect 23063 17765 23075 17768
rect 23017 17759 23075 17765
rect 23106 17756 23112 17768
rect 23164 17756 23170 17808
rect 24596 17796 24624 17827
rect 24854 17824 24860 17876
rect 24912 17864 24918 17876
rect 25041 17867 25099 17873
rect 25041 17864 25053 17867
rect 24912 17836 25053 17864
rect 24912 17824 24918 17836
rect 25041 17833 25053 17836
rect 25087 17833 25099 17867
rect 25041 17827 25099 17833
rect 25409 17799 25467 17805
rect 25409 17796 25421 17799
rect 24596 17768 25421 17796
rect 25409 17765 25421 17768
rect 25455 17765 25467 17799
rect 25409 17759 25467 17765
rect 24394 17728 24400 17740
rect 20496 17700 21496 17728
rect 24355 17700 24400 17728
rect 20496 17688 20502 17700
rect 24394 17688 24400 17700
rect 24452 17728 24458 17740
rect 24854 17728 24860 17740
rect 24452 17700 24860 17728
rect 24452 17688 24458 17700
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 25038 17688 25044 17740
rect 25096 17728 25102 17740
rect 25777 17731 25835 17737
rect 25777 17728 25789 17731
rect 25096 17700 25789 17728
rect 25096 17688 25102 17700
rect 25777 17697 25789 17700
rect 25823 17697 25835 17731
rect 25777 17691 25835 17697
rect 11885 17663 11943 17669
rect 11885 17629 11897 17663
rect 11931 17629 11943 17663
rect 11885 17623 11943 17629
rect 11900 17592 11928 17623
rect 13446 17620 13452 17672
rect 13504 17660 13510 17672
rect 13541 17663 13599 17669
rect 13541 17660 13553 17663
rect 13504 17632 13553 17660
rect 13504 17620 13510 17632
rect 13541 17629 13553 17632
rect 13587 17629 13599 17663
rect 13541 17623 13599 17629
rect 12158 17592 12164 17604
rect 11900 17564 12164 17592
rect 12158 17552 12164 17564
rect 12216 17552 12222 17604
rect 12986 17524 12992 17536
rect 11195 17496 11560 17524
rect 12899 17496 12992 17524
rect 11195 17493 11207 17496
rect 11149 17487 11207 17493
rect 12986 17484 12992 17496
rect 13044 17524 13050 17536
rect 13909 17527 13967 17533
rect 13909 17524 13921 17527
rect 13044 17496 13921 17524
rect 13044 17484 13050 17496
rect 13909 17493 13921 17496
rect 13955 17493 13967 17527
rect 13909 17487 13967 17493
rect 14182 17484 14188 17536
rect 14240 17524 14246 17536
rect 14292 17524 14320 17688
rect 14369 17595 14427 17601
rect 14369 17561 14381 17595
rect 14415 17592 14427 17595
rect 14568 17592 14596 17688
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 15712 17632 16252 17660
rect 15712 17620 15718 17632
rect 15930 17592 15936 17604
rect 14415 17564 15936 17592
rect 14415 17561 14427 17564
rect 14369 17555 14427 17561
rect 15930 17552 15936 17564
rect 15988 17552 15994 17604
rect 16224 17601 16252 17632
rect 18874 17620 18880 17672
rect 18932 17660 18938 17672
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 18932 17632 19717 17660
rect 18932 17620 18938 17632
rect 19705 17629 19717 17632
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 20898 17620 20904 17672
rect 20956 17660 20962 17672
rect 21174 17660 21180 17672
rect 20956 17632 21180 17660
rect 20956 17620 20962 17632
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 21542 17660 21548 17672
rect 21503 17632 21548 17660
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17629 23167 17663
rect 24670 17660 24676 17672
rect 24631 17632 24676 17660
rect 23109 17623 23167 17629
rect 16209 17595 16267 17601
rect 16209 17561 16221 17595
rect 16255 17592 16267 17595
rect 19061 17595 19119 17601
rect 16255 17564 16712 17592
rect 16255 17561 16267 17564
rect 16209 17555 16267 17561
rect 14642 17524 14648 17536
rect 14240 17496 14320 17524
rect 14603 17496 14648 17524
rect 14240 17484 14246 17496
rect 14642 17484 14648 17496
rect 14700 17484 14706 17536
rect 16574 17524 16580 17536
rect 16535 17496 16580 17524
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 16684 17524 16712 17564
rect 19061 17561 19073 17595
rect 19107 17592 19119 17595
rect 19610 17592 19616 17604
rect 19107 17564 19616 17592
rect 19107 17561 19119 17564
rect 19061 17555 19119 17561
rect 19610 17552 19616 17564
rect 19668 17552 19674 17604
rect 20349 17595 20407 17601
rect 20349 17561 20361 17595
rect 20395 17592 20407 17595
rect 21082 17592 21088 17604
rect 20395 17564 21088 17592
rect 20395 17561 20407 17564
rect 20349 17555 20407 17561
rect 21082 17552 21088 17564
rect 21140 17552 21146 17604
rect 21560 17592 21588 17620
rect 23124 17592 23152 17623
rect 24670 17620 24676 17632
rect 24728 17620 24734 17672
rect 24118 17592 24124 17604
rect 21560 17564 23152 17592
rect 24079 17564 24124 17592
rect 24118 17552 24124 17564
rect 24176 17552 24182 17604
rect 18966 17524 18972 17536
rect 16684 17496 18972 17524
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19337 17527 19395 17533
rect 19337 17493 19349 17527
rect 19383 17524 19395 17527
rect 20530 17524 20536 17536
rect 19383 17496 20536 17524
rect 19383 17493 19395 17496
rect 19337 17487 19395 17493
rect 20530 17484 20536 17496
rect 20588 17484 20594 17536
rect 20714 17484 20720 17536
rect 20772 17524 20778 17536
rect 20993 17527 21051 17533
rect 20993 17524 21005 17527
rect 20772 17496 21005 17524
rect 20772 17484 20778 17496
rect 20993 17493 21005 17496
rect 21039 17493 21051 17527
rect 22554 17524 22560 17536
rect 22515 17496 22560 17524
rect 20993 17487 21051 17493
rect 22554 17484 22560 17496
rect 22612 17484 22618 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2406 17280 2412 17332
rect 2464 17320 2470 17332
rect 3602 17320 3608 17332
rect 2464 17292 3608 17320
rect 2464 17280 2470 17292
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 4338 17320 4344 17332
rect 4299 17292 4344 17320
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 5261 17323 5319 17329
rect 5261 17320 5273 17323
rect 5224 17292 5273 17320
rect 5224 17280 5230 17292
rect 5261 17289 5273 17292
rect 5307 17289 5319 17323
rect 6914 17320 6920 17332
rect 6875 17292 6920 17320
rect 5261 17283 5319 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 7006 17280 7012 17332
rect 7064 17320 7070 17332
rect 7926 17320 7932 17332
rect 7064 17292 7932 17320
rect 7064 17280 7070 17292
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8938 17320 8944 17332
rect 8772 17292 8944 17320
rect 2777 17255 2835 17261
rect 2777 17221 2789 17255
rect 2823 17252 2835 17255
rect 3234 17252 3240 17264
rect 2823 17224 3240 17252
rect 2823 17221 2835 17224
rect 2777 17215 2835 17221
rect 3234 17212 3240 17224
rect 3292 17212 3298 17264
rect 4157 17255 4215 17261
rect 4157 17252 4169 17255
rect 3988 17224 4169 17252
rect 3878 17184 3884 17196
rect 1412 17156 3884 17184
rect 1412 17125 1440 17156
rect 3878 17144 3884 17156
rect 3936 17144 3942 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17085 1455 17119
rect 1397 17079 1455 17085
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 1762 17116 1768 17128
rect 1719 17088 1768 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 2501 17119 2559 17125
rect 2501 17085 2513 17119
rect 2547 17116 2559 17119
rect 2866 17116 2872 17128
rect 2547 17088 2872 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 2866 17076 2872 17088
rect 2924 17116 2930 17128
rect 3510 17116 3516 17128
rect 2924 17088 3516 17116
rect 2924 17076 2930 17088
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 2774 17008 2780 17060
rect 2832 17008 2838 17060
rect 3050 17048 3056 17060
rect 3011 17020 3056 17048
rect 3050 17008 3056 17020
rect 3108 17008 3114 17060
rect 3237 17051 3295 17057
rect 3237 17048 3249 17051
rect 3160 17020 3249 17048
rect 2792 16980 2820 17008
rect 3160 16980 3188 17020
rect 3237 17017 3249 17020
rect 3283 17017 3295 17051
rect 3237 17011 3295 17017
rect 3329 17051 3387 17057
rect 3329 17017 3341 17051
rect 3375 17048 3387 17051
rect 3602 17048 3608 17060
rect 3375 17020 3608 17048
rect 3375 17017 3387 17020
rect 3329 17011 3387 17017
rect 3602 17008 3608 17020
rect 3660 17048 3666 17060
rect 3988 17048 4016 17224
rect 4157 17221 4169 17224
rect 4203 17252 4215 17255
rect 5626 17252 5632 17264
rect 4203 17224 5632 17252
rect 4203 17221 4215 17224
rect 4157 17215 4215 17221
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 7190 17212 7196 17264
rect 7248 17252 7254 17264
rect 8573 17255 8631 17261
rect 8573 17252 8585 17255
rect 7248 17224 8585 17252
rect 7248 17212 7254 17224
rect 8573 17221 8585 17224
rect 8619 17252 8631 17255
rect 8772 17252 8800 17292
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 12526 17320 12532 17332
rect 12487 17292 12532 17320
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 13538 17320 13544 17332
rect 13499 17292 13544 17320
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 14093 17323 14151 17329
rect 14093 17289 14105 17323
rect 14139 17320 14151 17323
rect 14182 17320 14188 17332
rect 14139 17292 14188 17320
rect 14139 17289 14151 17292
rect 14093 17283 14151 17289
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 14366 17280 14372 17332
rect 14424 17320 14430 17332
rect 14826 17320 14832 17332
rect 14424 17292 14832 17320
rect 14424 17280 14430 17292
rect 14826 17280 14832 17292
rect 14884 17280 14890 17332
rect 16206 17320 16212 17332
rect 16167 17292 16212 17320
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 17037 17323 17095 17329
rect 17037 17289 17049 17323
rect 17083 17320 17095 17323
rect 17586 17320 17592 17332
rect 17083 17292 17592 17320
rect 17083 17289 17095 17292
rect 17037 17283 17095 17289
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 19794 17320 19800 17332
rect 17972 17292 19800 17320
rect 8619 17224 8800 17252
rect 8619 17221 8631 17224
rect 8573 17215 8631 17221
rect 4798 17184 4804 17196
rect 4759 17156 4804 17184
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 6273 17187 6331 17193
rect 6273 17184 6285 17187
rect 5500 17156 6285 17184
rect 5500 17144 5506 17156
rect 6273 17153 6285 17156
rect 6319 17184 6331 17187
rect 7466 17184 7472 17196
rect 6319 17156 7472 17184
rect 6319 17153 6331 17156
rect 6273 17147 6331 17153
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 8772 17193 8800 17224
rect 10137 17255 10195 17261
rect 10137 17221 10149 17255
rect 10183 17252 10195 17255
rect 10962 17252 10968 17264
rect 10183 17224 10968 17252
rect 10183 17221 10195 17224
rect 10137 17215 10195 17221
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 12158 17252 12164 17264
rect 12119 17224 12164 17252
rect 12158 17212 12164 17224
rect 12216 17212 12222 17264
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17153 8815 17187
rect 11330 17184 11336 17196
rect 11291 17156 11336 17184
rect 8757 17147 8815 17153
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 12066 17184 12072 17196
rect 12027 17156 12072 17184
rect 12066 17144 12072 17156
rect 12124 17144 12130 17196
rect 12710 17144 12716 17196
rect 12768 17144 12774 17196
rect 12989 17187 13047 17193
rect 12989 17153 13001 17187
rect 13035 17184 13047 17187
rect 13170 17184 13176 17196
rect 13035 17156 13176 17184
rect 13035 17153 13047 17156
rect 12989 17147 13047 17153
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 14200 17193 14228 17280
rect 15565 17255 15623 17261
rect 15565 17221 15577 17255
rect 15611 17252 15623 17255
rect 15930 17252 15936 17264
rect 15611 17224 15936 17252
rect 15611 17221 15623 17224
rect 15565 17215 15623 17221
rect 15930 17212 15936 17224
rect 15988 17212 15994 17264
rect 16761 17255 16819 17261
rect 16761 17221 16773 17255
rect 16807 17252 16819 17255
rect 17218 17252 17224 17264
rect 16807 17224 17224 17252
rect 16807 17221 16819 17224
rect 16761 17215 16819 17221
rect 17218 17212 17224 17224
rect 17276 17212 17282 17264
rect 17497 17255 17555 17261
rect 17497 17221 17509 17255
rect 17543 17252 17555 17255
rect 17862 17252 17868 17264
rect 17543 17224 17868 17252
rect 17543 17221 17555 17224
rect 17497 17215 17555 17221
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17153 14243 17187
rect 17972 17184 18000 17292
rect 19794 17280 19800 17292
rect 19852 17320 19858 17332
rect 19981 17323 20039 17329
rect 19981 17320 19993 17323
rect 19852 17292 19993 17320
rect 19852 17280 19858 17292
rect 19981 17289 19993 17292
rect 20027 17320 20039 17323
rect 20714 17320 20720 17332
rect 20027 17292 20720 17320
rect 20027 17289 20039 17292
rect 19981 17283 20039 17289
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 21266 17320 21272 17332
rect 20864 17292 21272 17320
rect 20864 17280 20870 17292
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 22554 17320 22560 17332
rect 22112 17292 22560 17320
rect 19061 17255 19119 17261
rect 19061 17221 19073 17255
rect 19107 17252 19119 17255
rect 19107 17224 20484 17252
rect 19107 17221 19119 17224
rect 19061 17215 19119 17221
rect 18782 17184 18788 17196
rect 14185 17147 14243 17153
rect 16500 17156 18000 17184
rect 18064 17156 18788 17184
rect 4706 17076 4712 17128
rect 4764 17116 4770 17128
rect 4893 17119 4951 17125
rect 4893 17116 4905 17119
rect 4764 17088 4905 17116
rect 4764 17076 4770 17088
rect 4893 17085 4905 17088
rect 4939 17085 4951 17119
rect 4893 17079 4951 17085
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 12728 17116 12756 17144
rect 16500 17116 16528 17156
rect 10008 17088 12756 17116
rect 14292 17088 16528 17116
rect 10008 17076 10014 17088
rect 4798 17048 4804 17060
rect 3660 17020 4016 17048
rect 4759 17020 4804 17048
rect 3660 17008 3666 17020
rect 4798 17008 4804 17020
rect 4856 17008 4862 17060
rect 6914 17008 6920 17060
rect 6972 17048 6978 17060
rect 7193 17051 7251 17057
rect 7193 17048 7205 17051
rect 6972 17020 7205 17048
rect 6972 17008 6978 17020
rect 7193 17017 7205 17020
rect 7239 17017 7251 17051
rect 7374 17048 7380 17060
rect 7335 17020 7380 17048
rect 7193 17011 7251 17017
rect 7374 17008 7380 17020
rect 7432 17008 7438 17060
rect 7929 17051 7987 17057
rect 7929 17017 7941 17051
rect 7975 17048 7987 17051
rect 8110 17048 8116 17060
rect 7975 17020 8116 17048
rect 7975 17017 7987 17020
rect 7929 17011 7987 17017
rect 8110 17008 8116 17020
rect 8168 17048 8174 17060
rect 8297 17051 8355 17057
rect 8297 17048 8309 17051
rect 8168 17020 8309 17048
rect 8168 17008 8174 17020
rect 8297 17017 8309 17020
rect 8343 17048 8355 17051
rect 9024 17051 9082 17057
rect 9024 17048 9036 17051
rect 8343 17020 9036 17048
rect 8343 17017 8355 17020
rect 8297 17011 8355 17017
rect 9024 17017 9036 17020
rect 9070 17048 9082 17051
rect 9122 17048 9128 17060
rect 9070 17020 9128 17048
rect 9070 17017 9082 17020
rect 9024 17011 9082 17017
rect 9122 17008 9128 17020
rect 9180 17008 9186 17060
rect 12342 17008 12348 17060
rect 12400 17048 12406 17060
rect 12434 17048 12440 17060
rect 12400 17020 12440 17048
rect 12400 17008 12406 17020
rect 12434 17008 12440 17020
rect 12492 17008 12498 17060
rect 12986 17048 12992 17060
rect 12947 17020 12992 17048
rect 12986 17008 12992 17020
rect 13044 17008 13050 17060
rect 13078 17008 13084 17060
rect 13136 17048 13142 17060
rect 13136 17020 13181 17048
rect 13136 17008 13142 17020
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 14292 17048 14320 17088
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 16724 17088 16865 17116
rect 16724 17076 16730 17088
rect 16853 17085 16865 17088
rect 16899 17085 16911 17119
rect 16853 17079 16911 17085
rect 17034 17076 17040 17128
rect 17092 17116 17098 17128
rect 18064 17116 18092 17156
rect 18782 17144 18788 17156
rect 18840 17144 18846 17196
rect 19518 17184 19524 17196
rect 19479 17156 19524 17184
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 20346 17184 20352 17196
rect 19668 17156 20352 17184
rect 19668 17144 19674 17156
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 19886 17116 19892 17128
rect 17092 17088 18092 17116
rect 18984 17088 19892 17116
rect 17092 17076 17098 17088
rect 13596 17020 14320 17048
rect 13596 17008 13602 17020
rect 14366 17008 14372 17060
rect 14424 17057 14430 17060
rect 14424 17051 14488 17057
rect 14424 17017 14442 17051
rect 14476 17017 14488 17051
rect 14424 17011 14488 17017
rect 14424 17008 14430 17011
rect 16942 17008 16948 17060
rect 17000 17048 17006 17060
rect 18984 17048 19012 17088
rect 19886 17076 19892 17088
rect 19944 17076 19950 17128
rect 17000 17020 19012 17048
rect 17000 17008 17006 17020
rect 3694 16980 3700 16992
rect 2792 16952 3188 16980
rect 3655 16952 3700 16980
rect 3694 16940 3700 16952
rect 3752 16940 3758 16992
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 4706 16980 4712 16992
rect 4304 16952 4712 16980
rect 4304 16940 4310 16952
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 5629 16983 5687 16989
rect 5629 16980 5641 16983
rect 5592 16952 5641 16980
rect 5592 16940 5598 16952
rect 5629 16949 5641 16952
rect 5675 16949 5687 16983
rect 5629 16943 5687 16949
rect 6641 16983 6699 16989
rect 6641 16949 6653 16983
rect 6687 16980 6699 16983
rect 7392 16980 7420 17008
rect 6687 16952 7420 16980
rect 10873 16983 10931 16989
rect 6687 16949 6699 16952
rect 6641 16943 6699 16949
rect 10873 16949 10885 16983
rect 10919 16980 10931 16983
rect 11054 16980 11060 16992
rect 10919 16952 11060 16980
rect 10919 16949 10931 16952
rect 10873 16943 10931 16949
rect 11054 16940 11060 16952
rect 11112 16980 11118 16992
rect 11149 16983 11207 16989
rect 11149 16980 11161 16983
rect 11112 16952 11161 16980
rect 11112 16940 11118 16952
rect 11149 16949 11161 16952
rect 11195 16949 11207 16983
rect 11149 16943 11207 16949
rect 11238 16940 11244 16992
rect 11296 16980 11302 16992
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11296 16952 11805 16980
rect 11296 16940 11302 16952
rect 11793 16949 11805 16952
rect 11839 16980 11851 16983
rect 12069 16983 12127 16989
rect 12069 16980 12081 16983
rect 11839 16952 12081 16980
rect 11839 16949 11851 16952
rect 11793 16943 11851 16949
rect 12069 16949 12081 16952
rect 12115 16949 12127 16983
rect 12069 16943 12127 16949
rect 14182 16940 14188 16992
rect 14240 16980 14246 16992
rect 17770 16980 17776 16992
rect 14240 16952 17776 16980
rect 14240 16940 14246 16952
rect 17770 16940 17776 16952
rect 17828 16940 17834 16992
rect 17865 16983 17923 16989
rect 17865 16949 17877 16983
rect 17911 16980 17923 16983
rect 18230 16980 18236 16992
rect 17911 16952 18236 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 18509 16983 18567 16989
rect 18509 16949 18521 16983
rect 18555 16980 18567 16983
rect 19242 16980 19248 16992
rect 18555 16952 19248 16980
rect 18555 16949 18567 16952
rect 18509 16943 18567 16949
rect 19242 16940 19248 16952
rect 19300 16980 19306 16992
rect 19521 16983 19579 16989
rect 19521 16980 19533 16983
rect 19300 16952 19533 16980
rect 19300 16940 19306 16952
rect 19521 16949 19533 16952
rect 19567 16949 19579 16983
rect 19521 16943 19579 16949
rect 19978 16940 19984 16992
rect 20036 16980 20042 16992
rect 20349 16983 20407 16989
rect 20349 16980 20361 16983
rect 20036 16952 20361 16980
rect 20036 16940 20042 16952
rect 20349 16949 20361 16952
rect 20395 16949 20407 16983
rect 20456 16980 20484 17224
rect 20530 17212 20536 17264
rect 20588 17252 20594 17264
rect 20625 17255 20683 17261
rect 20625 17252 20637 17255
rect 20588 17224 20637 17252
rect 20588 17212 20594 17224
rect 20625 17221 20637 17224
rect 20671 17221 20683 17255
rect 20625 17215 20683 17221
rect 20990 17212 20996 17264
rect 21048 17252 21054 17264
rect 22112 17252 22140 17292
rect 22554 17280 22560 17292
rect 22612 17280 22618 17332
rect 22830 17280 22836 17332
rect 22888 17320 22894 17332
rect 23017 17323 23075 17329
rect 23017 17320 23029 17323
rect 22888 17292 23029 17320
rect 22888 17280 22894 17292
rect 23017 17289 23029 17292
rect 23063 17289 23075 17323
rect 23750 17320 23756 17332
rect 23711 17292 23756 17320
rect 23017 17283 23075 17289
rect 23750 17280 23756 17292
rect 23808 17280 23814 17332
rect 25409 17323 25467 17329
rect 25409 17289 25421 17323
rect 25455 17320 25467 17323
rect 25682 17320 25688 17332
rect 25455 17292 25688 17320
rect 25455 17289 25467 17292
rect 25409 17283 25467 17289
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 21048 17224 22140 17252
rect 21048 17212 21054 17224
rect 22186 17212 22192 17264
rect 22244 17252 22250 17264
rect 24670 17252 24676 17264
rect 22244 17224 23612 17252
rect 24631 17224 24676 17252
rect 22244 17212 22250 17224
rect 21082 17184 21088 17196
rect 21043 17156 21088 17184
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 22370 17144 22376 17196
rect 22428 17184 22434 17196
rect 22465 17187 22523 17193
rect 22465 17184 22477 17187
rect 22428 17156 22477 17184
rect 22428 17144 22434 17156
rect 22465 17153 22477 17156
rect 22511 17153 22523 17187
rect 22465 17147 22523 17153
rect 21174 17116 21180 17128
rect 21135 17088 21180 17116
rect 21174 17076 21180 17088
rect 21232 17076 21238 17128
rect 21450 17076 21456 17128
rect 21508 17116 21514 17128
rect 22278 17116 22284 17128
rect 21508 17088 22284 17116
rect 21508 17076 21514 17088
rect 22278 17076 22284 17088
rect 22336 17076 22342 17128
rect 23584 17116 23612 17224
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 25314 17212 25320 17264
rect 25372 17252 25378 17264
rect 25866 17252 25872 17264
rect 25372 17224 25872 17252
rect 25372 17212 25378 17224
rect 25866 17212 25872 17224
rect 25924 17212 25930 17264
rect 23658 17144 23664 17196
rect 23716 17184 23722 17196
rect 24121 17187 24179 17193
rect 24121 17184 24133 17187
rect 23716 17156 24133 17184
rect 23716 17144 23722 17156
rect 24121 17153 24133 17156
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 23584 17088 25237 17116
rect 25225 17085 25237 17088
rect 25271 17116 25283 17119
rect 25777 17119 25835 17125
rect 25777 17116 25789 17119
rect 25271 17088 25789 17116
rect 25271 17085 25283 17088
rect 25225 17079 25283 17085
rect 25777 17085 25789 17088
rect 25823 17085 25835 17119
rect 25777 17079 25835 17085
rect 24305 17051 24363 17057
rect 24305 17048 24317 17051
rect 22112 17020 24317 17048
rect 20530 16980 20536 16992
rect 20456 16952 20536 16980
rect 20349 16943 20407 16949
rect 20530 16940 20536 16952
rect 20588 16980 20594 16992
rect 21085 16983 21143 16989
rect 21085 16980 21097 16983
rect 20588 16952 21097 16980
rect 20588 16940 20594 16952
rect 21085 16949 21097 16952
rect 21131 16949 21143 16983
rect 21542 16980 21548 16992
rect 21503 16952 21548 16980
rect 21085 16943 21143 16949
rect 21542 16940 21548 16952
rect 21600 16980 21606 16992
rect 22112 16989 22140 17020
rect 24305 17017 24317 17020
rect 24351 17048 24363 17051
rect 24670 17048 24676 17060
rect 24351 17020 24676 17048
rect 24351 17017 24363 17020
rect 24305 17011 24363 17017
rect 24670 17008 24676 17020
rect 24728 17048 24734 17060
rect 25041 17051 25099 17057
rect 25041 17048 25053 17051
rect 24728 17020 25053 17048
rect 24728 17008 24734 17020
rect 25041 17017 25053 17020
rect 25087 17017 25099 17051
rect 25041 17011 25099 17017
rect 22097 16983 22155 16989
rect 22097 16980 22109 16983
rect 21600 16952 22109 16980
rect 21600 16940 21606 16952
rect 22097 16949 22109 16952
rect 22143 16949 22155 16983
rect 22097 16943 22155 16949
rect 23014 16940 23020 16992
rect 23072 16980 23078 16992
rect 23477 16983 23535 16989
rect 23477 16980 23489 16983
rect 23072 16952 23489 16980
rect 23072 16940 23078 16952
rect 23477 16949 23489 16952
rect 23523 16980 23535 16983
rect 24210 16980 24216 16992
rect 23523 16952 24216 16980
rect 23523 16949 23535 16952
rect 23477 16943 23535 16949
rect 24210 16940 24216 16952
rect 24268 16940 24274 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2317 16779 2375 16785
rect 2317 16745 2329 16779
rect 2363 16776 2375 16779
rect 2406 16776 2412 16788
rect 2363 16748 2412 16776
rect 2363 16745 2375 16748
rect 2317 16739 2375 16745
rect 2406 16736 2412 16748
rect 2464 16736 2470 16788
rect 3050 16736 3056 16788
rect 3108 16776 3114 16788
rect 3418 16776 3424 16788
rect 3108 16748 3424 16776
rect 3108 16736 3114 16748
rect 3418 16736 3424 16748
rect 3476 16736 3482 16788
rect 3878 16776 3884 16788
rect 3791 16748 3884 16776
rect 3878 16736 3884 16748
rect 3936 16776 3942 16788
rect 5442 16776 5448 16788
rect 3936 16748 4292 16776
rect 5403 16748 5448 16776
rect 3936 16736 3942 16748
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 2961 16711 3019 16717
rect 2961 16708 2973 16711
rect 2648 16680 2973 16708
rect 2648 16668 2654 16680
rect 2961 16677 2973 16680
rect 3007 16708 3019 16711
rect 3970 16708 3976 16720
rect 3007 16680 3976 16708
rect 3007 16677 3019 16680
rect 2961 16671 3019 16677
rect 3970 16668 3976 16680
rect 4028 16668 4034 16720
rect 4264 16708 4292 16748
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 6914 16776 6920 16788
rect 6875 16748 6920 16776
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 8481 16779 8539 16785
rect 8481 16745 8493 16779
rect 8527 16745 8539 16779
rect 9858 16776 9864 16788
rect 9819 16748 9864 16776
rect 8481 16739 8539 16745
rect 5994 16708 6000 16720
rect 4264 16680 6000 16708
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 6178 16668 6184 16720
rect 6236 16708 6242 16720
rect 7346 16711 7404 16717
rect 7346 16708 7358 16711
rect 6236 16680 7358 16708
rect 6236 16668 6242 16680
rect 7346 16677 7358 16680
rect 7392 16677 7404 16711
rect 8496 16708 8524 16739
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 10686 16776 10692 16788
rect 10647 16748 10692 16776
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 12437 16779 12495 16785
rect 12437 16776 12449 16779
rect 11112 16748 12449 16776
rect 11112 16736 11118 16748
rect 12437 16745 12449 16748
rect 12483 16776 12495 16779
rect 13078 16776 13084 16788
rect 12483 16748 13084 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 13170 16736 13176 16788
rect 13228 16776 13234 16788
rect 13623 16779 13681 16785
rect 13623 16776 13635 16779
rect 13228 16748 13635 16776
rect 13228 16736 13234 16748
rect 13623 16745 13635 16748
rect 13669 16776 13681 16779
rect 14642 16776 14648 16788
rect 13669 16748 14648 16776
rect 13669 16745 13681 16748
rect 13623 16739 13681 16745
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 15010 16776 15016 16788
rect 14971 16748 15016 16776
rect 15010 16736 15016 16748
rect 15068 16776 15074 16788
rect 15838 16776 15844 16788
rect 15068 16748 15700 16776
rect 15799 16748 15844 16776
rect 15068 16736 15074 16748
rect 8846 16708 8852 16720
rect 8496 16680 8852 16708
rect 7346 16671 7404 16677
rect 8846 16668 8852 16680
rect 8904 16708 8910 16720
rect 8904 16680 10364 16708
rect 8904 16668 8910 16680
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 1762 16640 1768 16652
rect 1443 16612 1768 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 4338 16649 4344 16652
rect 2777 16643 2835 16649
rect 2777 16640 2789 16643
rect 2700 16612 2789 16640
rect 2498 16532 2504 16584
rect 2556 16572 2562 16584
rect 2700 16572 2728 16612
rect 2777 16609 2789 16612
rect 2823 16609 2835 16643
rect 2777 16603 2835 16609
rect 3053 16643 3111 16649
rect 3053 16609 3065 16643
rect 3099 16640 3111 16643
rect 4332 16640 4344 16649
rect 3099 16612 4344 16640
rect 3099 16609 3111 16612
rect 3053 16603 3111 16609
rect 4332 16603 4344 16612
rect 4338 16600 4344 16603
rect 4396 16600 4402 16652
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 6822 16640 6828 16652
rect 6595 16612 6828 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16640 7159 16643
rect 7190 16640 7196 16652
rect 7147 16612 7196 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 8202 16600 8208 16652
rect 8260 16640 8266 16652
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 8260 16612 9045 16640
rect 8260 16600 8266 16612
rect 9033 16609 9045 16612
rect 9079 16609 9091 16643
rect 9033 16603 9091 16609
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16640 9551 16643
rect 9677 16643 9735 16649
rect 9539 16612 9628 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 2556 16544 2728 16572
rect 4065 16575 4123 16581
rect 2556 16532 2562 16544
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 9600 16572 9628 16612
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 10226 16640 10232 16652
rect 9723 16612 10232 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 9858 16572 9864 16584
rect 9600 16544 9864 16572
rect 4065 16535 4123 16541
rect 2130 16464 2136 16516
rect 2188 16504 2194 16516
rect 2682 16504 2688 16516
rect 2188 16476 2688 16504
rect 2188 16464 2194 16476
rect 2682 16464 2688 16476
rect 2740 16464 2746 16516
rect 1946 16436 1952 16448
rect 1907 16408 1952 16436
rect 1946 16396 1952 16408
rect 2004 16396 2010 16448
rect 2501 16439 2559 16445
rect 2501 16405 2513 16439
rect 2547 16436 2559 16439
rect 2866 16436 2872 16448
rect 2547 16408 2872 16436
rect 2547 16405 2559 16408
rect 2501 16399 2559 16405
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 4080 16436 4108 16535
rect 9858 16532 9864 16544
rect 9916 16532 9922 16584
rect 4246 16436 4252 16448
rect 4080 16408 4252 16436
rect 4246 16396 4252 16408
rect 4304 16436 4310 16448
rect 5166 16436 5172 16448
rect 4304 16408 5172 16436
rect 4304 16396 4310 16408
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 5994 16436 6000 16448
rect 5955 16408 6000 16436
rect 5994 16396 6000 16408
rect 6052 16396 6058 16448
rect 10336 16445 10364 16680
rect 10962 16668 10968 16720
rect 11020 16708 11026 16720
rect 11302 16711 11360 16717
rect 11302 16708 11314 16711
rect 11020 16680 11314 16708
rect 11020 16668 11026 16680
rect 11302 16677 11314 16680
rect 11348 16708 11360 16711
rect 13446 16708 13452 16720
rect 11348 16680 13452 16708
rect 11348 16677 11360 16680
rect 11302 16671 11360 16677
rect 13446 16668 13452 16680
rect 13504 16668 13510 16720
rect 13814 16668 13820 16720
rect 13872 16708 13878 16720
rect 15672 16717 15700 16748
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 18414 16736 18420 16788
rect 18472 16776 18478 16788
rect 18877 16779 18935 16785
rect 18877 16776 18889 16779
rect 18472 16748 18889 16776
rect 18472 16736 18478 16748
rect 18877 16745 18889 16748
rect 18923 16745 18935 16779
rect 19426 16776 19432 16788
rect 19387 16748 19432 16776
rect 18877 16739 18935 16745
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 20530 16776 20536 16788
rect 20491 16748 20536 16776
rect 20530 16736 20536 16748
rect 20588 16736 20594 16788
rect 21174 16776 21180 16788
rect 20916 16748 21180 16776
rect 14093 16711 14151 16717
rect 14093 16708 14105 16711
rect 13872 16680 14105 16708
rect 13872 16668 13878 16680
rect 14093 16677 14105 16680
rect 14139 16677 14151 16711
rect 14093 16671 14151 16677
rect 15657 16711 15715 16717
rect 15657 16677 15669 16711
rect 15703 16677 15715 16711
rect 15657 16671 15715 16677
rect 17218 16668 17224 16720
rect 17276 16708 17282 16720
rect 17764 16711 17822 16717
rect 17764 16708 17776 16711
rect 17276 16680 17776 16708
rect 17276 16668 17282 16680
rect 17764 16677 17776 16680
rect 17810 16708 17822 16711
rect 18046 16708 18052 16720
rect 17810 16680 18052 16708
rect 17810 16677 17822 16680
rect 17764 16671 17822 16677
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 20257 16711 20315 16717
rect 20257 16677 20269 16711
rect 20303 16708 20315 16711
rect 20438 16708 20444 16720
rect 20303 16680 20444 16708
rect 20303 16677 20315 16680
rect 20257 16671 20315 16677
rect 20438 16668 20444 16680
rect 20496 16668 20502 16720
rect 12710 16600 12716 16652
rect 12768 16640 12774 16652
rect 12989 16643 13047 16649
rect 12989 16640 13001 16643
rect 12768 16612 13001 16640
rect 12768 16600 12774 16612
rect 12989 16609 13001 16612
rect 13035 16609 13047 16643
rect 13464 16640 13492 16668
rect 14185 16643 14243 16649
rect 14185 16640 14197 16643
rect 13464 16612 14197 16640
rect 12989 16603 13047 16609
rect 14185 16609 14197 16612
rect 14231 16609 14243 16643
rect 14918 16640 14924 16652
rect 14185 16603 14243 16609
rect 14292 16612 14924 16640
rect 10778 16532 10784 16584
rect 10836 16572 10842 16584
rect 11057 16575 11115 16581
rect 11057 16572 11069 16575
rect 10836 16544 11069 16572
rect 10836 16532 10842 16544
rect 11057 16541 11069 16544
rect 11103 16541 11115 16575
rect 11057 16535 11115 16541
rect 10321 16439 10379 16445
rect 10321 16405 10333 16439
rect 10367 16436 10379 16439
rect 10870 16436 10876 16448
rect 10367 16408 10876 16436
rect 10367 16405 10379 16408
rect 10321 16399 10379 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11072 16436 11100 16535
rect 13078 16532 13084 16584
rect 13136 16572 13142 16584
rect 13630 16572 13636 16584
rect 13136 16544 13636 16572
rect 13136 16532 13142 16544
rect 13630 16532 13636 16544
rect 13688 16572 13694 16584
rect 14001 16575 14059 16581
rect 14001 16572 14013 16575
rect 13688 16544 14013 16572
rect 13688 16532 13694 16544
rect 14001 16541 14013 16544
rect 14047 16572 14059 16575
rect 14292 16572 14320 16612
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 15396 16612 16313 16640
rect 14047 16544 14320 16572
rect 14047 16541 14059 16544
rect 14001 16535 14059 16541
rect 14090 16464 14096 16516
rect 14148 16504 14154 16516
rect 15396 16513 15424 16612
rect 16301 16609 16313 16612
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 16482 16600 16488 16652
rect 16540 16640 16546 16652
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 16540 16612 16681 16640
rect 16540 16600 16546 16612
rect 16669 16609 16681 16612
rect 16715 16609 16727 16643
rect 16669 16603 16727 16609
rect 17310 16600 17316 16652
rect 17368 16640 17374 16652
rect 17497 16643 17555 16649
rect 17497 16640 17509 16643
rect 17368 16612 17509 16640
rect 17368 16600 17374 16612
rect 17497 16609 17509 16612
rect 17543 16640 17555 16643
rect 18322 16640 18328 16652
rect 17543 16612 18328 16640
rect 17543 16609 17555 16612
rect 17497 16603 17555 16609
rect 18322 16600 18328 16612
rect 18380 16600 18386 16652
rect 19978 16600 19984 16652
rect 20036 16640 20042 16652
rect 20916 16640 20944 16748
rect 21174 16736 21180 16748
rect 21232 16776 21238 16788
rect 22002 16776 22008 16788
rect 21232 16748 22008 16776
rect 21232 16736 21238 16748
rect 22002 16736 22008 16748
rect 22060 16736 22066 16788
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 22833 16779 22891 16785
rect 22833 16776 22845 16779
rect 22336 16748 22845 16776
rect 22336 16736 22342 16748
rect 22833 16745 22845 16748
rect 22879 16745 22891 16779
rect 23934 16776 23940 16788
rect 23895 16748 23940 16776
rect 22833 16739 22891 16745
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 24854 16776 24860 16788
rect 24815 16748 24860 16776
rect 24854 16736 24860 16748
rect 24912 16736 24918 16788
rect 25130 16776 25136 16788
rect 25091 16748 25136 16776
rect 25130 16736 25136 16748
rect 25188 16736 25194 16788
rect 20990 16668 20996 16720
rect 21048 16708 21054 16720
rect 21542 16708 21548 16720
rect 21048 16680 21548 16708
rect 21048 16668 21054 16680
rect 21542 16668 21548 16680
rect 21600 16668 21606 16720
rect 22370 16668 22376 16720
rect 22428 16708 22434 16720
rect 23382 16708 23388 16720
rect 22428 16680 23388 16708
rect 22428 16668 22434 16680
rect 23382 16668 23388 16680
rect 23440 16668 23446 16720
rect 21174 16649 21180 16652
rect 21168 16640 21180 16649
rect 20036 16612 20944 16640
rect 21135 16612 21180 16640
rect 20036 16600 20042 16612
rect 21168 16603 21180 16612
rect 21174 16600 21180 16603
rect 21232 16600 21238 16652
rect 22554 16600 22560 16652
rect 22612 16640 22618 16652
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 22612 16612 23765 16640
rect 22612 16600 22618 16612
rect 23753 16609 23765 16612
rect 23799 16640 23811 16643
rect 24946 16640 24952 16652
rect 23799 16612 24952 16640
rect 23799 16609 23811 16612
rect 23753 16603 23811 16609
rect 24946 16600 24952 16612
rect 25004 16600 25010 16652
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16572 15991 16575
rect 16390 16572 16396 16584
rect 15979 16544 16396 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 20438 16532 20444 16584
rect 20496 16572 20502 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20496 16544 20913 16572
rect 20496 16532 20502 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 22830 16532 22836 16584
rect 22888 16572 22894 16584
rect 23290 16572 23296 16584
rect 22888 16544 23296 16572
rect 22888 16532 22894 16544
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 24029 16575 24087 16581
rect 24029 16541 24041 16575
rect 24075 16541 24087 16575
rect 24029 16535 24087 16541
rect 15381 16507 15439 16513
rect 15381 16504 15393 16507
rect 14148 16476 15393 16504
rect 14148 16464 14154 16476
rect 15381 16473 15393 16476
rect 15427 16473 15439 16507
rect 15381 16467 15439 16473
rect 15654 16464 15660 16516
rect 15712 16504 15718 16516
rect 17037 16507 17095 16513
rect 17037 16504 17049 16507
rect 15712 16476 17049 16504
rect 15712 16464 15718 16476
rect 17037 16473 17049 16476
rect 17083 16473 17095 16507
rect 17037 16467 17095 16473
rect 19518 16464 19524 16516
rect 19576 16504 19582 16516
rect 19889 16507 19947 16513
rect 19889 16504 19901 16507
rect 19576 16476 19901 16504
rect 19576 16464 19582 16476
rect 19889 16473 19901 16476
rect 19935 16504 19947 16507
rect 20530 16504 20536 16516
rect 19935 16476 20536 16504
rect 19935 16473 19947 16476
rect 19889 16467 19947 16473
rect 20530 16464 20536 16476
rect 20588 16464 20594 16516
rect 24044 16504 24072 16535
rect 24210 16504 24216 16516
rect 23216 16476 24216 16504
rect 23216 16448 23244 16476
rect 24210 16464 24216 16476
rect 24268 16504 24274 16516
rect 24397 16507 24455 16513
rect 24397 16504 24409 16507
rect 24268 16476 24409 16504
rect 24268 16464 24274 16476
rect 24397 16473 24409 16476
rect 24443 16473 24455 16507
rect 24397 16467 24455 16473
rect 11422 16436 11428 16448
rect 11072 16408 11428 16436
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 14366 16396 14372 16448
rect 14424 16436 14430 16448
rect 14645 16439 14703 16445
rect 14645 16436 14657 16439
rect 14424 16408 14657 16436
rect 14424 16396 14430 16408
rect 14645 16405 14657 16408
rect 14691 16436 14703 16439
rect 16022 16436 16028 16448
rect 14691 16408 16028 16436
rect 14691 16405 14703 16408
rect 14645 16399 14703 16405
rect 16022 16396 16028 16408
rect 16080 16396 16086 16448
rect 21174 16396 21180 16448
rect 21232 16436 21238 16448
rect 22281 16439 22339 16445
rect 22281 16436 22293 16439
rect 21232 16408 22293 16436
rect 21232 16396 21238 16408
rect 22281 16405 22293 16408
rect 22327 16405 22339 16439
rect 23198 16436 23204 16448
rect 23159 16408 23204 16436
rect 22281 16399 22339 16405
rect 23198 16396 23204 16408
rect 23256 16396 23262 16448
rect 23290 16396 23296 16448
rect 23348 16436 23354 16448
rect 23477 16439 23535 16445
rect 23477 16436 23489 16439
rect 23348 16408 23489 16436
rect 23348 16396 23354 16408
rect 23477 16405 23489 16408
rect 23523 16405 23535 16439
rect 23477 16399 23535 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1581 16235 1639 16241
rect 1581 16201 1593 16235
rect 1627 16232 1639 16235
rect 1670 16232 1676 16244
rect 1627 16204 1676 16232
rect 1627 16201 1639 16204
rect 1581 16195 1639 16201
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 2498 16232 2504 16244
rect 2459 16204 2504 16232
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 4525 16235 4583 16241
rect 4525 16232 4537 16235
rect 4304 16204 4537 16232
rect 4304 16192 4310 16204
rect 4525 16201 4537 16204
rect 4571 16201 4583 16235
rect 4525 16195 4583 16201
rect 4798 16192 4804 16244
rect 4856 16232 4862 16244
rect 5169 16235 5227 16241
rect 5169 16232 5181 16235
rect 4856 16204 5181 16232
rect 4856 16192 4862 16204
rect 5169 16201 5181 16204
rect 5215 16201 5227 16235
rect 5169 16195 5227 16201
rect 6178 16192 6184 16244
rect 6236 16232 6242 16244
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6236 16204 6561 16232
rect 6236 16192 6242 16204
rect 6549 16201 6561 16204
rect 6595 16201 6607 16235
rect 9122 16232 9128 16244
rect 9083 16204 9128 16232
rect 6549 16195 6607 16201
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 12158 16232 12164 16244
rect 12119 16204 12164 16232
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 13078 16192 13084 16244
rect 13136 16232 13142 16244
rect 13541 16235 13599 16241
rect 13541 16232 13553 16235
rect 13136 16204 13553 16232
rect 13136 16192 13142 16204
rect 13541 16201 13553 16204
rect 13587 16201 13599 16235
rect 13541 16195 13599 16201
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 13909 16235 13967 16241
rect 13909 16232 13921 16235
rect 13872 16204 13921 16232
rect 13872 16192 13878 16204
rect 13909 16201 13921 16204
rect 13955 16232 13967 16235
rect 14182 16232 14188 16244
rect 13955 16204 14188 16232
rect 13955 16201 13967 16204
rect 13909 16195 13967 16201
rect 14182 16192 14188 16204
rect 14240 16192 14246 16244
rect 14366 16192 14372 16244
rect 14424 16232 14430 16244
rect 16022 16232 16028 16244
rect 14424 16204 15884 16232
rect 15983 16204 16028 16232
rect 14424 16192 14430 16204
rect 2133 16167 2191 16173
rect 2133 16133 2145 16167
rect 2179 16164 2191 16167
rect 2590 16164 2596 16176
rect 2179 16136 2596 16164
rect 2179 16133 2191 16136
rect 2133 16127 2191 16133
rect 2590 16124 2596 16136
rect 2648 16124 2654 16176
rect 8754 16124 8760 16176
rect 8812 16164 8818 16176
rect 10321 16167 10379 16173
rect 10321 16164 10333 16167
rect 8812 16136 10333 16164
rect 8812 16124 8818 16136
rect 10321 16133 10333 16136
rect 10367 16133 10379 16167
rect 12526 16164 12532 16176
rect 12487 16136 12532 16164
rect 10321 16127 10379 16133
rect 12526 16124 12532 16136
rect 12584 16124 12590 16176
rect 15856 16164 15884 16204
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 17218 16232 17224 16244
rect 17179 16204 17224 16232
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17368 16204 17509 16232
rect 17368 16192 17374 16204
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 19150 16232 19156 16244
rect 17497 16195 17555 16201
rect 18309 16204 19156 16232
rect 18309 16164 18337 16204
rect 19150 16192 19156 16204
rect 19208 16232 19214 16244
rect 19208 16204 22048 16232
rect 19208 16192 19214 16204
rect 15856 16136 18337 16164
rect 4798 16056 4804 16108
rect 4856 16096 4862 16108
rect 4982 16096 4988 16108
rect 4856 16068 4988 16096
rect 4856 16056 4862 16068
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5592 16068 5733 16096
rect 5592 16056 5598 16068
rect 5721 16065 5733 16068
rect 5767 16096 5779 16099
rect 6089 16099 6147 16105
rect 6089 16096 6101 16099
rect 5767 16068 6101 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 6089 16065 6101 16068
rect 6135 16065 6147 16099
rect 6089 16059 6147 16065
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 10870 16096 10876 16108
rect 9824 16068 10640 16096
rect 10831 16068 10876 16096
rect 9824 16056 9830 16068
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 16028 1458 16040
rect 1578 16028 1584 16040
rect 1452 16000 1584 16028
rect 1452 15988 1458 16000
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 2590 16028 2596 16040
rect 2503 16000 2596 16028
rect 2590 15988 2596 16000
rect 2648 16028 2654 16040
rect 4154 16028 4160 16040
rect 2648 16000 4160 16028
rect 2648 15988 2654 16000
rect 4154 15988 4160 16000
rect 4212 15988 4218 16040
rect 4614 15988 4620 16040
rect 4672 16028 4678 16040
rect 5445 16031 5503 16037
rect 5445 16028 5457 16031
rect 4672 16000 5457 16028
rect 4672 15988 4678 16000
rect 5445 15997 5457 16000
rect 5491 15997 5503 16031
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 5445 15991 5503 15997
rect 7576 16000 7757 16028
rect 1946 15920 1952 15972
rect 2004 15960 2010 15972
rect 2838 15963 2896 15969
rect 2838 15960 2850 15963
rect 2004 15932 2850 15960
rect 2004 15920 2010 15932
rect 2838 15929 2850 15932
rect 2884 15929 2896 15963
rect 4338 15960 4344 15972
rect 2838 15923 2896 15929
rect 3988 15932 4344 15960
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 3988 15901 4016 15932
rect 4338 15920 4344 15932
rect 4396 15960 4402 15972
rect 4396 15932 5028 15960
rect 4396 15920 4402 15932
rect 5000 15904 5028 15932
rect 5534 15920 5540 15972
rect 5592 15960 5598 15972
rect 5629 15963 5687 15969
rect 5629 15960 5641 15963
rect 5592 15932 5641 15960
rect 5592 15920 5598 15932
rect 5629 15929 5641 15932
rect 5675 15960 5687 15963
rect 6086 15960 6092 15972
rect 5675 15932 6092 15960
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 6086 15920 6092 15932
rect 6144 15920 6150 15972
rect 3973 15895 4031 15901
rect 3973 15892 3985 15895
rect 3936 15864 3985 15892
rect 3936 15852 3942 15864
rect 3973 15861 3985 15864
rect 4019 15861 4031 15895
rect 4982 15892 4988 15904
rect 4943 15864 4988 15892
rect 3973 15855 4031 15861
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 7190 15892 7196 15904
rect 7151 15864 7196 15892
rect 7190 15852 7196 15864
rect 7248 15892 7254 15904
rect 7576 15901 7604 16000
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 8570 15988 8576 16040
rect 8628 16028 8634 16040
rect 9122 16028 9128 16040
rect 8628 16000 9128 16028
rect 8628 15988 8634 16000
rect 9122 15988 9128 16000
rect 9180 15988 9186 16040
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 16028 10195 16031
rect 10318 16028 10324 16040
rect 10183 16000 10324 16028
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 10318 15988 10324 16000
rect 10376 16028 10382 16040
rect 10612 16037 10640 16068
rect 10870 16056 10876 16068
rect 10928 16056 10934 16108
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16096 13139 16099
rect 13446 16096 13452 16108
rect 13127 16068 13452 16096
rect 13127 16065 13139 16068
rect 13081 16059 13139 16065
rect 13446 16056 13452 16068
rect 13504 16056 13510 16108
rect 13740 16068 14780 16096
rect 10597 16031 10655 16037
rect 10376 16000 10548 16028
rect 10376 15988 10382 16000
rect 7650 15920 7656 15972
rect 7708 15960 7714 15972
rect 7990 15963 8048 15969
rect 7990 15960 8002 15963
rect 7708 15932 8002 15960
rect 7708 15920 7714 15932
rect 7990 15929 8002 15932
rect 8036 15929 8048 15963
rect 7990 15923 8048 15929
rect 10226 15920 10232 15972
rect 10284 15920 10290 15972
rect 10520 15960 10548 16000
rect 10597 15997 10609 16031
rect 10643 16028 10655 16031
rect 10686 16028 10692 16040
rect 10643 16000 10692 16028
rect 10643 15997 10655 16000
rect 10597 15991 10655 15997
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 11882 15960 11888 15972
rect 10520 15932 10824 15960
rect 11795 15932 11888 15960
rect 7561 15895 7619 15901
rect 7561 15892 7573 15895
rect 7248 15864 7573 15892
rect 7248 15852 7254 15864
rect 7561 15861 7573 15864
rect 7607 15861 7619 15895
rect 7561 15855 7619 15861
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 9677 15895 9735 15901
rect 9677 15892 9689 15895
rect 9640 15864 9689 15892
rect 9640 15852 9646 15864
rect 9677 15861 9689 15864
rect 9723 15892 9735 15895
rect 10244 15892 10272 15920
rect 10796 15901 10824 15932
rect 9723 15864 10272 15892
rect 10781 15895 10839 15901
rect 9723 15861 9735 15864
rect 9677 15855 9735 15861
rect 10781 15861 10793 15895
rect 10827 15892 10839 15895
rect 10870 15892 10876 15904
rect 10827 15864 10876 15892
rect 10827 15861 10839 15864
rect 10781 15855 10839 15861
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 11333 15895 11391 15901
rect 11333 15861 11345 15895
rect 11379 15892 11391 15895
rect 11422 15892 11428 15904
rect 11379 15864 11428 15892
rect 11379 15861 11391 15864
rect 11333 15855 11391 15861
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 11808 15901 11836 15932
rect 11882 15920 11888 15932
rect 11940 15960 11946 15972
rect 12805 15963 12863 15969
rect 12805 15960 12817 15963
rect 11940 15932 12817 15960
rect 11940 15920 11946 15932
rect 12805 15929 12817 15932
rect 12851 15929 12863 15963
rect 12805 15923 12863 15929
rect 11793 15895 11851 15901
rect 11793 15892 11805 15895
rect 11756 15864 11805 15892
rect 11756 15852 11762 15864
rect 11793 15861 11805 15864
rect 11839 15861 11851 15895
rect 11793 15855 11851 15861
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 12989 15895 13047 15901
rect 12989 15892 13001 15895
rect 12216 15864 13001 15892
rect 12216 15852 12222 15864
rect 12989 15861 13001 15864
rect 13035 15892 13047 15895
rect 13740 15892 13768 16068
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 16028 14611 16031
rect 14642 16028 14648 16040
rect 14599 16000 14648 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 14752 16028 14780 16068
rect 15378 16028 15384 16040
rect 14752 16000 15384 16028
rect 15378 15988 15384 16000
rect 15436 15988 15442 16040
rect 18322 16028 18328 16040
rect 18235 16000 18328 16028
rect 18322 15988 18328 16000
rect 18380 16028 18386 16040
rect 21174 16037 21180 16040
rect 18417 16031 18475 16037
rect 18417 16028 18429 16031
rect 18380 16000 18429 16028
rect 18380 15988 18386 16000
rect 18417 15997 18429 16000
rect 18463 16028 18475 16031
rect 20901 16031 20959 16037
rect 18463 16000 20484 16028
rect 18463 15997 18475 16000
rect 18417 15991 18475 15997
rect 18800 15972 18828 16000
rect 20456 15972 20484 16000
rect 20901 15997 20913 16031
rect 20947 16028 20959 16031
rect 21168 16028 21180 16037
rect 20947 16000 20981 16028
rect 21135 16000 21180 16028
rect 20947 15997 20959 16000
rect 20901 15991 20959 15997
rect 21168 15991 21180 16000
rect 14918 15969 14924 15972
rect 14912 15960 14924 15969
rect 14879 15932 14924 15960
rect 14912 15923 14924 15932
rect 14918 15920 14924 15923
rect 14976 15920 14982 15972
rect 18662 15963 18720 15969
rect 18662 15960 18674 15963
rect 18432 15932 18674 15960
rect 18432 15904 18460 15932
rect 18662 15929 18674 15932
rect 18708 15929 18720 15963
rect 18662 15923 18720 15929
rect 18782 15920 18788 15972
rect 18840 15920 18846 15972
rect 19242 15920 19248 15972
rect 19300 15960 19306 15972
rect 20438 15960 20444 15972
rect 19300 15932 19932 15960
rect 20351 15932 20444 15960
rect 19300 15920 19306 15932
rect 13035 15864 13768 15892
rect 13035 15861 13047 15864
rect 12989 15855 13047 15861
rect 15194 15852 15200 15904
rect 15252 15892 15258 15904
rect 15654 15892 15660 15904
rect 15252 15864 15660 15892
rect 15252 15852 15258 15864
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 16577 15895 16635 15901
rect 16577 15892 16589 15895
rect 16448 15864 16589 15892
rect 16448 15852 16454 15864
rect 16577 15861 16589 15864
rect 16623 15861 16635 15895
rect 16577 15855 16635 15861
rect 18414 15852 18420 15904
rect 18472 15852 18478 15904
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 19797 15895 19855 15901
rect 19797 15892 19809 15895
rect 19392 15864 19809 15892
rect 19392 15852 19398 15864
rect 19797 15861 19809 15864
rect 19843 15861 19855 15895
rect 19904 15892 19932 15932
rect 20438 15920 20444 15932
rect 20496 15960 20502 15972
rect 20809 15963 20867 15969
rect 20809 15960 20821 15963
rect 20496 15932 20821 15960
rect 20496 15920 20502 15932
rect 20809 15929 20821 15932
rect 20855 15960 20867 15963
rect 20916 15960 20944 15991
rect 21174 15988 21180 15991
rect 21232 15988 21238 16040
rect 22020 16028 22048 16204
rect 22094 16192 22100 16244
rect 22152 16232 22158 16244
rect 22281 16235 22339 16241
rect 22281 16232 22293 16235
rect 22152 16204 22293 16232
rect 22152 16192 22158 16204
rect 22281 16201 22293 16204
rect 22327 16201 22339 16235
rect 22281 16195 22339 16201
rect 22554 16192 22560 16244
rect 22612 16232 22618 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 22612 16204 23029 16232
rect 22612 16192 22618 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 23474 16232 23480 16244
rect 23435 16204 23480 16232
rect 23017 16195 23075 16201
rect 23474 16192 23480 16204
rect 23532 16192 23538 16244
rect 24946 16232 24952 16244
rect 24907 16204 24952 16232
rect 24946 16192 24952 16204
rect 25004 16192 25010 16244
rect 25409 16235 25467 16241
rect 25409 16201 25421 16235
rect 25455 16232 25467 16235
rect 25498 16232 25504 16244
rect 25455 16204 25504 16232
rect 25455 16201 25467 16204
rect 25409 16195 25467 16201
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 23382 16124 23388 16176
rect 23440 16164 23446 16176
rect 23753 16167 23811 16173
rect 23753 16164 23765 16167
rect 23440 16136 23765 16164
rect 23440 16124 23446 16136
rect 23753 16133 23765 16136
rect 23799 16133 23811 16167
rect 24394 16164 24400 16176
rect 23753 16127 23811 16133
rect 24136 16136 24400 16164
rect 24136 16105 24164 16136
rect 24394 16124 24400 16136
rect 24452 16164 24458 16176
rect 25222 16164 25228 16176
rect 24452 16136 25228 16164
rect 24452 16124 24458 16136
rect 25222 16124 25228 16136
rect 25280 16124 25286 16176
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 24210 16056 24216 16108
rect 24268 16096 24274 16108
rect 24305 16099 24363 16105
rect 24305 16096 24317 16099
rect 24268 16068 24317 16096
rect 24268 16056 24274 16068
rect 24305 16065 24317 16068
rect 24351 16065 24363 16099
rect 24305 16059 24363 16065
rect 24946 16028 24952 16040
rect 22020 16000 24952 16028
rect 24946 15988 24952 16000
rect 25004 15988 25010 16040
rect 25225 16031 25283 16037
rect 25225 15997 25237 16031
rect 25271 16028 25283 16031
rect 25777 16031 25835 16037
rect 25777 16028 25789 16031
rect 25271 16000 25789 16028
rect 25271 15997 25283 16000
rect 25225 15991 25283 15997
rect 25777 15997 25789 16000
rect 25823 16028 25835 16031
rect 26142 16028 26148 16040
rect 25823 16000 26148 16028
rect 25823 15997 25835 16000
rect 25777 15991 25835 15997
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 21450 15960 21456 15972
rect 20855 15932 21456 15960
rect 20855 15929 20867 15932
rect 20809 15923 20867 15929
rect 21450 15920 21456 15932
rect 21508 15920 21514 15972
rect 23566 15960 23572 15972
rect 21744 15932 23572 15960
rect 21744 15892 21772 15932
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 19904 15864 21772 15892
rect 19797 15855 19855 15861
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 23014 15892 23020 15904
rect 22152 15864 23020 15892
rect 22152 15852 22158 15864
rect 23014 15852 23020 15864
rect 23072 15852 23078 15904
rect 23474 15852 23480 15904
rect 23532 15892 23538 15904
rect 24213 15895 24271 15901
rect 24213 15892 24225 15895
rect 23532 15864 24225 15892
rect 23532 15852 23538 15864
rect 24213 15861 24225 15864
rect 24259 15861 24271 15895
rect 24213 15855 24271 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 3878 15688 3884 15700
rect 3839 15660 3884 15688
rect 3878 15648 3884 15660
rect 3936 15648 3942 15700
rect 4246 15688 4252 15700
rect 4207 15660 4252 15688
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 4890 15648 4896 15700
rect 4948 15688 4954 15700
rect 5169 15691 5227 15697
rect 5169 15688 5181 15691
rect 4948 15660 5181 15688
rect 4948 15648 4954 15660
rect 5169 15657 5181 15660
rect 5215 15657 5227 15691
rect 5442 15688 5448 15700
rect 5169 15651 5227 15657
rect 5276 15660 5448 15688
rect 2961 15623 3019 15629
rect 2961 15589 2973 15623
rect 3007 15620 3019 15623
rect 3142 15620 3148 15632
rect 3007 15592 3148 15620
rect 3007 15589 3019 15592
rect 2961 15583 3019 15589
rect 3142 15580 3148 15592
rect 3200 15580 3206 15632
rect 3513 15623 3571 15629
rect 3513 15589 3525 15623
rect 3559 15620 3571 15623
rect 4154 15620 4160 15632
rect 3559 15592 4160 15620
rect 3559 15589 3571 15592
rect 3513 15583 3571 15589
rect 4154 15580 4160 15592
rect 4212 15580 4218 15632
rect 4338 15580 4344 15632
rect 4396 15620 4402 15632
rect 5276 15629 5304 15660
rect 5442 15648 5448 15660
rect 5500 15688 5506 15700
rect 5629 15691 5687 15697
rect 5629 15688 5641 15691
rect 5500 15660 5641 15688
rect 5500 15648 5506 15660
rect 5629 15657 5641 15660
rect 5675 15657 5687 15691
rect 5629 15651 5687 15657
rect 6454 15648 6460 15700
rect 6512 15688 6518 15700
rect 6730 15688 6736 15700
rect 6512 15660 6736 15688
rect 6512 15648 6518 15660
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 7285 15691 7343 15697
rect 7285 15657 7297 15691
rect 7331 15688 7343 15691
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 7331 15660 8309 15688
rect 7331 15657 7343 15660
rect 7285 15651 7343 15657
rect 8297 15657 8309 15660
rect 8343 15688 8355 15691
rect 8754 15688 8760 15700
rect 8343 15660 8760 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9824 15660 9873 15688
rect 9824 15648 9830 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 9861 15651 9919 15657
rect 10321 15691 10379 15697
rect 10321 15657 10333 15691
rect 10367 15688 10379 15691
rect 10686 15688 10692 15700
rect 10367 15660 10692 15688
rect 10367 15657 10379 15660
rect 10321 15651 10379 15657
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 10962 15688 10968 15700
rect 10923 15660 10968 15688
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 13081 15691 13139 15697
rect 13081 15657 13093 15691
rect 13127 15688 13139 15691
rect 13446 15688 13452 15700
rect 13127 15660 13452 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 14090 15688 14096 15700
rect 14051 15660 14096 15688
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 14734 15648 14740 15700
rect 14792 15688 14798 15700
rect 15013 15691 15071 15697
rect 15013 15688 15025 15691
rect 14792 15660 15025 15688
rect 14792 15648 14798 15660
rect 15013 15657 15025 15660
rect 15059 15657 15071 15691
rect 17129 15691 17187 15697
rect 17129 15688 17141 15691
rect 15013 15651 15071 15657
rect 15672 15660 17141 15688
rect 15672 15632 15700 15660
rect 17129 15657 17141 15660
rect 17175 15657 17187 15691
rect 17862 15688 17868 15700
rect 17823 15660 17868 15688
rect 17129 15651 17187 15657
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 18414 15688 18420 15700
rect 18375 15660 18420 15688
rect 18414 15648 18420 15660
rect 18472 15648 18478 15700
rect 20346 15648 20352 15700
rect 20404 15688 20410 15700
rect 21174 15688 21180 15700
rect 20404 15660 21180 15688
rect 20404 15648 20410 15660
rect 21174 15648 21180 15660
rect 21232 15688 21238 15700
rect 21453 15691 21511 15697
rect 21453 15688 21465 15691
rect 21232 15660 21465 15688
rect 21232 15648 21238 15660
rect 21453 15657 21465 15660
rect 21499 15657 21511 15691
rect 21453 15651 21511 15657
rect 23017 15691 23075 15697
rect 23017 15657 23029 15691
rect 23063 15688 23075 15691
rect 23198 15688 23204 15700
rect 23063 15660 23204 15688
rect 23063 15657 23075 15660
rect 23017 15651 23075 15657
rect 5261 15623 5319 15629
rect 5261 15620 5273 15623
rect 4396 15592 5273 15620
rect 4396 15580 4402 15592
rect 5261 15589 5273 15592
rect 5307 15589 5319 15623
rect 5261 15583 5319 15589
rect 6362 15580 6368 15632
rect 6420 15620 6426 15632
rect 6549 15623 6607 15629
rect 6549 15620 6561 15623
rect 6420 15592 6561 15620
rect 6420 15580 6426 15592
rect 6549 15589 6561 15592
rect 6595 15620 6607 15623
rect 6638 15620 6644 15632
rect 6595 15592 6644 15620
rect 6595 15589 6607 15592
rect 6549 15583 6607 15589
rect 6638 15580 6644 15592
rect 6696 15580 6702 15632
rect 9692 15592 11468 15620
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 3050 15552 3056 15564
rect 2963 15524 3056 15552
rect 3050 15512 3056 15524
rect 3108 15552 3114 15564
rect 3970 15552 3976 15564
rect 3108 15524 3976 15552
rect 3108 15512 3114 15524
rect 3970 15512 3976 15524
rect 4028 15552 4034 15564
rect 6178 15552 6184 15564
rect 4028 15524 6184 15552
rect 4028 15512 4034 15524
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 9692 15561 9720 15592
rect 10704 15564 10732 15592
rect 8113 15555 8171 15561
rect 8113 15552 8125 15555
rect 6288 15524 8125 15552
rect 2682 15444 2688 15496
rect 2740 15484 2746 15496
rect 2869 15487 2927 15493
rect 2869 15484 2881 15487
rect 2740 15456 2881 15484
rect 2740 15444 2746 15456
rect 2869 15453 2881 15456
rect 2915 15453 2927 15487
rect 2869 15447 2927 15453
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15484 5227 15487
rect 5258 15484 5264 15496
rect 5215 15456 5264 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 2498 15416 2504 15428
rect 2459 15388 2504 15416
rect 2498 15376 2504 15388
rect 2556 15376 2562 15428
rect 4614 15376 4620 15428
rect 4672 15416 4678 15428
rect 6288 15425 6316 15524
rect 8113 15521 8125 15524
rect 8159 15552 8171 15555
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 8159 15524 9137 15552
rect 8159 15521 8171 15524
rect 8113 15515 8171 15521
rect 9125 15521 9137 15524
rect 9171 15521 9183 15555
rect 9125 15515 9183 15521
rect 9677 15555 9735 15561
rect 9677 15521 9689 15555
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 10686 15512 10692 15564
rect 10744 15512 10750 15564
rect 11146 15512 11152 15564
rect 11204 15552 11210 15564
rect 11313 15555 11371 15561
rect 11313 15552 11325 15555
rect 11204 15524 11325 15552
rect 11204 15512 11210 15524
rect 11313 15521 11325 15524
rect 11359 15521 11371 15555
rect 11440 15552 11468 15592
rect 13814 15580 13820 15632
rect 13872 15620 13878 15632
rect 14185 15623 14243 15629
rect 14185 15620 14197 15623
rect 13872 15592 14197 15620
rect 13872 15580 13878 15592
rect 14185 15589 14197 15592
rect 14231 15620 14243 15623
rect 14550 15620 14556 15632
rect 14231 15592 14556 15620
rect 14231 15589 14243 15592
rect 14185 15583 14243 15589
rect 14550 15580 14556 15592
rect 14608 15580 14614 15632
rect 15194 15620 15200 15632
rect 14660 15592 15200 15620
rect 14660 15552 14688 15592
rect 15194 15580 15200 15592
rect 15252 15580 15258 15632
rect 15654 15620 15660 15632
rect 15615 15592 15660 15620
rect 15654 15580 15660 15592
rect 15712 15580 15718 15632
rect 15838 15620 15844 15632
rect 15799 15592 15844 15620
rect 15838 15580 15844 15592
rect 15896 15620 15902 15632
rect 16761 15623 16819 15629
rect 16761 15620 16773 15623
rect 15896 15592 16773 15620
rect 15896 15580 15902 15592
rect 16761 15589 16773 15592
rect 16807 15589 16819 15623
rect 16761 15583 16819 15589
rect 17586 15580 17592 15632
rect 17644 15620 17650 15632
rect 17681 15623 17739 15629
rect 17681 15620 17693 15623
rect 17644 15592 17693 15620
rect 17644 15580 17650 15592
rect 17681 15589 17693 15592
rect 17727 15589 17739 15623
rect 19426 15620 19432 15632
rect 19387 15592 19432 15620
rect 17681 15583 17739 15589
rect 19426 15580 19432 15592
rect 19484 15580 19490 15632
rect 21266 15580 21272 15632
rect 21324 15620 21330 15632
rect 23032 15620 23060 15651
rect 23198 15648 23204 15660
rect 23256 15648 23262 15700
rect 23661 15691 23719 15697
rect 23661 15657 23673 15691
rect 23707 15688 23719 15691
rect 23934 15688 23940 15700
rect 23707 15660 23940 15688
rect 23707 15657 23719 15660
rect 23661 15651 23719 15657
rect 23934 15648 23940 15660
rect 23992 15648 23998 15700
rect 24029 15691 24087 15697
rect 24029 15657 24041 15691
rect 24075 15688 24087 15691
rect 24394 15688 24400 15700
rect 24075 15660 24400 15688
rect 24075 15657 24087 15660
rect 24029 15651 24087 15657
rect 24394 15648 24400 15660
rect 24452 15648 24458 15700
rect 21324 15592 23060 15620
rect 21324 15580 21330 15592
rect 23750 15580 23756 15632
rect 23808 15620 23814 15632
rect 24673 15623 24731 15629
rect 24673 15620 24685 15623
rect 23808 15592 24685 15620
rect 23808 15580 23814 15592
rect 24673 15589 24685 15592
rect 24719 15620 24731 15623
rect 25133 15623 25191 15629
rect 25133 15620 25145 15623
rect 24719 15592 25145 15620
rect 24719 15589 24731 15592
rect 24673 15583 24731 15589
rect 25133 15589 25145 15592
rect 25179 15589 25191 15623
rect 25133 15583 25191 15589
rect 11440 15524 14688 15552
rect 14737 15555 14795 15561
rect 11313 15515 11371 15521
rect 14737 15521 14749 15555
rect 14783 15552 14795 15555
rect 14918 15552 14924 15564
rect 14783 15524 14924 15552
rect 14783 15521 14795 15524
rect 14737 15515 14795 15521
rect 14918 15512 14924 15524
rect 14976 15512 14982 15564
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 15933 15555 15991 15561
rect 15933 15552 15945 15555
rect 15436 15524 15945 15552
rect 15436 15512 15442 15524
rect 15933 15521 15945 15524
rect 15979 15552 15991 15555
rect 16390 15552 16396 15564
rect 15979 15524 16396 15552
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 20438 15552 20444 15564
rect 19352 15524 20444 15552
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6788 15456 6837 15484
rect 6788 15444 6794 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 7834 15484 7840 15496
rect 6825 15447 6883 15453
rect 7392 15456 7840 15484
rect 4709 15419 4767 15425
rect 4709 15416 4721 15419
rect 4672 15388 4721 15416
rect 4672 15376 4678 15388
rect 4709 15385 4721 15388
rect 4755 15385 4767 15419
rect 4709 15379 4767 15385
rect 6273 15419 6331 15425
rect 6273 15385 6285 15419
rect 6319 15385 6331 15419
rect 6273 15379 6331 15385
rect 7392 15360 7420 15456
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8478 15484 8484 15496
rect 8435 15456 8484 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 8478 15444 8484 15456
rect 8536 15484 8542 15496
rect 8757 15487 8815 15493
rect 8757 15484 8769 15487
rect 8536 15456 8769 15484
rect 8536 15444 8542 15456
rect 8757 15453 8769 15456
rect 8803 15453 8815 15487
rect 8757 15447 8815 15453
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15453 11115 15487
rect 11057 15447 11115 15453
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 6086 15348 6092 15360
rect 6047 15320 6092 15348
rect 6086 15308 6092 15320
rect 6144 15308 6150 15360
rect 7374 15308 7380 15360
rect 7432 15308 7438 15360
rect 7650 15348 7656 15360
rect 7611 15320 7656 15348
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 7834 15348 7840 15360
rect 7795 15320 7840 15348
rect 7834 15308 7840 15320
rect 7892 15308 7898 15360
rect 11072 15348 11100 15447
rect 13630 15416 13636 15428
rect 13591 15388 13636 15416
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 14108 15416 14136 15447
rect 14642 15444 14648 15496
rect 14700 15484 14706 15496
rect 16666 15484 16672 15496
rect 14700 15456 16672 15484
rect 14700 15444 14706 15456
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15484 18015 15487
rect 18046 15484 18052 15496
rect 18003 15456 18052 15484
rect 18003 15453 18015 15456
rect 17957 15447 18015 15453
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 19352 15493 19380 15524
rect 20438 15512 20444 15524
rect 20496 15512 20502 15564
rect 21893 15555 21951 15561
rect 21893 15552 21905 15555
rect 21008 15524 21905 15552
rect 21008 15496 21036 15524
rect 21893 15521 21905 15524
rect 21939 15521 21951 15555
rect 21893 15515 21951 15521
rect 24578 15512 24584 15564
rect 24636 15552 24642 15564
rect 24765 15555 24823 15561
rect 24765 15552 24777 15555
rect 24636 15524 24777 15552
rect 24636 15512 24642 15524
rect 24765 15521 24777 15524
rect 24811 15552 24823 15555
rect 24811 15524 25176 15552
rect 24811 15521 24823 15524
rect 24765 15515 24823 15521
rect 25148 15496 25176 15524
rect 19337 15487 19395 15493
rect 19337 15484 19349 15487
rect 18564 15456 19349 15484
rect 18564 15444 18570 15456
rect 19337 15453 19349 15456
rect 19383 15453 19395 15487
rect 19337 15447 19395 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15484 19579 15487
rect 19889 15487 19947 15493
rect 19889 15484 19901 15487
rect 19567 15456 19901 15484
rect 19567 15453 19579 15456
rect 19521 15447 19579 15453
rect 19889 15453 19901 15456
rect 19935 15484 19947 15487
rect 20990 15484 20996 15496
rect 19935 15456 20996 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 20990 15444 20996 15456
rect 21048 15444 21054 15496
rect 21450 15444 21456 15496
rect 21508 15484 21514 15496
rect 21637 15487 21695 15493
rect 21637 15484 21649 15487
rect 21508 15456 21649 15484
rect 21508 15444 21514 15456
rect 21637 15453 21649 15456
rect 21683 15453 21695 15487
rect 24670 15484 24676 15496
rect 24631 15456 24676 15484
rect 21637 15447 21695 15453
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 25130 15444 25136 15496
rect 25188 15444 25194 15496
rect 15381 15419 15439 15425
rect 15381 15416 15393 15419
rect 14108 15388 15393 15416
rect 15381 15385 15393 15388
rect 15427 15416 15439 15419
rect 16482 15416 16488 15428
rect 15427 15388 16488 15416
rect 15427 15385 15439 15388
rect 15381 15379 15439 15385
rect 16482 15376 16488 15388
rect 16540 15376 16546 15428
rect 16684 15416 16712 15444
rect 16684 15388 16896 15416
rect 16868 15360 16896 15388
rect 19242 15376 19248 15428
rect 19300 15416 19306 15428
rect 20257 15419 20315 15425
rect 20257 15416 20269 15419
rect 19300 15388 20269 15416
rect 19300 15376 19306 15388
rect 20257 15385 20269 15388
rect 20303 15385 20315 15419
rect 20257 15379 20315 15385
rect 20717 15419 20775 15425
rect 20717 15385 20729 15419
rect 20763 15416 20775 15419
rect 24210 15416 24216 15428
rect 20763 15388 21680 15416
rect 24171 15388 24216 15416
rect 20763 15385 20775 15388
rect 20717 15379 20775 15385
rect 11422 15348 11428 15360
rect 11072 15320 11428 15348
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 12434 15348 12440 15360
rect 12395 15320 12440 15348
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 16393 15351 16451 15357
rect 16393 15317 16405 15351
rect 16439 15348 16451 15351
rect 16666 15348 16672 15360
rect 16439 15320 16672 15348
rect 16439 15317 16451 15320
rect 16393 15311 16451 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 16850 15308 16856 15360
rect 16908 15308 16914 15360
rect 17405 15351 17463 15357
rect 17405 15317 17417 15351
rect 17451 15348 17463 15351
rect 17862 15348 17868 15360
rect 17451 15320 17868 15348
rect 17451 15317 17463 15320
rect 17405 15311 17463 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 18966 15348 18972 15360
rect 18927 15320 18972 15348
rect 18966 15308 18972 15320
rect 19024 15308 19030 15360
rect 21177 15351 21235 15357
rect 21177 15317 21189 15351
rect 21223 15348 21235 15351
rect 21266 15348 21272 15360
rect 21223 15320 21272 15348
rect 21223 15317 21235 15320
rect 21177 15311 21235 15317
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 21652 15348 21680 15388
rect 24210 15376 24216 15388
rect 24268 15376 24274 15428
rect 22002 15348 22008 15360
rect 21652 15320 22008 15348
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1762 15144 1768 15156
rect 1723 15116 1768 15144
rect 1762 15104 1768 15116
rect 1820 15144 1826 15156
rect 2682 15144 2688 15156
rect 1820 15116 2688 15144
rect 1820 15104 1826 15116
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 3050 15104 3056 15156
rect 3108 15144 3114 15156
rect 3329 15147 3387 15153
rect 3329 15144 3341 15147
rect 3108 15116 3341 15144
rect 3108 15104 3114 15116
rect 3329 15113 3341 15116
rect 3375 15113 3387 15147
rect 4338 15144 4344 15156
rect 4299 15116 4344 15144
rect 3329 15107 3387 15113
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 4893 15147 4951 15153
rect 4893 15113 4905 15147
rect 4939 15144 4951 15147
rect 5442 15144 5448 15156
rect 4939 15116 5448 15144
rect 4939 15113 4951 15116
rect 4893 15107 4951 15113
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 6273 15147 6331 15153
rect 6273 15113 6285 15147
rect 6319 15144 6331 15147
rect 6362 15144 6368 15156
rect 6319 15116 6368 15144
rect 6319 15113 6331 15116
rect 6273 15107 6331 15113
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 6454 15104 6460 15156
rect 6512 15144 6518 15156
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 6512 15116 6561 15144
rect 6512 15104 6518 15116
rect 6549 15113 6561 15116
rect 6595 15113 6607 15147
rect 6549 15107 6607 15113
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 7009 15147 7067 15153
rect 7009 15144 7021 15147
rect 6972 15116 7021 15144
rect 6972 15104 6978 15116
rect 7009 15113 7021 15116
rect 7055 15113 7067 15147
rect 7009 15107 7067 15113
rect 7469 15147 7527 15153
rect 7469 15113 7481 15147
rect 7515 15144 7527 15147
rect 7926 15144 7932 15156
rect 7515 15116 7932 15144
rect 7515 15113 7527 15116
rect 7469 15107 7527 15113
rect 2041 15079 2099 15085
rect 2041 15045 2053 15079
rect 2087 15076 2099 15079
rect 4706 15076 4712 15088
rect 2087 15048 3556 15076
rect 4619 15048 4712 15076
rect 2087 15045 2099 15048
rect 2041 15039 2099 15045
rect 1946 14968 1952 15020
rect 2004 15008 2010 15020
rect 2593 15011 2651 15017
rect 2593 15008 2605 15011
rect 2004 14980 2605 15008
rect 2004 14968 2010 14980
rect 2593 14977 2605 14980
rect 2639 15008 2651 15011
rect 2866 15008 2872 15020
rect 2639 14980 2872 15008
rect 2639 14977 2651 14980
rect 2593 14971 2651 14977
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 2314 14940 2320 14952
rect 2275 14912 2320 14940
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 3528 14949 3556 15048
rect 4706 15036 4712 15048
rect 4764 15076 4770 15088
rect 5258 15076 5264 15088
rect 4764 15048 5264 15076
rect 4764 15036 4770 15048
rect 5258 15036 5264 15048
rect 5316 15036 5322 15088
rect 3786 14968 3792 15020
rect 3844 14968 3850 15020
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 5445 15011 5503 15017
rect 5445 15008 5457 15011
rect 5408 14980 5457 15008
rect 5408 14968 5414 14980
rect 5445 14977 5457 14980
rect 5491 14977 5503 15011
rect 5445 14971 5503 14977
rect 3513 14943 3571 14949
rect 3513 14909 3525 14943
rect 3559 14940 3571 14943
rect 3804 14940 3832 14968
rect 3559 14912 3832 14940
rect 3559 14909 3571 14912
rect 3513 14903 3571 14909
rect 5074 14900 5080 14952
rect 5132 14940 5138 14952
rect 5169 14943 5227 14949
rect 5169 14940 5181 14943
rect 5132 14912 5181 14940
rect 5132 14900 5138 14912
rect 5169 14909 5181 14912
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6512 14912 6837 14940
rect 6512 14900 6518 14912
rect 6825 14909 6837 14912
rect 6871 14940 6883 14943
rect 7484 14940 7512 15107
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10505 15147 10563 15153
rect 10505 15144 10517 15147
rect 10192 15116 10517 15144
rect 10192 15104 10198 15116
rect 10505 15113 10517 15116
rect 10551 15113 10563 15147
rect 10505 15107 10563 15113
rect 10778 15104 10784 15156
rect 10836 15144 10842 15156
rect 13633 15147 13691 15153
rect 10836 15116 13584 15144
rect 10836 15104 10842 15116
rect 12526 15076 12532 15088
rect 12487 15048 12532 15076
rect 12526 15036 12532 15048
rect 12584 15036 12590 15088
rect 13556 15076 13584 15116
rect 13633 15113 13645 15147
rect 13679 15144 13691 15147
rect 13814 15144 13820 15156
rect 13679 15116 13820 15144
rect 13679 15113 13691 15116
rect 13633 15107 13691 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 14090 15144 14096 15156
rect 14051 15116 14096 15144
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 15197 15147 15255 15153
rect 15197 15113 15209 15147
rect 15243 15144 15255 15147
rect 16942 15144 16948 15156
rect 15243 15116 16948 15144
rect 15243 15113 15255 15116
rect 15197 15107 15255 15113
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17497 15147 17555 15153
rect 17497 15113 17509 15147
rect 17543 15144 17555 15147
rect 17586 15144 17592 15156
rect 17543 15116 17592 15144
rect 17543 15113 17555 15116
rect 17497 15107 17555 15113
rect 17586 15104 17592 15116
rect 17644 15104 17650 15156
rect 17770 15144 17776 15156
rect 17731 15116 17776 15144
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 18969 15147 19027 15153
rect 18969 15113 18981 15147
rect 19015 15144 19027 15147
rect 19058 15144 19064 15156
rect 19015 15116 19064 15144
rect 19015 15113 19027 15116
rect 18969 15107 19027 15113
rect 19058 15104 19064 15116
rect 19116 15104 19122 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 20990 15144 20996 15156
rect 20772 15116 20996 15144
rect 20772 15104 20778 15116
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 21082 15104 21088 15156
rect 21140 15144 21146 15156
rect 21637 15147 21695 15153
rect 21637 15144 21649 15147
rect 21140 15116 21649 15144
rect 21140 15104 21146 15116
rect 21637 15113 21649 15116
rect 21683 15113 21695 15147
rect 23014 15144 23020 15156
rect 22975 15116 23020 15144
rect 21637 15107 21695 15113
rect 23014 15104 23020 15116
rect 23072 15104 23078 15156
rect 23198 15104 23204 15156
rect 23256 15144 23262 15156
rect 23385 15147 23443 15153
rect 23385 15144 23397 15147
rect 23256 15116 23397 15144
rect 23256 15104 23262 15116
rect 23385 15113 23397 15116
rect 23431 15113 23443 15147
rect 23385 15107 23443 15113
rect 18506 15076 18512 15088
rect 13556 15048 18512 15076
rect 18506 15036 18512 15048
rect 18564 15036 18570 15088
rect 23400 15076 23428 15107
rect 23566 15104 23572 15156
rect 23624 15144 23630 15156
rect 23753 15147 23811 15153
rect 23753 15144 23765 15147
rect 23624 15116 23765 15144
rect 23624 15104 23630 15116
rect 23753 15113 23765 15116
rect 23799 15113 23811 15147
rect 23753 15107 23811 15113
rect 24765 15147 24823 15153
rect 24765 15113 24777 15147
rect 24811 15144 24823 15147
rect 25130 15144 25136 15156
rect 24811 15116 25136 15144
rect 24811 15113 24823 15116
rect 24765 15107 24823 15113
rect 25130 15104 25136 15116
rect 25188 15104 25194 15156
rect 23400 15048 24348 15076
rect 9953 15011 10011 15017
rect 6871 14912 7512 14940
rect 7576 14980 8044 15008
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 2222 14832 2228 14884
rect 2280 14872 2286 14884
rect 2501 14875 2559 14881
rect 2501 14872 2513 14875
rect 2280 14844 2513 14872
rect 2280 14832 2286 14844
rect 2501 14841 2513 14844
rect 2547 14841 2559 14875
rect 3786 14872 3792 14884
rect 3747 14844 3792 14872
rect 2501 14835 2559 14841
rect 3786 14832 3792 14844
rect 3844 14832 3850 14884
rect 3878 14832 3884 14884
rect 3936 14872 3942 14884
rect 5905 14875 5963 14881
rect 3936 14844 5488 14872
rect 3936 14832 3942 14844
rect 3053 14807 3111 14813
rect 3053 14773 3065 14807
rect 3099 14804 3111 14807
rect 3142 14804 3148 14816
rect 3099 14776 3148 14804
rect 3099 14773 3111 14776
rect 3053 14767 3111 14773
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 5166 14764 5172 14816
rect 5224 14804 5230 14816
rect 5353 14807 5411 14813
rect 5353 14804 5365 14807
rect 5224 14776 5365 14804
rect 5224 14764 5230 14776
rect 5353 14773 5365 14776
rect 5399 14773 5411 14807
rect 5460 14804 5488 14844
rect 5905 14841 5917 14875
rect 5951 14872 5963 14875
rect 6730 14872 6736 14884
rect 5951 14844 6736 14872
rect 5951 14841 5963 14844
rect 5905 14835 5963 14841
rect 6730 14832 6736 14844
rect 6788 14832 6794 14884
rect 7576 14872 7604 14980
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14909 7987 14943
rect 8016 14940 8044 14980
rect 9953 14977 9965 15011
rect 9999 15008 10011 15011
rect 11054 15008 11060 15020
rect 9999 14980 11060 15008
rect 9999 14977 10011 14980
rect 9953 14971 10011 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 12894 15008 12900 15020
rect 11931 14980 12900 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 15654 15008 15660 15020
rect 13504 14980 15660 15008
rect 13504 14968 13510 14980
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 16666 14968 16672 15020
rect 16724 15008 16730 15020
rect 16945 15011 17003 15017
rect 16945 15008 16957 15011
rect 16724 14980 16957 15008
rect 16724 14968 16730 14980
rect 16945 14977 16957 14980
rect 16991 15008 17003 15011
rect 17034 15008 17040 15020
rect 16991 14980 17040 15008
rect 16991 14977 17003 14980
rect 16945 14971 17003 14977
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18049 15011 18107 15017
rect 18049 15008 18061 15011
rect 18012 14980 18061 15008
rect 18012 14968 18018 14980
rect 18049 14977 18061 14980
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 20438 14968 20444 15020
rect 20496 15008 20502 15020
rect 21634 15008 21640 15020
rect 20496 14980 21640 15008
rect 20496 14968 20502 14980
rect 21634 14968 21640 14980
rect 21692 14968 21698 15020
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 23382 15008 23388 15020
rect 22143 14980 23388 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 23382 14968 23388 14980
rect 23440 14968 23446 15020
rect 24320 15017 24348 15048
rect 24305 15011 24363 15017
rect 24305 14977 24317 15011
rect 24351 14977 24363 15011
rect 24305 14971 24363 14977
rect 9582 14940 9588 14952
rect 8016 14912 9588 14940
rect 7929 14903 7987 14909
rect 6840 14844 7604 14872
rect 6840 14804 6868 14844
rect 7944 14816 7972 14903
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 9916 14912 11008 14940
rect 9916 14900 9922 14912
rect 8196 14875 8254 14881
rect 8196 14841 8208 14875
rect 8242 14872 8254 14875
rect 8478 14872 8484 14884
rect 8242 14844 8484 14872
rect 8242 14841 8254 14844
rect 8196 14835 8254 14841
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 10321 14875 10379 14881
rect 10321 14841 10333 14875
rect 10367 14872 10379 14875
rect 10778 14872 10784 14884
rect 10367 14844 10784 14872
rect 10367 14841 10379 14844
rect 10321 14835 10379 14841
rect 10778 14832 10784 14844
rect 10836 14832 10842 14884
rect 10980 14881 11008 14912
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 13081 14943 13139 14949
rect 13081 14940 13093 14943
rect 12124 14912 13093 14940
rect 12124 14900 12130 14912
rect 13081 14909 13093 14912
rect 13127 14909 13139 14943
rect 13081 14903 13139 14909
rect 15933 14943 15991 14949
rect 15933 14909 15945 14943
rect 15979 14940 15991 14943
rect 15979 14912 17080 14940
rect 15979 14909 15991 14912
rect 15933 14903 15991 14909
rect 10965 14875 11023 14881
rect 10965 14841 10977 14875
rect 11011 14841 11023 14875
rect 12250 14872 12256 14884
rect 12163 14844 12256 14872
rect 10965 14835 11023 14841
rect 12250 14832 12256 14844
rect 12308 14872 12314 14884
rect 12989 14875 13047 14881
rect 12989 14872 13001 14875
rect 12308 14844 13001 14872
rect 12308 14832 12314 14844
rect 12989 14841 13001 14844
rect 13035 14872 13047 14875
rect 14366 14872 14372 14884
rect 13035 14844 14372 14872
rect 13035 14841 13047 14844
rect 12989 14835 13047 14841
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 14642 14872 14648 14884
rect 14603 14844 14648 14872
rect 14642 14832 14648 14844
rect 14700 14872 14706 14884
rect 15013 14875 15071 14881
rect 15013 14872 15025 14875
rect 14700 14844 15025 14872
rect 14700 14832 14706 14844
rect 15013 14841 15025 14844
rect 15059 14841 15071 14875
rect 15013 14835 15071 14841
rect 16467 14875 16525 14881
rect 16467 14841 16479 14875
rect 16513 14872 16525 14875
rect 16666 14872 16672 14884
rect 16513 14844 16672 14872
rect 16513 14841 16525 14844
rect 16467 14835 16525 14841
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 16942 14872 16948 14884
rect 16903 14844 16948 14872
rect 16942 14832 16948 14844
rect 17000 14832 17006 14884
rect 17052 14881 17080 14912
rect 18782 14900 18788 14952
rect 18840 14940 18846 14952
rect 19061 14943 19119 14949
rect 19061 14940 19073 14943
rect 18840 14912 19073 14940
rect 18840 14900 18846 14912
rect 19061 14909 19073 14912
rect 19107 14909 19119 14943
rect 19061 14903 19119 14909
rect 21174 14900 21180 14952
rect 21232 14940 21238 14952
rect 22189 14943 22247 14949
rect 22189 14940 22201 14943
rect 21232 14912 22201 14940
rect 21232 14900 21238 14912
rect 22189 14909 22201 14912
rect 22235 14940 22247 14943
rect 22557 14943 22615 14949
rect 22557 14940 22569 14943
rect 22235 14912 22569 14940
rect 22235 14909 22247 14912
rect 22189 14903 22247 14909
rect 22557 14909 22569 14912
rect 22603 14909 22615 14943
rect 23290 14940 23296 14952
rect 22557 14903 22615 14909
rect 22664 14912 23296 14940
rect 17037 14875 17095 14881
rect 17037 14841 17049 14875
rect 17083 14872 17095 14875
rect 17218 14872 17224 14884
rect 17083 14844 17224 14872
rect 17083 14841 17095 14844
rect 17037 14835 17095 14841
rect 17218 14832 17224 14844
rect 17276 14832 17282 14884
rect 19328 14875 19386 14881
rect 19328 14841 19340 14875
rect 19374 14872 19386 14875
rect 19426 14872 19432 14884
rect 19374 14844 19432 14872
rect 19374 14841 19386 14844
rect 19328 14835 19386 14841
rect 19426 14832 19432 14844
rect 19484 14872 19490 14884
rect 19886 14872 19892 14884
rect 19484 14844 19892 14872
rect 19484 14832 19490 14844
rect 19886 14832 19892 14844
rect 19944 14832 19950 14884
rect 22002 14832 22008 14884
rect 22060 14872 22066 14884
rect 22097 14875 22155 14881
rect 22097 14872 22109 14875
rect 22060 14844 22109 14872
rect 22060 14832 22066 14844
rect 22097 14841 22109 14844
rect 22143 14872 22155 14875
rect 22664 14872 22692 14912
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 25041 14943 25099 14949
rect 25041 14940 25053 14943
rect 24044 14912 25053 14940
rect 24044 14884 24072 14912
rect 25041 14909 25053 14912
rect 25087 14909 25099 14943
rect 25041 14903 25099 14909
rect 25130 14900 25136 14952
rect 25188 14940 25194 14952
rect 25225 14943 25283 14949
rect 25225 14940 25237 14943
rect 25188 14912 25237 14940
rect 25188 14900 25194 14912
rect 25225 14909 25237 14912
rect 25271 14940 25283 14943
rect 25961 14943 26019 14949
rect 25961 14940 25973 14943
rect 25271 14912 25973 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25961 14909 25973 14912
rect 26007 14909 26019 14943
rect 25961 14903 26019 14909
rect 22143 14844 22692 14872
rect 22143 14841 22155 14844
rect 22097 14835 22155 14841
rect 23014 14832 23020 14884
rect 23072 14872 23078 14884
rect 24026 14872 24032 14884
rect 23072 14844 23520 14872
rect 23987 14844 24032 14872
rect 23072 14832 23078 14844
rect 5460 14776 6868 14804
rect 5353 14767 5411 14773
rect 7190 14764 7196 14816
rect 7248 14804 7254 14816
rect 7837 14807 7895 14813
rect 7837 14804 7849 14807
rect 7248 14776 7849 14804
rect 7248 14764 7254 14776
rect 7837 14773 7849 14776
rect 7883 14804 7895 14807
rect 7926 14804 7932 14816
rect 7883 14776 7932 14804
rect 7883 14773 7895 14776
rect 7837 14767 7895 14773
rect 7926 14764 7932 14776
rect 7984 14764 7990 14816
rect 9306 14804 9312 14816
rect 9267 14776 9312 14804
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 11517 14807 11575 14813
rect 11517 14804 11529 14807
rect 11480 14776 11529 14804
rect 11480 14764 11486 14776
rect 11517 14773 11529 14776
rect 11563 14804 11575 14807
rect 11882 14804 11888 14816
rect 11563 14776 11888 14804
rect 11563 14773 11575 14776
rect 11517 14767 11575 14773
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 14274 14764 14280 14816
rect 14332 14804 14338 14816
rect 14553 14807 14611 14813
rect 14553 14804 14565 14807
rect 14332 14776 14565 14804
rect 14332 14764 14338 14776
rect 14553 14773 14565 14776
rect 14599 14804 14611 14807
rect 15197 14807 15255 14813
rect 15197 14804 15209 14807
rect 14599 14776 15209 14804
rect 14599 14773 14611 14776
rect 14553 14767 14611 14773
rect 15197 14773 15209 14776
rect 15243 14773 15255 14807
rect 15378 14804 15384 14816
rect 15339 14776 15384 14804
rect 15197 14767 15255 14773
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 16301 14807 16359 14813
rect 16301 14773 16313 14807
rect 16347 14804 16359 14807
rect 16960 14804 16988 14832
rect 16347 14776 16988 14804
rect 16347 14773 16359 14776
rect 16301 14767 16359 14773
rect 20070 14764 20076 14816
rect 20128 14804 20134 14816
rect 20441 14807 20499 14813
rect 20441 14804 20453 14807
rect 20128 14776 20453 14804
rect 20128 14764 20134 14776
rect 20441 14773 20453 14776
rect 20487 14773 20499 14807
rect 21450 14804 21456 14816
rect 21363 14776 21456 14804
rect 20441 14767 20499 14773
rect 21450 14764 21456 14776
rect 21508 14804 21514 14816
rect 22646 14804 22652 14816
rect 21508 14776 22652 14804
rect 21508 14764 21514 14776
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 22738 14764 22744 14816
rect 22796 14804 22802 14816
rect 23290 14804 23296 14816
rect 22796 14776 23296 14804
rect 22796 14764 22802 14776
rect 23290 14764 23296 14776
rect 23348 14764 23354 14816
rect 23492 14804 23520 14844
rect 24026 14832 24032 14844
rect 24084 14832 24090 14884
rect 25498 14872 25504 14884
rect 25459 14844 25504 14872
rect 25498 14832 25504 14844
rect 25556 14832 25562 14884
rect 24213 14807 24271 14813
rect 24213 14804 24225 14807
rect 23492 14776 24225 14804
rect 24213 14773 24225 14776
rect 24259 14773 24271 14807
rect 24213 14767 24271 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2866 14600 2872 14612
rect 2827 14572 2872 14600
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 5166 14600 5172 14612
rect 4764 14572 5172 14600
rect 4764 14560 4770 14572
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 6638 14600 6644 14612
rect 6599 14572 6644 14600
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 6914 14600 6920 14612
rect 6875 14572 6920 14600
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 8846 14600 8852 14612
rect 8807 14572 8852 14600
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10229 14603 10287 14609
rect 10229 14600 10241 14603
rect 9824 14572 10241 14600
rect 9824 14560 9830 14572
rect 10229 14569 10241 14572
rect 10275 14569 10287 14603
rect 11146 14600 11152 14612
rect 11107 14572 11152 14600
rect 10229 14563 10287 14569
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 11422 14560 11428 14612
rect 11480 14600 11486 14612
rect 11698 14600 11704 14612
rect 11480 14572 11704 14600
rect 11480 14560 11486 14572
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 11793 14603 11851 14609
rect 11793 14569 11805 14603
rect 11839 14600 11851 14603
rect 12066 14600 12072 14612
rect 11839 14572 12072 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 1670 14532 1676 14544
rect 1504 14504 1676 14532
rect 1504 14473 1532 14504
rect 1670 14492 1676 14504
rect 1728 14532 1734 14544
rect 2590 14532 2596 14544
rect 1728 14504 2596 14532
rect 1728 14492 1734 14504
rect 2590 14492 2596 14504
rect 2648 14492 2654 14544
rect 4338 14492 4344 14544
rect 4396 14532 4402 14544
rect 5442 14532 5448 14544
rect 4396 14504 5448 14532
rect 4396 14492 4402 14504
rect 5442 14492 5448 14504
rect 5500 14532 5506 14544
rect 5721 14535 5779 14541
rect 5721 14532 5733 14535
rect 5500 14504 5733 14532
rect 5500 14492 5506 14504
rect 5721 14501 5733 14504
rect 5767 14501 5779 14535
rect 5721 14495 5779 14501
rect 8294 14492 8300 14544
rect 8352 14532 8358 14544
rect 8389 14535 8447 14541
rect 8389 14532 8401 14535
rect 8352 14504 8401 14532
rect 8352 14492 8358 14504
rect 8389 14501 8401 14504
rect 8435 14532 8447 14535
rect 9217 14535 9275 14541
rect 9217 14532 9229 14535
rect 8435 14504 9229 14532
rect 8435 14501 8447 14504
rect 8389 14495 8447 14501
rect 9217 14501 9229 14504
rect 9263 14501 9275 14535
rect 9217 14495 9275 14501
rect 10042 14492 10048 14544
rect 10100 14532 10106 14544
rect 11808 14532 11836 14563
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 16669 14603 16727 14609
rect 16669 14569 16681 14603
rect 16715 14600 16727 14603
rect 16758 14600 16764 14612
rect 16715 14572 16764 14600
rect 16715 14569 16727 14572
rect 16669 14563 16727 14569
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 17954 14560 17960 14612
rect 18012 14600 18018 14612
rect 18325 14603 18383 14609
rect 18325 14600 18337 14603
rect 18012 14572 18337 14600
rect 18012 14560 18018 14572
rect 18325 14569 18337 14572
rect 18371 14600 18383 14603
rect 19242 14600 19248 14612
rect 18371 14572 19248 14600
rect 18371 14569 18383 14572
rect 18325 14563 18383 14569
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19426 14600 19432 14612
rect 19387 14572 19432 14600
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 19889 14603 19947 14609
rect 19889 14569 19901 14603
rect 19935 14600 19947 14603
rect 19978 14600 19984 14612
rect 19935 14572 19984 14600
rect 19935 14569 19947 14572
rect 19889 14563 19947 14569
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20254 14600 20260 14612
rect 20215 14572 20260 14600
rect 20254 14560 20260 14572
rect 20312 14560 20318 14612
rect 20714 14600 20720 14612
rect 20675 14572 20720 14600
rect 20714 14560 20720 14572
rect 20772 14600 20778 14612
rect 20772 14572 21588 14600
rect 20772 14560 20778 14572
rect 10100 14504 11836 14532
rect 10100 14492 10106 14504
rect 15194 14492 15200 14544
rect 15252 14532 15258 14544
rect 15534 14535 15592 14541
rect 15534 14532 15546 14535
rect 15252 14504 15546 14532
rect 15252 14492 15258 14504
rect 15534 14501 15546 14504
rect 15580 14532 15592 14535
rect 15654 14532 15660 14544
rect 15580 14504 15660 14532
rect 15580 14501 15592 14504
rect 15534 14495 15592 14501
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 17862 14492 17868 14544
rect 17920 14532 17926 14544
rect 17920 14504 20760 14532
rect 17920 14492 17926 14504
rect 20732 14476 20760 14504
rect 21358 14492 21364 14544
rect 21416 14532 21422 14544
rect 21560 14541 21588 14572
rect 21726 14560 21732 14612
rect 21784 14600 21790 14612
rect 22002 14600 22008 14612
rect 21784 14572 22008 14600
rect 21784 14560 21790 14572
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 22741 14603 22799 14609
rect 22741 14569 22753 14603
rect 22787 14600 22799 14603
rect 23382 14600 23388 14612
rect 22787 14572 23388 14600
rect 22787 14569 22799 14572
rect 22741 14563 22799 14569
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 24673 14603 24731 14609
rect 24673 14569 24685 14603
rect 24719 14569 24731 14603
rect 24673 14563 24731 14569
rect 21453 14535 21511 14541
rect 21453 14532 21465 14535
rect 21416 14504 21465 14532
rect 21416 14492 21422 14504
rect 21453 14501 21465 14504
rect 21499 14501 21511 14535
rect 21453 14495 21511 14501
rect 21545 14535 21603 14541
rect 21545 14501 21557 14535
rect 21591 14532 21603 14535
rect 21634 14532 21640 14544
rect 21591 14504 21640 14532
rect 21591 14501 21603 14504
rect 21545 14495 21603 14501
rect 21634 14492 21640 14504
rect 21692 14532 21698 14544
rect 21913 14535 21971 14541
rect 21913 14532 21925 14535
rect 21692 14504 21925 14532
rect 21692 14492 21698 14504
rect 21913 14501 21925 14504
rect 21959 14532 21971 14535
rect 24688 14532 24716 14563
rect 21959 14504 24716 14532
rect 21959 14501 21971 14504
rect 21913 14495 21971 14501
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14433 1547 14467
rect 1489 14427 1547 14433
rect 1756 14467 1814 14473
rect 1756 14433 1768 14467
rect 1802 14464 1814 14467
rect 3050 14464 3056 14476
rect 1802 14436 3056 14464
rect 1802 14433 1814 14436
rect 1756 14427 1814 14433
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4706 14464 4712 14476
rect 4111 14436 4712 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14464 5595 14467
rect 6086 14464 6092 14476
rect 5583 14436 6092 14464
rect 5583 14433 5595 14436
rect 5537 14427 5595 14433
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 6638 14424 6644 14476
rect 6696 14464 6702 14476
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 6696 14436 6745 14464
rect 6696 14424 6702 14436
rect 6733 14433 6745 14436
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 7377 14467 7435 14473
rect 7377 14433 7389 14467
rect 7423 14464 7435 14467
rect 7650 14464 7656 14476
rect 7423 14436 7656 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 7650 14424 7656 14436
rect 7708 14464 7714 14476
rect 9306 14464 9312 14476
rect 7708 14436 9312 14464
rect 7708 14424 7714 14436
rect 9306 14424 9312 14436
rect 9364 14464 9370 14476
rect 9364 14436 10364 14464
rect 9364 14424 9370 14436
rect 3142 14356 3148 14408
rect 3200 14396 3206 14408
rect 3200 14368 4844 14396
rect 3200 14356 3206 14368
rect 3881 14331 3939 14337
rect 3881 14297 3893 14331
rect 3927 14328 3939 14331
rect 4154 14328 4160 14340
rect 3927 14300 4160 14328
rect 3927 14297 3939 14300
rect 3881 14291 3939 14297
rect 4154 14288 4160 14300
rect 4212 14288 4218 14340
rect 3050 14220 3056 14272
rect 3108 14260 3114 14272
rect 3421 14263 3479 14269
rect 3421 14260 3433 14263
rect 3108 14232 3433 14260
rect 3108 14220 3114 14232
rect 3421 14229 3433 14232
rect 3467 14229 3479 14263
rect 4246 14260 4252 14272
rect 4207 14232 4252 14260
rect 3421 14223 3479 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 4706 14260 4712 14272
rect 4667 14232 4712 14260
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 4816 14260 4844 14368
rect 4982 14356 4988 14408
rect 5040 14396 5046 14408
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 5040 14368 5089 14396
rect 5040 14356 5046 14368
rect 5077 14365 5089 14368
rect 5123 14396 5135 14399
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 5123 14368 5825 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5813 14365 5825 14368
rect 5859 14396 5871 14399
rect 6178 14396 6184 14408
rect 5859 14368 6184 14396
rect 5859 14365 5871 14368
rect 5813 14359 5871 14365
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 8386 14396 8392 14408
rect 8347 14368 8392 14396
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 10336 14405 10364 14436
rect 11146 14424 11152 14476
rect 11204 14464 11210 14476
rect 12141 14467 12199 14473
rect 12141 14464 12153 14467
rect 11204 14436 12153 14464
rect 11204 14424 11210 14436
rect 12141 14433 12153 14436
rect 12187 14464 12199 14467
rect 12434 14464 12440 14476
rect 12187 14436 12440 14464
rect 12187 14433 12199 14436
rect 12141 14427 12199 14433
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 14734 14424 14740 14476
rect 14792 14464 14798 14476
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 14792 14436 15301 14464
rect 14792 14424 14798 14436
rect 15289 14433 15301 14436
rect 15335 14464 15347 14467
rect 15378 14464 15384 14476
rect 15335 14436 15384 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 19702 14464 19708 14476
rect 19663 14436 19708 14464
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 20162 14424 20168 14476
rect 20220 14464 20226 14476
rect 20438 14464 20444 14476
rect 20220 14436 20444 14464
rect 20220 14424 20226 14436
rect 20438 14424 20444 14436
rect 20496 14424 20502 14476
rect 20714 14424 20720 14476
rect 20772 14424 20778 14476
rect 23382 14424 23388 14476
rect 23440 14464 23446 14476
rect 23549 14467 23607 14473
rect 23549 14464 23561 14467
rect 23440 14436 23561 14464
rect 23440 14424 23446 14436
rect 23549 14433 23561 14436
rect 23595 14433 23607 14467
rect 23549 14427 23607 14433
rect 10137 14399 10195 14405
rect 8536 14368 8581 14396
rect 8536 14356 8542 14368
rect 10137 14365 10149 14399
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10502 14396 10508 14408
rect 10367 14368 10508 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 4890 14288 4896 14340
rect 4948 14328 4954 14340
rect 5261 14331 5319 14337
rect 5261 14328 5273 14331
rect 4948 14300 5273 14328
rect 4948 14288 4954 14300
rect 5261 14297 5273 14300
rect 5307 14297 5319 14331
rect 5261 14291 5319 14297
rect 6273 14331 6331 14337
rect 6273 14297 6285 14331
rect 6319 14328 6331 14331
rect 7929 14331 7987 14337
rect 7929 14328 7941 14331
rect 6319 14300 7941 14328
rect 6319 14297 6331 14300
rect 6273 14291 6331 14297
rect 7929 14297 7941 14300
rect 7975 14328 7987 14331
rect 10152 14328 10180 14359
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 11882 14396 11888 14408
rect 11843 14368 11888 14396
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 18230 14396 18236 14408
rect 18191 14368 18236 14396
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 18414 14396 18420 14408
rect 18375 14368 18420 14396
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 21453 14399 21511 14405
rect 21453 14365 21465 14399
rect 21499 14396 21511 14399
rect 21726 14396 21732 14408
rect 21499 14368 21732 14396
rect 21499 14365 21511 14368
rect 21453 14359 21511 14365
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 22646 14356 22652 14408
rect 22704 14396 22710 14408
rect 23293 14399 23351 14405
rect 23293 14396 23305 14399
rect 22704 14368 23305 14396
rect 22704 14356 22710 14368
rect 23293 14365 23305 14368
rect 23339 14365 23351 14399
rect 23293 14359 23351 14365
rect 7975 14300 10180 14328
rect 7975 14297 7987 14300
rect 7929 14291 7987 14297
rect 14366 14288 14372 14340
rect 14424 14328 14430 14340
rect 14461 14331 14519 14337
rect 14461 14328 14473 14331
rect 14424 14300 14473 14328
rect 14424 14288 14430 14300
rect 14461 14297 14473 14300
rect 14507 14328 14519 14331
rect 15194 14328 15200 14340
rect 14507 14300 15200 14328
rect 14507 14297 14519 14300
rect 14461 14291 14519 14297
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 17405 14331 17463 14337
rect 17405 14297 17417 14331
rect 17451 14328 17463 14331
rect 18046 14328 18052 14340
rect 17451 14300 18052 14328
rect 17451 14297 17463 14300
rect 17405 14291 17463 14297
rect 18046 14288 18052 14300
rect 18104 14328 18110 14340
rect 18966 14328 18972 14340
rect 18104 14300 18972 14328
rect 18104 14288 18110 14300
rect 18966 14288 18972 14300
rect 19024 14288 19030 14340
rect 20990 14328 20996 14340
rect 20951 14300 20996 14328
rect 20990 14288 20996 14300
rect 21048 14288 21054 14340
rect 7190 14260 7196 14272
rect 4816 14232 7196 14260
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 7745 14263 7803 14269
rect 7745 14229 7757 14263
rect 7791 14260 7803 14263
rect 7834 14260 7840 14272
rect 7791 14232 7840 14260
rect 7791 14229 7803 14232
rect 7745 14223 7803 14229
rect 7834 14220 7840 14232
rect 7892 14260 7898 14272
rect 8478 14260 8484 14272
rect 7892 14232 8484 14260
rect 7892 14220 7898 14232
rect 8478 14220 8484 14232
rect 8536 14220 8542 14272
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 9769 14263 9827 14269
rect 9769 14260 9781 14263
rect 9732 14232 9781 14260
rect 9732 14220 9738 14232
rect 9769 14229 9781 14232
rect 9815 14229 9827 14263
rect 9769 14223 9827 14229
rect 10781 14263 10839 14269
rect 10781 14229 10793 14263
rect 10827 14260 10839 14263
rect 10962 14260 10968 14272
rect 10827 14232 10968 14260
rect 10827 14229 10839 14232
rect 10781 14223 10839 14229
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 12066 14260 12072 14272
rect 11388 14232 12072 14260
rect 11388 14220 11394 14232
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 13170 14220 13176 14272
rect 13228 14260 13234 14272
rect 13265 14263 13323 14269
rect 13265 14260 13277 14263
rect 13228 14232 13277 14260
rect 13228 14220 13234 14232
rect 13265 14229 13277 14232
rect 13311 14229 13323 14263
rect 13265 14223 13323 14229
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 14001 14263 14059 14269
rect 14001 14260 14013 14263
rect 13504 14232 14013 14260
rect 13504 14220 13510 14232
rect 14001 14229 14013 14232
rect 14047 14260 14059 14263
rect 14274 14260 14280 14272
rect 14047 14232 14280 14260
rect 14047 14229 14059 14232
rect 14001 14223 14059 14229
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 14734 14260 14740 14272
rect 14695 14232 14740 14260
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 16758 14220 16764 14272
rect 16816 14260 16822 14272
rect 17865 14263 17923 14269
rect 17865 14260 17877 14263
rect 16816 14232 17877 14260
rect 16816 14220 16822 14232
rect 17865 14229 17877 14232
rect 17911 14229 17923 14263
rect 17865 14223 17923 14229
rect 18782 14220 18788 14272
rect 18840 14260 18846 14272
rect 19061 14263 19119 14269
rect 19061 14260 19073 14263
rect 18840 14232 19073 14260
rect 18840 14220 18846 14232
rect 19061 14229 19073 14232
rect 19107 14229 19119 14263
rect 22278 14260 22284 14272
rect 22239 14232 22284 14260
rect 19061 14223 19119 14229
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 23017 14263 23075 14269
rect 23017 14260 23029 14263
rect 22796 14232 23029 14260
rect 22796 14220 22802 14232
rect 23017 14229 23029 14232
rect 23063 14229 23075 14263
rect 25222 14260 25228 14272
rect 25183 14232 25228 14260
rect 23017 14223 23075 14229
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 3050 14056 3056 14068
rect 3011 14028 3056 14056
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 3697 14059 3755 14065
rect 3697 14025 3709 14059
rect 3743 14056 3755 14059
rect 3970 14056 3976 14068
rect 3743 14028 3976 14056
rect 3743 14025 3755 14028
rect 3697 14019 3755 14025
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4890 14016 4896 14068
rect 4948 14056 4954 14068
rect 5258 14056 5264 14068
rect 4948 14028 5264 14056
rect 4948 14016 4954 14028
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 6638 14056 6644 14068
rect 6599 14028 6644 14056
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 7101 14059 7159 14065
rect 7101 14025 7113 14059
rect 7147 14056 7159 14059
rect 8202 14056 8208 14068
rect 7147 14028 8208 14056
rect 7147 14025 7159 14028
rect 7101 14019 7159 14025
rect 8202 14016 8208 14028
rect 8260 14016 8266 14068
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 9953 14059 10011 14065
rect 9953 14056 9965 14059
rect 8536 14028 9965 14056
rect 8536 14016 8542 14028
rect 9953 14025 9965 14028
rect 9999 14056 10011 14059
rect 10042 14056 10048 14068
rect 9999 14028 10048 14056
rect 9999 14025 10011 14028
rect 9953 14019 10011 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10502 14056 10508 14068
rect 10463 14028 10508 14056
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 13078 14056 13084 14068
rect 12952 14028 13084 14056
rect 12952 14016 12958 14028
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 14461 14059 14519 14065
rect 14461 14025 14473 14059
rect 14507 14056 14519 14059
rect 14550 14056 14556 14068
rect 14507 14028 14556 14056
rect 14507 14025 14519 14028
rect 14461 14019 14519 14025
rect 14550 14016 14556 14028
rect 14608 14016 14614 14068
rect 16482 14056 16488 14068
rect 16443 14028 16488 14056
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 18506 14056 18512 14068
rect 18419 14028 18512 14056
rect 18506 14016 18512 14028
rect 18564 14056 18570 14068
rect 18782 14056 18788 14068
rect 18564 14028 18788 14056
rect 18564 14016 18570 14028
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19702 14016 19708 14068
rect 19760 14056 19766 14068
rect 20625 14059 20683 14065
rect 20625 14056 20637 14059
rect 19760 14028 20637 14056
rect 19760 14016 19766 14028
rect 20625 14025 20637 14028
rect 20671 14056 20683 14059
rect 21082 14056 21088 14068
rect 20671 14028 21088 14056
rect 20671 14025 20683 14028
rect 20625 14019 20683 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 21177 14059 21235 14065
rect 21177 14025 21189 14059
rect 21223 14056 21235 14059
rect 21450 14056 21456 14068
rect 21223 14028 21456 14056
rect 21223 14025 21235 14028
rect 21177 14019 21235 14025
rect 21450 14016 21456 14028
rect 21508 14056 21514 14068
rect 22278 14056 22284 14068
rect 21508 14028 22284 14056
rect 21508 14016 21514 14028
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 23014 14056 23020 14068
rect 22975 14028 23020 14056
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 23753 14059 23811 14065
rect 23753 14025 23765 14059
rect 23799 14056 23811 14059
rect 24670 14056 24676 14068
rect 23799 14028 24676 14056
rect 23799 14025 23811 14028
rect 23753 14019 23811 14025
rect 24670 14016 24676 14028
rect 24728 14056 24734 14068
rect 25222 14056 25228 14068
rect 24728 14028 25228 14056
rect 24728 14016 24734 14028
rect 25222 14016 25228 14028
rect 25280 14016 25286 14068
rect 25406 14056 25412 14068
rect 25367 14028 25412 14056
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 5902 13948 5908 14000
rect 5960 13988 5966 14000
rect 8018 13988 8024 14000
rect 5960 13960 8024 13988
rect 5960 13948 5966 13960
rect 8018 13948 8024 13960
rect 8076 13948 8082 14000
rect 8113 13991 8171 13997
rect 8113 13957 8125 13991
rect 8159 13988 8171 13991
rect 8386 13988 8392 14000
rect 8159 13960 8392 13988
rect 8159 13957 8171 13960
rect 8113 13951 8171 13957
rect 8386 13948 8392 13960
rect 8444 13948 8450 14000
rect 16206 13948 16212 14000
rect 16264 13988 16270 14000
rect 17405 13991 17463 13997
rect 17405 13988 17417 13991
rect 16264 13960 17417 13988
rect 16264 13948 16270 13960
rect 17405 13957 17417 13960
rect 17451 13957 17463 13991
rect 17405 13951 17463 13957
rect 21358 13948 21364 14000
rect 21416 13988 21422 14000
rect 22097 13991 22155 13997
rect 22097 13988 22109 13991
rect 21416 13960 22109 13988
rect 21416 13948 21422 13960
rect 22097 13957 22109 13960
rect 22143 13957 22155 13991
rect 22097 13951 22155 13957
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 4065 13923 4123 13929
rect 4065 13889 4077 13923
rect 4111 13920 4123 13923
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 4111 13892 4169 13920
rect 4111 13889 4123 13892
rect 4065 13883 4123 13889
rect 4157 13889 4169 13892
rect 4203 13889 4215 13923
rect 7650 13920 7656 13932
rect 4157 13883 4215 13889
rect 6564 13892 7512 13920
rect 7611 13892 7656 13920
rect 4172 13852 4200 13883
rect 6564 13852 6592 13892
rect 4172 13824 6592 13852
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 7484 13852 7512 13892
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 16298 13920 16304 13932
rect 16211 13892 16304 13920
rect 16298 13880 16304 13892
rect 16356 13920 16362 13932
rect 16942 13920 16948 13932
rect 16356 13892 16948 13920
rect 16356 13880 16362 13892
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17218 13920 17224 13932
rect 17083 13892 17224 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 7926 13852 7932 13864
rect 6696 13824 6960 13852
rect 7484 13824 7932 13852
rect 6696 13812 6702 13824
rect 1946 13793 1952 13796
rect 1940 13784 1952 13793
rect 1907 13756 1952 13784
rect 1940 13747 1952 13756
rect 1946 13744 1952 13747
rect 2004 13744 2010 13796
rect 2038 13744 2044 13796
rect 2096 13784 2102 13796
rect 2406 13784 2412 13796
rect 2096 13756 2412 13784
rect 2096 13744 2102 13756
rect 2406 13744 2412 13756
rect 2464 13744 2470 13796
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 4402 13787 4460 13793
rect 4402 13784 4414 13787
rect 4028 13756 4414 13784
rect 4028 13744 4034 13756
rect 4402 13753 4414 13756
rect 4448 13753 4460 13787
rect 4402 13747 4460 13753
rect 4614 13744 4620 13796
rect 4672 13784 4678 13796
rect 4982 13784 4988 13796
rect 4672 13756 4988 13784
rect 4672 13744 4678 13756
rect 4982 13744 4988 13756
rect 5040 13744 5046 13796
rect 6932 13784 6960 13824
rect 7926 13812 7932 13824
rect 7984 13852 7990 13864
rect 8846 13861 8852 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 7984 13824 8401 13852
rect 7984 13812 7990 13824
rect 8389 13821 8401 13824
rect 8435 13852 8447 13855
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8435 13824 8585 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8840 13852 8852 13861
rect 8807 13824 8852 13852
rect 8573 13815 8631 13821
rect 8840 13815 8852 13824
rect 8846 13812 8852 13815
rect 8904 13812 8910 13864
rect 12250 13852 12256 13864
rect 11256 13824 12256 13852
rect 7377 13787 7435 13793
rect 7377 13784 7389 13787
rect 6932 13756 7389 13784
rect 7377 13753 7389 13756
rect 7423 13753 7435 13787
rect 7558 13784 7564 13796
rect 7519 13756 7564 13784
rect 7377 13747 7435 13753
rect 7558 13744 7564 13756
rect 7616 13744 7622 13796
rect 7650 13744 7656 13796
rect 7708 13784 7714 13796
rect 11256 13784 11284 13824
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 15933 13855 15991 13861
rect 15933 13821 15945 13855
rect 15979 13852 15991 13855
rect 17052 13852 17080 13883
rect 17218 13880 17224 13892
rect 17276 13920 17282 13932
rect 17865 13923 17923 13929
rect 17865 13920 17877 13923
rect 17276 13892 17877 13920
rect 17276 13880 17282 13892
rect 17865 13889 17877 13892
rect 17911 13920 17923 13923
rect 18414 13920 18420 13932
rect 17911 13892 18420 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 18414 13880 18420 13892
rect 18472 13920 18478 13932
rect 20993 13923 21051 13929
rect 18472 13892 18736 13920
rect 18472 13880 18478 13892
rect 15979 13824 17080 13852
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 7708 13756 11284 13784
rect 11333 13787 11391 13793
rect 7708 13744 7714 13756
rect 11333 13753 11345 13787
rect 11379 13784 11391 13787
rect 11514 13784 11520 13796
rect 11379 13756 11520 13784
rect 11379 13753 11391 13756
rect 11333 13747 11391 13753
rect 11514 13744 11520 13756
rect 11572 13744 11578 13796
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 6086 13716 6092 13728
rect 6047 13688 6092 13716
rect 6086 13676 6092 13688
rect 6144 13676 6150 13728
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 7098 13716 7104 13728
rect 6880 13688 7104 13716
rect 6880 13676 6886 13688
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 8110 13676 8116 13728
rect 8168 13716 8174 13728
rect 9582 13716 9588 13728
rect 8168 13688 9588 13716
rect 8168 13676 8174 13688
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 11146 13716 11152 13728
rect 11107 13688 11152 13716
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11882 13676 11888 13728
rect 11940 13716 11946 13728
rect 11977 13719 12035 13725
rect 11977 13716 11989 13719
rect 11940 13688 11989 13716
rect 11940 13676 11946 13688
rect 11977 13685 11989 13688
rect 12023 13716 12035 13719
rect 12989 13719 13047 13725
rect 12989 13716 13001 13719
rect 12023 13688 13001 13716
rect 12023 13685 12035 13688
rect 11977 13679 12035 13685
rect 12989 13685 13001 13688
rect 13035 13716 13047 13719
rect 13096 13716 13124 13815
rect 18506 13812 18512 13864
rect 18564 13852 18570 13864
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18564 13824 18613 13852
rect 18564 13812 18570 13824
rect 18601 13821 18613 13824
rect 18647 13821 18659 13855
rect 18708 13852 18736 13892
rect 20993 13889 21005 13923
rect 21039 13920 21051 13923
rect 21542 13920 21548 13932
rect 21039 13892 21548 13920
rect 21039 13889 21051 13892
rect 20993 13883 21051 13889
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 21634 13880 21640 13932
rect 21692 13920 21698 13932
rect 21729 13923 21787 13929
rect 21729 13920 21741 13923
rect 21692 13892 21741 13920
rect 21692 13880 21698 13892
rect 21729 13889 21741 13892
rect 21775 13889 21787 13923
rect 23032 13920 23060 14016
rect 24121 13923 24179 13929
rect 24121 13920 24133 13923
rect 23032 13892 24133 13920
rect 21729 13883 21787 13889
rect 24121 13889 24133 13892
rect 24167 13889 24179 13923
rect 24121 13883 24179 13889
rect 18708 13824 20024 13852
rect 18601 13815 18659 13821
rect 13170 13744 13176 13796
rect 13228 13784 13234 13796
rect 13326 13787 13384 13793
rect 13326 13784 13338 13787
rect 13228 13756 13338 13784
rect 13228 13744 13234 13756
rect 13326 13753 13338 13756
rect 13372 13753 13384 13787
rect 13326 13747 13384 13753
rect 16482 13744 16488 13796
rect 16540 13784 16546 13796
rect 16945 13787 17003 13793
rect 16945 13784 16957 13787
rect 16540 13756 16957 13784
rect 16540 13744 16546 13756
rect 16945 13753 16957 13756
rect 16991 13784 17003 13787
rect 17126 13784 17132 13796
rect 16991 13756 17132 13784
rect 16991 13753 17003 13756
rect 16945 13747 17003 13753
rect 17126 13744 17132 13756
rect 17184 13744 17190 13796
rect 18868 13787 18926 13793
rect 18868 13753 18880 13787
rect 18914 13784 18926 13787
rect 18966 13784 18972 13796
rect 18914 13756 18972 13784
rect 18914 13753 18926 13756
rect 18868 13747 18926 13753
rect 18966 13744 18972 13756
rect 19024 13744 19030 13796
rect 15378 13716 15384 13728
rect 13035 13688 15384 13716
rect 13035 13685 13047 13688
rect 12989 13679 13047 13685
rect 15378 13676 15384 13688
rect 15436 13716 15442 13728
rect 15838 13716 15844 13728
rect 15436 13688 15844 13716
rect 15436 13676 15442 13688
rect 15838 13676 15844 13688
rect 15896 13716 15902 13728
rect 16850 13716 16856 13728
rect 15896 13688 16856 13716
rect 15896 13676 15902 13688
rect 16850 13676 16856 13688
rect 16908 13676 16914 13728
rect 19996 13725 20024 13824
rect 21082 13812 21088 13864
rect 21140 13852 21146 13864
rect 21818 13852 21824 13864
rect 21140 13824 21824 13852
rect 21140 13812 21146 13824
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 22646 13852 22652 13864
rect 22607 13824 22652 13852
rect 22646 13812 22652 13824
rect 22704 13812 22710 13864
rect 23934 13812 23940 13864
rect 23992 13852 23998 13864
rect 24305 13855 24363 13861
rect 24305 13852 24317 13855
rect 23992 13824 24317 13852
rect 23992 13812 23998 13824
rect 24305 13821 24317 13824
rect 24351 13852 24363 13855
rect 24670 13852 24676 13864
rect 24351 13824 24676 13852
rect 24351 13821 24363 13824
rect 24305 13815 24363 13821
rect 24670 13812 24676 13824
rect 24728 13852 24734 13864
rect 25041 13855 25099 13861
rect 25041 13852 25053 13855
rect 24728 13824 25053 13852
rect 24728 13812 24734 13824
rect 25041 13821 25053 13824
rect 25087 13821 25099 13855
rect 25041 13815 25099 13821
rect 25225 13855 25283 13861
rect 25225 13821 25237 13855
rect 25271 13852 25283 13855
rect 25774 13852 25780 13864
rect 25271 13824 25780 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 25774 13812 25780 13824
rect 25832 13812 25838 13864
rect 22186 13744 22192 13796
rect 22244 13784 22250 13796
rect 22922 13784 22928 13796
rect 22244 13756 22928 13784
rect 22244 13744 22250 13756
rect 22922 13744 22928 13756
rect 22980 13744 22986 13796
rect 19981 13719 20039 13725
rect 19981 13685 19993 13719
rect 20027 13716 20039 13719
rect 20162 13716 20168 13728
rect 20027 13688 20168 13716
rect 20027 13685 20039 13688
rect 19981 13679 20039 13685
rect 20162 13676 20168 13688
rect 20220 13676 20226 13728
rect 21637 13719 21695 13725
rect 21637 13685 21649 13719
rect 21683 13716 21695 13719
rect 22554 13716 22560 13728
rect 21683 13688 22560 13716
rect 21683 13685 21695 13688
rect 21637 13679 21695 13685
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 23474 13716 23480 13728
rect 23435 13688 23480 13716
rect 23474 13676 23480 13688
rect 23532 13716 23538 13728
rect 24213 13719 24271 13725
rect 24213 13716 24225 13719
rect 23532 13688 24225 13716
rect 23532 13676 23538 13688
rect 24213 13685 24225 13688
rect 24259 13685 24271 13719
rect 24213 13679 24271 13685
rect 24578 13676 24584 13728
rect 24636 13716 24642 13728
rect 24673 13719 24731 13725
rect 24673 13716 24685 13719
rect 24636 13688 24685 13716
rect 24636 13676 24642 13688
rect 24673 13685 24685 13688
rect 24719 13685 24731 13719
rect 24673 13679 24731 13685
rect 24762 13676 24768 13728
rect 24820 13716 24826 13728
rect 25958 13716 25964 13728
rect 24820 13688 25964 13716
rect 24820 13676 24826 13688
rect 25958 13676 25964 13688
rect 26016 13676 26022 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 1728 13484 1869 13512
rect 1728 13472 1734 13484
rect 1857 13481 1869 13484
rect 1903 13512 1915 13515
rect 2225 13515 2283 13521
rect 2225 13512 2237 13515
rect 1903 13484 2237 13512
rect 1903 13481 1915 13484
rect 1857 13475 1915 13481
rect 2225 13481 2237 13484
rect 2271 13512 2283 13515
rect 2590 13512 2596 13524
rect 2271 13484 2596 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 2682 13472 2688 13524
rect 2740 13512 2746 13524
rect 2961 13515 3019 13521
rect 2961 13512 2973 13515
rect 2740 13484 2973 13512
rect 2740 13472 2746 13484
rect 2961 13481 2973 13484
rect 3007 13512 3019 13515
rect 3326 13512 3332 13524
rect 3007 13484 3332 13512
rect 3007 13481 3019 13484
rect 2961 13475 3019 13481
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 5261 13515 5319 13521
rect 5261 13481 5273 13515
rect 5307 13512 5319 13515
rect 5442 13512 5448 13524
rect 5307 13484 5448 13512
rect 5307 13481 5319 13484
rect 5261 13475 5319 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5736 13484 7236 13512
rect 3050 13404 3056 13456
rect 3108 13444 3114 13456
rect 5736 13444 5764 13484
rect 5902 13444 5908 13456
rect 3108 13416 3153 13444
rect 3344 13416 5764 13444
rect 5863 13416 5908 13444
rect 3108 13404 3114 13416
rect 3344 13388 3372 13416
rect 5902 13404 5908 13416
rect 5960 13404 5966 13456
rect 6362 13404 6368 13456
rect 6420 13444 6426 13456
rect 6420 13416 6960 13444
rect 6420 13404 6426 13416
rect 1946 13336 1952 13388
rect 2004 13376 2010 13388
rect 2004 13348 3280 13376
rect 2004 13336 2010 13348
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 3142 13308 3148 13320
rect 3007 13280 3148 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 3252 13308 3280 13348
rect 3326 13336 3332 13388
rect 3384 13336 3390 13388
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 5534 13376 5540 13388
rect 4172 13348 5540 13376
rect 3513 13311 3571 13317
rect 3513 13308 3525 13311
rect 3252 13280 3525 13308
rect 3513 13277 3525 13280
rect 3559 13308 3571 13311
rect 4172 13308 4200 13348
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 5721 13379 5779 13385
rect 5721 13345 5733 13379
rect 5767 13376 5779 13379
rect 6454 13376 6460 13388
rect 5767 13348 6460 13376
rect 5767 13345 5779 13348
rect 5721 13339 5779 13345
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 6932 13385 6960 13416
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7098 13376 7104 13388
rect 6963 13348 7104 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 7208 13376 7236 13484
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 8110 13512 8116 13524
rect 7524 13484 8116 13512
rect 7524 13472 7530 13484
rect 8110 13472 8116 13484
rect 8168 13512 8174 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 8168 13484 8585 13512
rect 8168 13472 8174 13484
rect 8573 13481 8585 13484
rect 8619 13481 8631 13515
rect 8573 13475 8631 13481
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 9030 13512 9036 13524
rect 8904 13484 9036 13512
rect 8904 13472 8910 13484
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 9861 13515 9919 13521
rect 9861 13481 9873 13515
rect 9907 13512 9919 13515
rect 10042 13512 10048 13524
rect 9907 13484 10048 13512
rect 9907 13481 9919 13484
rect 9861 13475 9919 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 11422 13512 11428 13524
rect 10336 13484 11428 13512
rect 10336 13456 10364 13484
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 13170 13512 13176 13524
rect 13131 13484 13176 13512
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 14185 13515 14243 13521
rect 14185 13512 14197 13515
rect 14056 13484 14197 13512
rect 14056 13472 14062 13484
rect 14185 13481 14197 13484
rect 14231 13481 14243 13515
rect 16482 13512 16488 13524
rect 14185 13475 14243 13481
rect 15212 13484 16488 13512
rect 8665 13447 8723 13453
rect 8665 13413 8677 13447
rect 8711 13444 8723 13447
rect 8754 13444 8760 13456
rect 8711 13416 8760 13444
rect 8711 13413 8723 13416
rect 8665 13407 8723 13413
rect 8754 13404 8760 13416
rect 8812 13444 8818 13456
rect 9582 13444 9588 13456
rect 8812 13416 9588 13444
rect 8812 13404 8818 13416
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 10318 13404 10324 13456
rect 10376 13404 10382 13456
rect 11054 13444 11060 13456
rect 10520 13416 11060 13444
rect 7208 13348 9536 13376
rect 4338 13308 4344 13320
rect 3559 13280 4200 13308
rect 4299 13280 4344 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5997 13311 6055 13317
rect 5132 13280 5488 13308
rect 5132 13268 5138 13280
rect 2314 13200 2320 13252
rect 2372 13240 2378 13252
rect 2501 13243 2559 13249
rect 2501 13240 2513 13243
rect 2372 13212 2513 13240
rect 2372 13200 2378 13212
rect 2501 13209 2513 13212
rect 2547 13209 2559 13243
rect 2501 13203 2559 13209
rect 4893 13243 4951 13249
rect 4893 13209 4905 13243
rect 4939 13240 4951 13243
rect 5350 13240 5356 13252
rect 4939 13212 5356 13240
rect 4939 13209 4951 13212
rect 4893 13203 4951 13209
rect 5350 13200 5356 13212
rect 5408 13200 5414 13252
rect 5460 13249 5488 13280
rect 5997 13277 6009 13311
rect 6043 13308 6055 13311
rect 6178 13308 6184 13320
rect 6043 13280 6184 13308
rect 6043 13277 6055 13280
rect 5997 13271 6055 13277
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 8018 13308 8024 13320
rect 7524 13280 8024 13308
rect 7524 13268 7530 13280
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 8570 13308 8576 13320
rect 8531 13280 8576 13308
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 9508 13308 9536 13348
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 10520 13376 10548 13416
rect 11054 13404 11060 13416
rect 11112 13404 11118 13456
rect 11238 13404 11244 13456
rect 11296 13444 11302 13456
rect 11701 13447 11759 13453
rect 11701 13444 11713 13447
rect 11296 13416 11713 13444
rect 11296 13404 11302 13416
rect 9732 13348 10548 13376
rect 9732 13336 9738 13348
rect 10594 13336 10600 13388
rect 10652 13376 10658 13388
rect 11517 13379 11575 13385
rect 11517 13376 11529 13379
rect 10652 13348 11529 13376
rect 10652 13336 10658 13348
rect 11517 13345 11529 13348
rect 11563 13345 11575 13379
rect 11517 13339 11575 13345
rect 11624 13320 11652 13416
rect 11701 13413 11713 13416
rect 11747 13413 11759 13447
rect 11701 13407 11759 13413
rect 14090 13404 14096 13456
rect 14148 13444 14154 13456
rect 15212 13444 15240 13484
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 16758 13512 16764 13524
rect 16719 13484 16764 13512
rect 16758 13472 16764 13484
rect 16816 13472 16822 13524
rect 19426 13512 19432 13524
rect 19387 13484 19432 13512
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 21450 13512 21456 13524
rect 21411 13484 21456 13512
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 22278 13512 22284 13524
rect 22239 13484 22284 13512
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 22646 13472 22652 13524
rect 22704 13472 22710 13524
rect 23382 13472 23388 13524
rect 23440 13512 23446 13524
rect 24029 13515 24087 13521
rect 24029 13512 24041 13515
rect 23440 13484 24041 13512
rect 23440 13472 23446 13484
rect 24029 13481 24041 13484
rect 24075 13512 24087 13515
rect 24578 13512 24584 13524
rect 24075 13484 24584 13512
rect 24075 13481 24087 13484
rect 24029 13475 24087 13481
rect 24578 13472 24584 13484
rect 24636 13472 24642 13524
rect 24854 13472 24860 13524
rect 24912 13512 24918 13524
rect 25317 13515 25375 13521
rect 25317 13512 25329 13515
rect 24912 13484 25329 13512
rect 24912 13472 24918 13484
rect 25317 13481 25329 13484
rect 25363 13481 25375 13515
rect 25317 13475 25375 13481
rect 15930 13444 15936 13456
rect 14148 13416 15240 13444
rect 15891 13416 15936 13444
rect 14148 13404 14154 13416
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 17218 13453 17224 13456
rect 17212 13444 17224 13453
rect 17179 13416 17224 13444
rect 17212 13407 17224 13416
rect 17218 13404 17224 13407
rect 17276 13404 17282 13456
rect 18966 13444 18972 13456
rect 18879 13416 18972 13444
rect 18966 13404 18972 13416
rect 19024 13444 19030 13456
rect 20070 13444 20076 13456
rect 19024 13416 20076 13444
rect 19024 13404 19030 13416
rect 20070 13404 20076 13416
rect 20128 13404 20134 13456
rect 21174 13404 21180 13456
rect 21232 13444 21238 13456
rect 21269 13447 21327 13453
rect 21269 13444 21281 13447
rect 21232 13416 21281 13444
rect 21232 13404 21238 13416
rect 21269 13413 21281 13416
rect 21315 13413 21327 13447
rect 21269 13407 21327 13413
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 12400 13348 14657 13376
rect 12400 13336 12406 13348
rect 14645 13345 14657 13348
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 15105 13379 15163 13385
rect 15105 13376 15117 13379
rect 14792 13348 15117 13376
rect 14792 13336 14798 13348
rect 15105 13345 15117 13348
rect 15151 13376 15163 13379
rect 15654 13376 15660 13388
rect 15151 13348 15660 13376
rect 15151 13345 15163 13348
rect 15105 13339 15163 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 15749 13379 15807 13385
rect 15749 13345 15761 13379
rect 15795 13376 15807 13379
rect 16482 13376 16488 13388
rect 15795 13348 16488 13376
rect 15795 13345 15807 13348
rect 15749 13339 15807 13345
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 16945 13379 17003 13385
rect 16945 13376 16957 13379
rect 16908 13348 16957 13376
rect 16908 13336 16914 13348
rect 16945 13345 16957 13348
rect 16991 13376 17003 13379
rect 17494 13376 17500 13388
rect 16991 13348 17500 13376
rect 16991 13345 17003 13348
rect 16945 13339 17003 13345
rect 17494 13336 17500 13348
rect 17552 13376 17558 13388
rect 18506 13376 18512 13388
rect 17552 13348 18512 13376
rect 17552 13336 17558 13348
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 19242 13336 19248 13388
rect 19300 13376 19306 13388
rect 19426 13376 19432 13388
rect 19300 13348 19432 13376
rect 19300 13336 19306 13348
rect 19426 13336 19432 13348
rect 19484 13336 19490 13388
rect 22005 13379 22063 13385
rect 22005 13345 22017 13379
rect 22051 13376 22063 13379
rect 22554 13376 22560 13388
rect 22051 13348 22560 13376
rect 22051 13345 22063 13348
rect 22005 13339 22063 13345
rect 22554 13336 22560 13348
rect 22612 13336 22618 13388
rect 22664 13385 22692 13472
rect 22922 13453 22928 13456
rect 22916 13444 22928 13453
rect 22883 13416 22928 13444
rect 22916 13407 22928 13416
rect 22922 13404 22928 13407
rect 22980 13404 22986 13456
rect 22656 13379 22714 13385
rect 22656 13345 22668 13379
rect 22702 13345 22714 13379
rect 22656 13339 22714 13345
rect 23934 13336 23940 13388
rect 23992 13376 23998 13388
rect 25038 13376 25044 13388
rect 23992 13348 25044 13376
rect 23992 13336 23998 13348
rect 25038 13336 25044 13348
rect 25096 13376 25102 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 25096 13348 25145 13376
rect 25096 13336 25102 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 11606 13308 11612 13320
rect 9508 13280 11612 13308
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 11790 13308 11796 13320
rect 11751 13280 11796 13308
rect 11790 13268 11796 13280
rect 11848 13308 11854 13320
rect 12529 13311 12587 13317
rect 12529 13308 12541 13311
rect 11848 13280 12541 13308
rect 11848 13268 11854 13280
rect 12529 13277 12541 13280
rect 12575 13308 12587 13311
rect 13078 13308 13084 13320
rect 12575 13280 13084 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 13906 13268 13912 13320
rect 13964 13308 13970 13320
rect 14185 13311 14243 13317
rect 14185 13308 14197 13311
rect 13964 13280 14197 13308
rect 13964 13268 13970 13280
rect 14185 13277 14197 13280
rect 14231 13277 14243 13311
rect 14185 13271 14243 13277
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14550 13308 14556 13320
rect 14323 13280 14556 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 5445 13243 5503 13249
rect 5445 13209 5457 13243
rect 5491 13209 5503 13243
rect 5445 13203 5503 13209
rect 5902 13200 5908 13252
rect 5960 13200 5966 13252
rect 6086 13200 6092 13252
rect 6144 13240 6150 13252
rect 6733 13243 6791 13249
rect 6733 13240 6745 13243
rect 6144 13212 6745 13240
rect 6144 13200 6150 13212
rect 6733 13209 6745 13212
rect 6779 13209 6791 13243
rect 6733 13203 6791 13209
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 7101 13243 7159 13249
rect 7101 13240 7113 13243
rect 6880 13212 7113 13240
rect 6880 13200 6886 13212
rect 7101 13209 7113 13212
rect 7147 13209 7159 13243
rect 8113 13243 8171 13249
rect 7101 13203 7159 13209
rect 7576 13212 8064 13240
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 3970 13172 3976 13184
rect 3927 13144 3976 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 5074 13132 5080 13184
rect 5132 13172 5138 13184
rect 5920 13172 5948 13200
rect 7576 13184 7604 13212
rect 6362 13172 6368 13184
rect 5132 13144 5948 13172
rect 6323 13144 6368 13172
rect 5132 13132 5138 13144
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 7558 13172 7564 13184
rect 7519 13144 7564 13172
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 7834 13172 7840 13184
rect 7795 13144 7840 13172
rect 7834 13132 7840 13144
rect 7892 13132 7898 13184
rect 8036 13172 8064 13212
rect 8113 13209 8125 13243
rect 8159 13240 8171 13243
rect 8202 13240 8208 13252
rect 8159 13212 8208 13240
rect 8159 13209 8171 13212
rect 8113 13203 8171 13209
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 9493 13243 9551 13249
rect 9493 13209 9505 13243
rect 9539 13240 9551 13243
rect 11238 13240 11244 13252
rect 9539 13212 11244 13240
rect 9539 13209 9551 13212
rect 9493 13203 9551 13209
rect 11238 13200 11244 13212
rect 11296 13200 11302 13252
rect 13722 13240 13728 13252
rect 13683 13212 13728 13240
rect 13722 13200 13728 13212
rect 13780 13200 13786 13252
rect 14200 13240 14228 13271
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 16022 13308 16028 13320
rect 15983 13280 16028 13308
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 21450 13268 21456 13320
rect 21508 13308 21514 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 21508 13280 21557 13308
rect 21508 13268 21514 13280
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 24946 13308 24952 13320
rect 24907 13280 24952 13308
rect 21545 13271 21603 13277
rect 24946 13268 24952 13280
rect 25004 13268 25010 13320
rect 14734 13240 14740 13252
rect 14200 13212 14740 13240
rect 14734 13200 14740 13212
rect 14792 13200 14798 13252
rect 15473 13243 15531 13249
rect 15473 13209 15485 13243
rect 15519 13240 15531 13243
rect 15746 13240 15752 13252
rect 15519 13212 15752 13240
rect 15519 13209 15531 13212
rect 15473 13203 15531 13209
rect 15746 13200 15752 13212
rect 15804 13200 15810 13252
rect 20530 13200 20536 13252
rect 20588 13240 20594 13252
rect 20993 13243 21051 13249
rect 20993 13240 21005 13243
rect 20588 13212 21005 13240
rect 20588 13200 20594 13212
rect 20993 13209 21005 13212
rect 21039 13209 21051 13243
rect 20993 13203 21051 13209
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8036 13144 9045 13172
rect 9033 13141 9045 13144
rect 9079 13172 9091 13175
rect 9306 13172 9312 13184
rect 9079 13144 9312 13172
rect 9079 13141 9091 13144
rect 9033 13135 9091 13141
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 10502 13172 10508 13184
rect 10463 13144 10508 13172
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 10873 13175 10931 13181
rect 10873 13141 10885 13175
rect 10919 13172 10931 13175
rect 11422 13172 11428 13184
rect 10919 13144 11428 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 13538 13172 13544 13184
rect 13499 13144 13544 13172
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 18322 13172 18328 13184
rect 18283 13144 18328 13172
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 19334 13172 19340 13184
rect 19295 13144 19340 13172
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 20073 13175 20131 13181
rect 20073 13141 20085 13175
rect 20119 13172 20131 13175
rect 20162 13172 20168 13184
rect 20119 13144 20168 13172
rect 20119 13141 20131 13144
rect 20073 13135 20131 13141
rect 20162 13132 20168 13144
rect 20220 13132 20226 13184
rect 20717 13175 20775 13181
rect 20717 13141 20729 13175
rect 20763 13172 20775 13175
rect 21266 13172 21272 13184
rect 20763 13144 21272 13172
rect 20763 13141 20775 13144
rect 20717 13135 20775 13141
rect 21266 13132 21272 13144
rect 21324 13172 21330 13184
rect 21726 13172 21732 13184
rect 21324 13144 21732 13172
rect 21324 13132 21330 13144
rect 21726 13132 21732 13144
rect 21784 13132 21790 13184
rect 24118 13132 24124 13184
rect 24176 13172 24182 13184
rect 24581 13175 24639 13181
rect 24581 13172 24593 13175
rect 24176 13144 24593 13172
rect 24176 13132 24182 13144
rect 24581 13141 24593 13144
rect 24627 13141 24639 13175
rect 24581 13135 24639 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1765 12971 1823 12977
rect 1765 12937 1777 12971
rect 1811 12968 1823 12971
rect 2222 12968 2228 12980
rect 1811 12940 2228 12968
rect 1811 12937 1823 12940
rect 1765 12931 1823 12937
rect 2222 12928 2228 12940
rect 2280 12928 2286 12980
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 5261 12971 5319 12977
rect 5261 12968 5273 12971
rect 4212 12940 5273 12968
rect 4212 12928 4218 12940
rect 5261 12937 5273 12940
rect 5307 12937 5319 12971
rect 5261 12931 5319 12937
rect 5997 12971 6055 12977
rect 5997 12937 6009 12971
rect 6043 12968 6055 12971
rect 6178 12968 6184 12980
rect 6043 12940 6184 12968
rect 6043 12937 6055 12940
rect 5997 12931 6055 12937
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 6273 12971 6331 12977
rect 6273 12937 6285 12971
rect 6319 12968 6331 12971
rect 6454 12968 6460 12980
rect 6319 12940 6460 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 6454 12928 6460 12940
rect 6512 12968 6518 12980
rect 6638 12968 6644 12980
rect 6512 12940 6644 12968
rect 6512 12928 6518 12940
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 6972 12940 7205 12968
rect 6972 12928 6978 12940
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 8110 12968 8116 12980
rect 8071 12940 8116 12968
rect 7193 12931 7251 12937
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8570 12968 8576 12980
rect 8483 12940 8576 12968
rect 8570 12928 8576 12940
rect 8628 12968 8634 12980
rect 9214 12968 9220 12980
rect 8628 12940 9220 12968
rect 8628 12928 8634 12940
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 9677 12971 9735 12977
rect 9677 12968 9689 12971
rect 9640 12940 9689 12968
rect 9640 12928 9646 12940
rect 9677 12937 9689 12940
rect 9723 12937 9735 12971
rect 9677 12931 9735 12937
rect 10321 12971 10379 12977
rect 10321 12937 10333 12971
rect 10367 12968 10379 12971
rect 11790 12968 11796 12980
rect 10367 12940 11796 12968
rect 10367 12937 10379 12940
rect 10321 12931 10379 12937
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11940 12940 12173 12968
rect 11940 12928 11946 12940
rect 12161 12937 12173 12940
rect 12207 12968 12219 12971
rect 12207 12940 12940 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 3142 12860 3148 12912
rect 3200 12900 3206 12912
rect 3329 12903 3387 12909
rect 3329 12900 3341 12903
rect 3200 12872 3341 12900
rect 3200 12860 3206 12872
rect 3329 12869 3341 12872
rect 3375 12869 3387 12903
rect 5074 12900 5080 12912
rect 5035 12872 5080 12900
rect 3329 12863 3387 12869
rect 5074 12860 5080 12872
rect 5132 12860 5138 12912
rect 7834 12900 7840 12912
rect 5828 12872 7840 12900
rect 2314 12792 2320 12844
rect 2372 12832 2378 12844
rect 3050 12832 3056 12844
rect 2372 12804 3056 12832
rect 2372 12792 2378 12804
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 3602 12792 3608 12844
rect 3660 12832 3666 12844
rect 3878 12832 3884 12844
rect 3660 12804 3884 12832
rect 3660 12792 3666 12804
rect 3878 12792 3884 12804
rect 3936 12792 3942 12844
rect 5828 12841 5856 12872
rect 7834 12860 7840 12872
rect 7892 12860 7898 12912
rect 8754 12900 8760 12912
rect 8715 12872 8760 12900
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 9030 12860 9036 12912
rect 9088 12900 9094 12912
rect 10870 12900 10876 12912
rect 9088 12872 10456 12900
rect 10831 12872 10876 12900
rect 9088 12860 9094 12872
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12832 4399 12835
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 4387 12804 5825 12832
rect 4387 12801 4399 12804
rect 4341 12795 4399 12801
rect 5813 12801 5825 12804
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 7190 12832 7196 12844
rect 6512 12804 7196 12832
rect 6512 12792 6518 12804
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 7745 12835 7803 12841
rect 7745 12832 7757 12835
rect 7616 12804 7757 12832
rect 7616 12792 7622 12804
rect 7745 12801 7757 12804
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 9122 12832 9128 12844
rect 8628 12804 9128 12832
rect 8628 12792 8634 12804
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 2041 12767 2099 12773
rect 2041 12733 2053 12767
rect 2087 12764 2099 12767
rect 2774 12764 2780 12776
rect 2087 12736 2780 12764
rect 2087 12733 2099 12736
rect 2041 12727 2099 12733
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12764 4767 12767
rect 6822 12764 6828 12776
rect 4755 12736 6828 12764
rect 4755 12733 4767 12736
rect 4709 12727 4767 12733
rect 2314 12696 2320 12708
rect 2275 12668 2320 12696
rect 2314 12656 2320 12668
rect 2372 12656 2378 12708
rect 3145 12699 3203 12705
rect 3145 12665 3157 12699
rect 3191 12696 3203 12699
rect 3605 12699 3663 12705
rect 3605 12696 3617 12699
rect 3191 12668 3617 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 3605 12665 3617 12668
rect 3651 12696 3663 12699
rect 4062 12696 4068 12708
rect 3651 12668 4068 12696
rect 3651 12665 3663 12668
rect 3605 12659 3663 12665
rect 4062 12656 4068 12668
rect 4120 12696 4126 12708
rect 4246 12696 4252 12708
rect 4120 12668 4252 12696
rect 4120 12656 4126 12668
rect 4246 12656 4252 12668
rect 4304 12656 4310 12708
rect 5258 12656 5264 12708
rect 5316 12696 5322 12708
rect 5736 12705 5764 12736
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 7469 12767 7527 12773
rect 7469 12764 7481 12767
rect 7340 12736 7481 12764
rect 7340 12724 7346 12736
rect 7469 12733 7481 12736
rect 7515 12733 7527 12767
rect 7469 12727 7527 12733
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8720 12736 9045 12764
rect 8720 12724 8726 12736
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9306 12764 9312 12776
rect 9267 12736 9312 12764
rect 9033 12727 9091 12733
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 9582 12724 9588 12776
rect 9640 12764 9646 12776
rect 10318 12764 10324 12776
rect 9640 12736 10324 12764
rect 9640 12724 9646 12736
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 5537 12699 5595 12705
rect 5537 12696 5549 12699
rect 5316 12668 5549 12696
rect 5316 12656 5322 12668
rect 5537 12665 5549 12668
rect 5583 12665 5595 12699
rect 5537 12659 5595 12665
rect 5721 12699 5779 12705
rect 5721 12665 5733 12699
rect 5767 12665 5779 12699
rect 5994 12696 6000 12708
rect 5955 12668 6000 12696
rect 5721 12659 5779 12665
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 6641 12699 6699 12705
rect 6641 12665 6653 12699
rect 6687 12696 6699 12699
rect 7098 12696 7104 12708
rect 6687 12668 7104 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 7650 12696 7656 12708
rect 7611 12668 7656 12696
rect 7650 12656 7656 12668
rect 7708 12656 7714 12708
rect 9122 12656 9128 12708
rect 9180 12696 9186 12708
rect 9858 12696 9864 12708
rect 9180 12668 9864 12696
rect 9180 12656 9186 12668
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 2225 12631 2283 12637
rect 2225 12597 2237 12631
rect 2271 12628 2283 12631
rect 2406 12628 2412 12640
rect 2271 12600 2412 12628
rect 2271 12597 2283 12600
rect 2225 12591 2283 12597
rect 2406 12588 2412 12600
rect 2464 12588 2470 12640
rect 2777 12631 2835 12637
rect 2777 12597 2789 12631
rect 2823 12628 2835 12631
rect 3786 12628 3792 12640
rect 2823 12600 3792 12628
rect 2823 12597 2835 12600
rect 2777 12591 2835 12597
rect 3786 12588 3792 12600
rect 3844 12628 3850 12640
rect 5074 12628 5080 12640
rect 3844 12600 5080 12628
rect 3844 12588 3850 12600
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 7116 12628 7144 12656
rect 7926 12628 7932 12640
rect 7116 12600 7932 12628
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 9217 12631 9275 12637
rect 9217 12628 9229 12631
rect 8904 12600 9229 12628
rect 8904 12588 8910 12600
rect 9217 12597 9229 12600
rect 9263 12597 9275 12631
rect 10428 12628 10456 12872
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 11238 12832 11244 12844
rect 11199 12804 11244 12832
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11606 12792 11612 12844
rect 11664 12832 11670 12844
rect 12912 12841 12940 12940
rect 12986 12928 12992 12980
rect 13044 12968 13050 12980
rect 13449 12971 13507 12977
rect 13449 12968 13461 12971
rect 13044 12940 13461 12968
rect 13044 12928 13050 12940
rect 13449 12937 13461 12940
rect 13495 12937 13507 12971
rect 13449 12931 13507 12937
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11664 12804 11805 12832
rect 11664 12792 11670 12804
rect 11793 12801 11805 12804
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 13464 12832 13492 12931
rect 13538 12928 13544 12980
rect 13596 12968 13602 12980
rect 14093 12971 14151 12977
rect 14093 12968 14105 12971
rect 13596 12940 14105 12968
rect 13596 12928 13602 12940
rect 14093 12937 14105 12940
rect 14139 12937 14151 12971
rect 14093 12931 14151 12937
rect 15473 12971 15531 12977
rect 15473 12937 15485 12971
rect 15519 12968 15531 12971
rect 15746 12968 15752 12980
rect 15519 12940 15752 12968
rect 15519 12937 15531 12940
rect 15473 12931 15531 12937
rect 15746 12928 15752 12940
rect 15804 12968 15810 12980
rect 16022 12968 16028 12980
rect 15804 12940 16028 12968
rect 15804 12928 15810 12940
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 16482 12968 16488 12980
rect 16443 12940 16488 12968
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 17494 12968 17500 12980
rect 17455 12940 17500 12968
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 19426 12968 19432 12980
rect 19387 12940 19432 12968
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19518 12928 19524 12980
rect 19576 12968 19582 12980
rect 19705 12971 19763 12977
rect 19705 12968 19717 12971
rect 19576 12940 19717 12968
rect 19576 12928 19582 12940
rect 19705 12937 19717 12940
rect 19751 12968 19763 12971
rect 19797 12971 19855 12977
rect 19797 12968 19809 12971
rect 19751 12940 19809 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 19797 12937 19809 12940
rect 19843 12937 19855 12971
rect 19797 12931 19855 12937
rect 20714 12928 20720 12980
rect 20772 12968 20778 12980
rect 21637 12971 21695 12977
rect 21637 12968 21649 12971
rect 20772 12940 21649 12968
rect 20772 12928 20778 12940
rect 21637 12937 21649 12940
rect 21683 12937 21695 12971
rect 23750 12968 23756 12980
rect 23711 12940 23756 12968
rect 21637 12931 21695 12937
rect 23750 12928 23756 12940
rect 23808 12928 23814 12980
rect 24670 12968 24676 12980
rect 24320 12940 24676 12968
rect 13906 12900 13912 12912
rect 13867 12872 13912 12900
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 16301 12903 16359 12909
rect 16301 12869 16313 12903
rect 16347 12900 16359 12903
rect 17218 12900 17224 12912
rect 16347 12872 17224 12900
rect 16347 12869 16359 12872
rect 16301 12863 16359 12869
rect 17218 12860 17224 12872
rect 17276 12860 17282 12912
rect 18414 12860 18420 12912
rect 18472 12900 18478 12912
rect 18509 12903 18567 12909
rect 18509 12900 18521 12903
rect 18472 12872 18521 12900
rect 18472 12860 18478 12872
rect 18509 12869 18521 12872
rect 18555 12869 18567 12903
rect 18509 12863 18567 12869
rect 19150 12860 19156 12912
rect 19208 12900 19214 12912
rect 20073 12903 20131 12909
rect 20073 12900 20085 12903
rect 19208 12872 20085 12900
rect 19208 12860 19214 12872
rect 20073 12869 20085 12872
rect 20119 12869 20131 12903
rect 20073 12863 20131 12869
rect 21085 12903 21143 12909
rect 21085 12869 21097 12903
rect 21131 12900 21143 12903
rect 21174 12900 21180 12912
rect 21131 12872 21180 12900
rect 21131 12869 21143 12872
rect 21085 12863 21143 12869
rect 21174 12860 21180 12872
rect 21232 12860 21238 12912
rect 14461 12835 14519 12841
rect 14461 12832 14473 12835
rect 13464 12804 14473 12832
rect 12897 12795 12955 12801
rect 14461 12801 14473 12804
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 14550 12792 14556 12844
rect 14608 12832 14614 12844
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14608 12804 15117 12832
rect 14608 12792 14614 12804
rect 15105 12801 15117 12804
rect 15151 12832 15163 12835
rect 15654 12832 15660 12844
rect 15151 12804 15660 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 15654 12792 15660 12804
rect 15712 12832 15718 12844
rect 15933 12835 15991 12841
rect 15933 12832 15945 12835
rect 15712 12804 15945 12832
rect 15712 12792 15718 12804
rect 15933 12801 15945 12804
rect 15979 12832 15991 12835
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 15979 12804 17049 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 17037 12801 17049 12804
rect 17083 12832 17095 12835
rect 18322 12832 18328 12844
rect 17083 12804 18328 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12832 19119 12835
rect 19242 12832 19248 12844
rect 19107 12804 19248 12832
rect 19107 12801 19119 12804
rect 19061 12795 19119 12801
rect 10594 12764 10600 12776
rect 10555 12736 10600 12764
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 11422 12724 11428 12776
rect 11480 12764 11486 12776
rect 13538 12764 13544 12776
rect 11480 12736 11525 12764
rect 13004 12736 13544 12764
rect 11480 12724 11486 12736
rect 10502 12656 10508 12708
rect 10560 12696 10566 12708
rect 13004 12705 13032 12736
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 14332 12736 14657 12764
rect 14332 12724 14338 12736
rect 14645 12733 14657 12736
rect 14691 12733 14703 12767
rect 16758 12764 16764 12776
rect 16719 12736 16764 12764
rect 14645 12727 14703 12733
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 17862 12764 17868 12776
rect 17775 12736 17868 12764
rect 17862 12724 17868 12736
rect 17920 12764 17926 12776
rect 19076 12764 19104 12795
rect 19242 12792 19248 12804
rect 19300 12792 19306 12844
rect 20162 12792 20168 12844
rect 20220 12832 20226 12844
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20220 12804 20637 12832
rect 20220 12792 20226 12804
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12832 22247 12835
rect 22278 12832 22284 12844
rect 22235 12804 22284 12832
rect 22235 12801 22247 12804
rect 22189 12795 22247 12801
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 24320 12841 24348 12940
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 25409 12971 25467 12977
rect 25409 12937 25421 12971
rect 25455 12968 25467 12971
rect 25590 12968 25596 12980
rect 25455 12940 25596 12968
rect 25455 12937 25467 12940
rect 25409 12931 25467 12937
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 25038 12860 25044 12912
rect 25096 12900 25102 12912
rect 25777 12903 25835 12909
rect 25777 12900 25789 12903
rect 25096 12872 25789 12900
rect 25096 12860 25102 12872
rect 25777 12869 25789 12872
rect 25823 12869 25835 12903
rect 25777 12863 25835 12869
rect 24305 12835 24363 12841
rect 24305 12801 24317 12835
rect 24351 12801 24363 12835
rect 24305 12795 24363 12801
rect 17920 12736 19104 12764
rect 19705 12767 19763 12773
rect 17920 12724 17926 12736
rect 19705 12733 19717 12767
rect 19751 12764 19763 12767
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 19751 12736 20361 12764
rect 19751 12733 19763 12736
rect 19705 12727 19763 12733
rect 20349 12733 20361 12736
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 24210 12724 24216 12776
rect 24268 12764 24274 12776
rect 24670 12764 24676 12776
rect 24268 12736 24676 12764
rect 24268 12724 24274 12736
rect 24670 12724 24676 12736
rect 24728 12724 24734 12776
rect 25225 12767 25283 12773
rect 25225 12733 25237 12767
rect 25271 12764 25283 12767
rect 25498 12764 25504 12776
rect 25271 12736 25504 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 25498 12724 25504 12736
rect 25556 12764 25562 12776
rect 26145 12767 26203 12773
rect 26145 12764 26157 12767
rect 25556 12736 26157 12764
rect 25556 12724 25562 12736
rect 26145 12733 26157 12736
rect 26191 12733 26203 12767
rect 26145 12727 26203 12733
rect 11333 12699 11391 12705
rect 11333 12696 11345 12699
rect 10560 12668 11345 12696
rect 10560 12656 10566 12668
rect 11333 12665 11345 12668
rect 11379 12696 11391 12699
rect 12511 12699 12569 12705
rect 12511 12696 12523 12699
rect 11379 12668 12523 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 12511 12665 12523 12668
rect 12557 12665 12569 12699
rect 12511 12659 12569 12665
rect 12989 12699 13047 12705
rect 12989 12665 13001 12699
rect 13035 12665 13047 12699
rect 12989 12659 13047 12665
rect 13078 12656 13084 12708
rect 13136 12696 13142 12708
rect 13136 12668 13181 12696
rect 13136 12656 13142 12668
rect 13906 12656 13912 12708
rect 13964 12696 13970 12708
rect 14553 12699 14611 12705
rect 14553 12696 14565 12699
rect 13964 12668 14565 12696
rect 13964 12656 13970 12668
rect 14553 12665 14565 12668
rect 14599 12665 14611 12699
rect 14553 12659 14611 12665
rect 18046 12656 18052 12708
rect 18104 12696 18110 12708
rect 18325 12699 18383 12705
rect 18325 12696 18337 12699
rect 18104 12668 18337 12696
rect 18104 12656 18110 12668
rect 18325 12665 18337 12668
rect 18371 12696 18383 12699
rect 18785 12699 18843 12705
rect 18785 12696 18797 12699
rect 18371 12668 18797 12696
rect 18371 12665 18383 12668
rect 18325 12659 18383 12665
rect 18785 12665 18797 12668
rect 18831 12665 18843 12699
rect 19794 12696 19800 12708
rect 18785 12659 18843 12665
rect 19352 12668 19800 12696
rect 19352 12640 19380 12668
rect 19794 12656 19800 12668
rect 19852 12656 19858 12708
rect 21542 12656 21548 12708
rect 21600 12696 21606 12708
rect 21913 12699 21971 12705
rect 21913 12696 21925 12699
rect 21600 12668 21925 12696
rect 21600 12656 21606 12668
rect 21913 12665 21925 12668
rect 21959 12665 21971 12699
rect 24029 12699 24087 12705
rect 24029 12696 24041 12699
rect 21913 12659 21971 12665
rect 23308 12668 24041 12696
rect 23308 12640 23336 12668
rect 24029 12665 24041 12668
rect 24075 12665 24087 12699
rect 24029 12659 24087 12665
rect 11238 12628 11244 12640
rect 10428 12600 11244 12628
rect 9217 12591 9275 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 13538 12628 13544 12640
rect 13320 12600 13544 12628
rect 13320 12588 13326 12600
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 16945 12631 17003 12637
rect 16945 12628 16957 12631
rect 16632 12600 16957 12628
rect 16632 12588 16638 12600
rect 16945 12597 16957 12600
rect 16991 12597 17003 12631
rect 18966 12628 18972 12640
rect 18927 12600 18972 12628
rect 16945 12591 17003 12597
rect 18966 12588 18972 12600
rect 19024 12588 19030 12640
rect 19334 12588 19340 12640
rect 19392 12588 19398 12640
rect 20530 12628 20536 12640
rect 20491 12600 20536 12628
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 21358 12628 21364 12640
rect 21319 12600 21364 12628
rect 21358 12588 21364 12600
rect 21416 12628 21422 12640
rect 22097 12631 22155 12637
rect 22097 12628 22109 12631
rect 21416 12600 22109 12628
rect 21416 12588 21422 12600
rect 22097 12597 22109 12600
rect 22143 12597 22155 12631
rect 22646 12628 22652 12640
rect 22607 12600 22652 12628
rect 22097 12591 22155 12597
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 23109 12631 23167 12637
rect 23109 12597 23121 12631
rect 23155 12628 23167 12631
rect 23290 12628 23296 12640
rect 23155 12600 23296 12628
rect 23155 12597 23167 12600
rect 23109 12591 23167 12597
rect 23290 12588 23296 12600
rect 23348 12588 23354 12640
rect 23477 12631 23535 12637
rect 23477 12597 23489 12631
rect 23523 12628 23535 12631
rect 24210 12628 24216 12640
rect 23523 12600 24216 12628
rect 23523 12597 23535 12600
rect 23477 12591 23535 12597
rect 24210 12588 24216 12600
rect 24268 12588 24274 12640
rect 25038 12628 25044 12640
rect 24999 12600 25044 12628
rect 25038 12588 25044 12600
rect 25096 12588 25102 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1394 12424 1400 12436
rect 1355 12396 1400 12424
rect 1394 12384 1400 12396
rect 1452 12384 1458 12436
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2314 12424 2320 12436
rect 1995 12396 2320 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 3513 12427 3571 12433
rect 3513 12424 3525 12427
rect 3292 12396 3525 12424
rect 3292 12384 3298 12396
rect 3513 12393 3525 12396
rect 3559 12424 3571 12427
rect 3602 12424 3608 12436
rect 3559 12396 3608 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 3602 12384 3608 12396
rect 3660 12424 3666 12436
rect 4338 12424 4344 12436
rect 3660 12396 4344 12424
rect 3660 12384 3666 12396
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 5258 12424 5264 12436
rect 5219 12396 5264 12424
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 5721 12427 5779 12433
rect 5721 12393 5733 12427
rect 5767 12424 5779 12427
rect 5994 12424 6000 12436
rect 5767 12396 6000 12424
rect 5767 12393 5779 12396
rect 5721 12387 5779 12393
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 7193 12427 7251 12433
rect 7193 12393 7205 12427
rect 7239 12424 7251 12427
rect 7650 12424 7656 12436
rect 7239 12396 7656 12424
rect 7239 12393 7251 12396
rect 7193 12387 7251 12393
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 8662 12424 8668 12436
rect 8623 12396 8668 12424
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8904 12396 9045 12424
rect 8904 12384 8910 12396
rect 9033 12393 9045 12396
rect 9079 12424 9091 12427
rect 9309 12427 9367 12433
rect 9309 12424 9321 12427
rect 9079 12396 9321 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9309 12393 9321 12396
rect 9355 12393 9367 12427
rect 15654 12424 15660 12436
rect 15615 12396 15660 12424
rect 9309 12387 9367 12393
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 16482 12424 16488 12436
rect 15804 12396 16488 12424
rect 15804 12384 15810 12396
rect 16482 12384 16488 12396
rect 16540 12424 16546 12436
rect 17221 12427 17279 12433
rect 17221 12424 17233 12427
rect 16540 12396 17233 12424
rect 16540 12384 16546 12396
rect 17221 12393 17233 12396
rect 17267 12393 17279 12427
rect 18509 12427 18567 12433
rect 18509 12424 18521 12427
rect 17221 12387 17279 12393
rect 17604 12396 18521 12424
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2556 12328 2789 12356
rect 2556 12316 2562 12328
rect 2777 12325 2789 12328
rect 2823 12325 2835 12359
rect 2958 12356 2964 12368
rect 2919 12328 2964 12356
rect 2777 12319 2835 12325
rect 2958 12316 2964 12328
rect 3016 12316 3022 12368
rect 4614 12356 4620 12368
rect 4575 12328 4620 12356
rect 4614 12316 4620 12328
rect 4672 12316 4678 12368
rect 4798 12356 4804 12368
rect 4759 12328 4804 12356
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 4893 12359 4951 12365
rect 4893 12325 4905 12359
rect 4939 12356 4951 12359
rect 5534 12356 5540 12368
rect 4939 12328 5540 12356
rect 4939 12325 4951 12328
rect 4893 12319 4951 12325
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3326 12220 3332 12232
rect 3099 12192 3332 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3326 12180 3332 12192
rect 3384 12220 3390 12232
rect 4908 12220 4936 12319
rect 5534 12316 5540 12328
rect 5592 12316 5598 12368
rect 6365 12359 6423 12365
rect 6365 12325 6377 12359
rect 6411 12356 6423 12359
rect 6454 12356 6460 12368
rect 6411 12328 6460 12356
rect 6411 12325 6423 12328
rect 6365 12319 6423 12325
rect 5442 12248 5448 12300
rect 5500 12288 5506 12300
rect 5994 12288 6000 12300
rect 5500 12260 6000 12288
rect 5500 12248 5506 12260
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6178 12288 6184 12300
rect 6139 12260 6184 12288
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 6380 12288 6408 12319
rect 6454 12316 6460 12328
rect 6512 12316 6518 12368
rect 8202 12356 8208 12368
rect 8163 12328 8208 12356
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 9674 12356 9680 12368
rect 9635 12328 9680 12356
rect 9674 12316 9680 12328
rect 9732 12316 9738 12368
rect 12713 12359 12771 12365
rect 12713 12325 12725 12359
rect 12759 12356 12771 12359
rect 13722 12356 13728 12368
rect 12759 12328 13728 12356
rect 12759 12325 12771 12328
rect 12713 12319 12771 12325
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 15672 12356 15700 12384
rect 16086 12359 16144 12365
rect 16086 12356 16098 12359
rect 15672 12328 16098 12356
rect 16086 12325 16098 12328
rect 16132 12325 16144 12359
rect 16086 12319 16144 12325
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 17604 12356 17632 12396
rect 18509 12393 18521 12396
rect 18555 12424 18567 12427
rect 18966 12424 18972 12436
rect 18555 12396 18972 12424
rect 18555 12393 18567 12396
rect 18509 12387 18567 12393
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 20993 12427 21051 12433
rect 20993 12393 21005 12427
rect 21039 12424 21051 12427
rect 21082 12424 21088 12436
rect 21039 12396 21088 12424
rect 21039 12393 21051 12396
rect 20993 12387 21051 12393
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 22922 12384 22928 12436
rect 22980 12424 22986 12436
rect 23385 12427 23443 12433
rect 23385 12424 23397 12427
rect 22980 12396 23397 12424
rect 22980 12384 22986 12396
rect 23385 12393 23397 12396
rect 23431 12424 23443 12427
rect 23937 12427 23995 12433
rect 23937 12424 23949 12427
rect 23431 12396 23949 12424
rect 23431 12393 23443 12396
rect 23385 12387 23443 12393
rect 23937 12393 23949 12396
rect 23983 12393 23995 12427
rect 23937 12387 23995 12393
rect 16448 12328 17632 12356
rect 16448 12316 16454 12328
rect 18414 12316 18420 12368
rect 18472 12356 18478 12368
rect 19153 12359 19211 12365
rect 19153 12356 19165 12359
rect 18472 12328 19165 12356
rect 18472 12316 18478 12328
rect 19153 12325 19165 12328
rect 19199 12325 19211 12359
rect 20254 12356 20260 12368
rect 20215 12328 20260 12356
rect 19153 12319 19211 12325
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 20717 12359 20775 12365
rect 20717 12325 20729 12359
rect 20763 12356 20775 12359
rect 21450 12356 21456 12368
rect 20763 12328 21456 12356
rect 20763 12325 20775 12328
rect 20717 12319 20775 12325
rect 21450 12316 21456 12328
rect 21508 12316 21514 12368
rect 22646 12356 22652 12368
rect 22020 12328 22652 12356
rect 6288 12260 6408 12288
rect 3384 12192 4936 12220
rect 5537 12223 5595 12229
rect 3384 12180 3390 12192
rect 5537 12189 5549 12223
rect 5583 12220 5595 12223
rect 6288 12220 6316 12260
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 7374 12288 7380 12300
rect 6604 12260 7380 12288
rect 6604 12248 6610 12260
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 9030 12288 9036 12300
rect 8128 12260 9036 12288
rect 6454 12220 6460 12232
rect 5583 12192 6316 12220
rect 6415 12192 6460 12220
rect 5583 12189 5595 12192
rect 5537 12183 5595 12189
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 8128 12220 8156 12260
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 9950 12288 9956 12300
rect 9548 12260 9956 12288
rect 9548 12248 9554 12260
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10597 12291 10655 12297
rect 10597 12257 10609 12291
rect 10643 12288 10655 12291
rect 10778 12288 10784 12300
rect 10643 12260 10784 12288
rect 10643 12257 10655 12260
rect 10597 12251 10655 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 10956 12291 11014 12297
rect 10956 12257 10968 12291
rect 11002 12288 11014 12291
rect 11422 12288 11428 12300
rect 11002 12260 11428 12288
rect 11002 12257 11014 12260
rect 10956 12251 11014 12257
rect 11422 12248 11428 12260
rect 11480 12248 11486 12300
rect 13078 12288 13084 12300
rect 12991 12260 13084 12288
rect 13078 12248 13084 12260
rect 13136 12288 13142 12300
rect 13136 12260 13860 12288
rect 13136 12248 13142 12260
rect 8294 12220 8300 12232
rect 7024 12192 8156 12220
rect 8255 12192 8300 12220
rect 2501 12155 2559 12161
rect 2501 12121 2513 12155
rect 2547 12152 2559 12155
rect 2682 12152 2688 12164
rect 2547 12124 2688 12152
rect 2547 12121 2559 12124
rect 2501 12115 2559 12121
rect 2682 12112 2688 12124
rect 2740 12112 2746 12164
rect 4341 12155 4399 12161
rect 4341 12121 4353 12155
rect 4387 12152 4399 12155
rect 4430 12152 4436 12164
rect 4387 12124 4436 12152
rect 4387 12121 4399 12124
rect 4341 12115 4399 12121
rect 4430 12112 4436 12124
rect 4488 12112 4494 12164
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 7024 12152 7052 12192
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 10502 12180 10508 12232
rect 10560 12220 10566 12232
rect 10689 12223 10747 12229
rect 10689 12220 10701 12223
rect 10560 12192 10701 12220
rect 10560 12180 10566 12192
rect 10689 12189 10701 12192
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12250 12220 12256 12232
rect 12124 12192 12256 12220
rect 12124 12180 12130 12192
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 13722 12220 13728 12232
rect 13683 12192 13728 12220
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 13832 12229 13860 12260
rect 14458 12248 14464 12300
rect 14516 12288 14522 12300
rect 18046 12288 18052 12300
rect 14516 12260 18052 12288
rect 14516 12248 14522 12260
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 22020 12297 22048 12328
rect 22646 12316 22652 12328
rect 22704 12316 22710 12368
rect 25041 12359 25099 12365
rect 25041 12325 25053 12359
rect 25087 12356 25099 12359
rect 25498 12356 25504 12368
rect 25087 12328 25504 12356
rect 25087 12325 25099 12328
rect 25041 12319 25099 12325
rect 25498 12316 25504 12328
rect 25556 12316 25562 12368
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 18748 12260 19257 12288
rect 18748 12248 18754 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 22005 12291 22063 12297
rect 22005 12257 22017 12291
rect 22051 12257 22063 12291
rect 22272 12291 22330 12297
rect 22272 12288 22284 12291
rect 22005 12251 22063 12257
rect 22112 12260 22284 12288
rect 13817 12223 13875 12229
rect 13817 12189 13829 12223
rect 13863 12220 13875 12223
rect 13998 12220 14004 12232
rect 13863 12192 14004 12220
rect 13863 12189 13875 12192
rect 13817 12183 13875 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14918 12220 14924 12232
rect 14879 12192 14924 12220
rect 14918 12180 14924 12192
rect 14976 12180 14982 12232
rect 15838 12220 15844 12232
rect 15799 12192 15844 12220
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 19150 12220 19156 12232
rect 19111 12192 19156 12220
rect 19150 12180 19156 12192
rect 19208 12180 19214 12232
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 22112 12220 22140 12260
rect 22272 12257 22284 12260
rect 22318 12288 22330 12291
rect 22554 12288 22560 12300
rect 22318 12260 22560 12288
rect 22318 12257 22330 12260
rect 22272 12251 22330 12257
rect 22554 12248 22560 12260
rect 22612 12248 22618 12300
rect 23382 12248 23388 12300
rect 23440 12288 23446 12300
rect 23842 12288 23848 12300
rect 23440 12260 23848 12288
rect 23440 12248 23446 12260
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 24302 12220 24308 12232
rect 20772 12192 22140 12220
rect 24263 12192 24308 12220
rect 20772 12180 20778 12192
rect 24302 12180 24308 12192
rect 24360 12180 24366 12232
rect 24946 12220 24952 12232
rect 24907 12192 24952 12220
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 25133 12223 25191 12229
rect 25133 12189 25145 12223
rect 25179 12220 25191 12223
rect 25222 12220 25228 12232
rect 25179 12192 25228 12220
rect 25179 12189 25191 12192
rect 25133 12183 25191 12189
rect 25222 12180 25228 12192
rect 25280 12180 25286 12232
rect 4672 12124 7052 12152
rect 4672 12112 4678 12124
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 8720 12124 9413 12152
rect 8720 12112 8726 12124
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 13740 12152 13768 12180
rect 14553 12155 14611 12161
rect 14553 12152 14565 12155
rect 13740 12124 14565 12152
rect 9401 12115 9459 12121
rect 14553 12121 14565 12124
rect 14599 12121 14611 12155
rect 14553 12115 14611 12121
rect 18966 12112 18972 12164
rect 19024 12152 19030 12164
rect 21358 12152 21364 12164
rect 19024 12124 21364 12152
rect 19024 12112 19030 12124
rect 21358 12112 21364 12124
rect 21416 12112 21422 12164
rect 24964 12152 24992 12180
rect 25501 12155 25559 12161
rect 25501 12152 25513 12155
rect 24964 12124 25513 12152
rect 25501 12121 25513 12124
rect 25547 12121 25559 12155
rect 25501 12115 25559 12121
rect 3786 12084 3792 12096
rect 3747 12056 3792 12084
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 5537 12087 5595 12093
rect 5537 12084 5549 12087
rect 5500 12056 5549 12084
rect 5500 12044 5506 12056
rect 5537 12053 5549 12056
rect 5583 12053 5595 12087
rect 5537 12047 5595 12053
rect 5905 12087 5963 12093
rect 5905 12053 5917 12087
rect 5951 12084 5963 12087
rect 6546 12084 6552 12096
rect 5951 12056 6552 12084
rect 5951 12053 5963 12056
rect 5905 12047 5963 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 7561 12087 7619 12093
rect 7561 12084 7573 12087
rect 7248 12056 7573 12084
rect 7248 12044 7254 12056
rect 7561 12053 7573 12056
rect 7607 12084 7619 12087
rect 7650 12084 7656 12096
rect 7607 12056 7656 12084
rect 7607 12053 7619 12056
rect 7561 12047 7619 12053
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12084 7803 12087
rect 7834 12084 7840 12096
rect 7791 12056 7840 12084
rect 7791 12053 7803 12056
rect 7745 12047 7803 12053
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 9309 12087 9367 12093
rect 9309 12053 9321 12087
rect 9355 12084 9367 12087
rect 9490 12084 9496 12096
rect 9355 12056 9496 12084
rect 9355 12053 9367 12056
rect 9309 12047 9367 12053
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 10229 12087 10287 12093
rect 10229 12053 10241 12087
rect 10275 12084 10287 12087
rect 10686 12084 10692 12096
rect 10275 12056 10692 12084
rect 10275 12053 10287 12056
rect 10229 12047 10287 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 12066 12084 12072 12096
rect 12027 12056 12072 12084
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 13136 12056 13277 12084
rect 13136 12044 13142 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 14274 12084 14280 12096
rect 14235 12056 14280 12084
rect 13265 12047 13323 12053
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 17770 12084 17776 12096
rect 17731 12056 17776 12084
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 18693 12087 18751 12093
rect 18693 12053 18705 12087
rect 18739 12084 18751 12087
rect 19242 12084 19248 12096
rect 18739 12056 19248 12084
rect 18739 12053 18751 12056
rect 18693 12047 18751 12053
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 19981 12087 20039 12093
rect 19981 12053 19993 12087
rect 20027 12084 20039 12087
rect 20622 12084 20628 12096
rect 20027 12056 20628 12084
rect 20027 12053 20039 12056
rect 19981 12047 20039 12053
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 21542 12084 21548 12096
rect 21503 12056 21548 12084
rect 21542 12044 21548 12056
rect 21600 12044 21606 12096
rect 23750 12044 23756 12096
rect 23808 12084 23814 12096
rect 24581 12087 24639 12093
rect 24581 12084 24593 12087
rect 23808 12056 24593 12084
rect 23808 12044 23814 12056
rect 24581 12053 24593 12056
rect 24627 12053 24639 12087
rect 24581 12047 24639 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 2832 11852 2877 11880
rect 2832 11840 2838 11852
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 4488 11852 5641 11880
rect 4488 11840 4494 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 6362 11880 6368 11892
rect 6323 11852 6368 11880
rect 5629 11843 5687 11849
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 8202 11880 8208 11892
rect 7248 11852 8208 11880
rect 7248 11840 7254 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8478 11880 8484 11892
rect 8439 11852 8484 11880
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9582 11880 9588 11892
rect 9180 11852 9588 11880
rect 9180 11840 9186 11852
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 10134 11840 10140 11892
rect 10192 11840 10198 11892
rect 10502 11880 10508 11892
rect 10415 11852 10508 11880
rect 10502 11840 10508 11852
rect 10560 11880 10566 11892
rect 11330 11880 11336 11892
rect 10560 11852 11336 11880
rect 10560 11840 10566 11852
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 13998 11840 14004 11892
rect 14056 11880 14062 11892
rect 15197 11883 15255 11889
rect 15197 11880 15209 11883
rect 14056 11852 15209 11880
rect 14056 11840 14062 11852
rect 15197 11849 15209 11852
rect 15243 11849 15255 11883
rect 19426 11880 19432 11892
rect 19387 11852 19432 11880
rect 15197 11843 15255 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 21545 11883 21603 11889
rect 21545 11849 21557 11883
rect 21591 11880 21603 11883
rect 21634 11880 21640 11892
rect 21591 11852 21640 11880
rect 21591 11849 21603 11852
rect 21545 11843 21603 11849
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 22557 11883 22615 11889
rect 22557 11849 22569 11883
rect 22603 11880 22615 11883
rect 22646 11880 22652 11892
rect 22603 11852 22652 11880
rect 22603 11849 22615 11852
rect 22557 11843 22615 11849
rect 22646 11840 22652 11852
rect 22704 11880 22710 11892
rect 25038 11880 25044 11892
rect 22704 11852 23520 11880
rect 24951 11852 25044 11880
rect 22704 11840 22710 11852
rect 2590 11772 2596 11824
rect 2648 11812 2654 11824
rect 4157 11815 4215 11821
rect 4157 11812 4169 11815
rect 2648 11784 4169 11812
rect 2648 11772 2654 11784
rect 4157 11781 4169 11784
rect 4203 11812 4215 11815
rect 4203 11784 4292 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 3237 11747 3295 11753
rect 3237 11744 3249 11747
rect 2832 11716 3249 11744
rect 2832 11704 2838 11716
rect 3237 11713 3249 11716
rect 3283 11744 3295 11747
rect 4062 11744 4068 11756
rect 3283 11716 4068 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 4264 11753 4292 11784
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 6181 11815 6239 11821
rect 6181 11812 6193 11815
rect 5500 11784 6193 11812
rect 5500 11772 5506 11784
rect 6181 11781 6193 11784
rect 6227 11781 6239 11815
rect 6181 11775 6239 11781
rect 6917 11815 6975 11821
rect 6917 11781 6929 11815
rect 6963 11812 6975 11815
rect 7006 11812 7012 11824
rect 6963 11784 7012 11812
rect 6963 11781 6975 11784
rect 6917 11775 6975 11781
rect 7006 11772 7012 11784
rect 7064 11772 7070 11824
rect 7098 11772 7104 11824
rect 7156 11812 7162 11824
rect 7834 11812 7840 11824
rect 7156 11784 7840 11812
rect 7156 11772 7162 11784
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 10152 11812 10180 11840
rect 10321 11815 10379 11821
rect 10321 11812 10333 11815
rect 8496 11784 10333 11812
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1578 11676 1584 11688
rect 1443 11648 1584 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1578 11636 1584 11648
rect 1636 11636 1642 11688
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11676 2559 11679
rect 3326 11676 3332 11688
rect 2547 11648 3332 11676
rect 2547 11645 2559 11648
rect 2501 11639 2559 11645
rect 3326 11636 3332 11648
rect 3384 11636 3390 11688
rect 4264 11676 4292 11707
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 8496 11744 8524 11784
rect 10321 11781 10333 11784
rect 10367 11781 10379 11815
rect 10686 11812 10692 11824
rect 10647 11784 10692 11812
rect 10321 11775 10379 11781
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 15378 11772 15384 11824
rect 15436 11812 15442 11824
rect 16393 11815 16451 11821
rect 16393 11812 16405 11815
rect 15436 11784 16405 11812
rect 15436 11772 15442 11784
rect 16393 11781 16405 11784
rect 16439 11781 16451 11815
rect 16393 11775 16451 11781
rect 18417 11815 18475 11821
rect 18417 11781 18429 11815
rect 18463 11812 18475 11815
rect 18782 11812 18788 11824
rect 18463 11784 18788 11812
rect 18463 11781 18475 11784
rect 18417 11775 18475 11781
rect 18782 11772 18788 11784
rect 18840 11772 18846 11824
rect 19978 11812 19984 11824
rect 19939 11784 19984 11812
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 20070 11772 20076 11824
rect 20128 11812 20134 11824
rect 23290 11812 23296 11824
rect 20128 11784 23296 11812
rect 20128 11772 20134 11784
rect 23290 11772 23296 11784
rect 23348 11772 23354 11824
rect 5316 11716 8524 11744
rect 8941 11747 8999 11753
rect 5316 11704 5322 11716
rect 8941 11713 8953 11747
rect 8987 11744 8999 11747
rect 9582 11744 9588 11756
rect 8987 11716 9588 11744
rect 8987 11713 8999 11716
rect 8941 11707 8999 11713
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 10134 11744 10140 11756
rect 10047 11716 10140 11744
rect 10134 11704 10140 11716
rect 10192 11744 10198 11756
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 10192 11716 11253 11744
rect 10192 11704 10198 11716
rect 11241 11713 11253 11716
rect 11287 11744 11299 11747
rect 11606 11744 11612 11756
rect 11287 11716 11612 11744
rect 11287 11713 11299 11716
rect 11241 11707 11299 11713
rect 11606 11704 11612 11716
rect 11664 11744 11670 11756
rect 12066 11744 12072 11756
rect 11664 11716 12072 11744
rect 11664 11704 11670 11716
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16298 11744 16304 11756
rect 15887 11716 16304 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16298 11704 16304 11716
rect 16356 11744 16362 11756
rect 16761 11747 16819 11753
rect 16761 11744 16773 11747
rect 16356 11716 16773 11744
rect 16356 11704 16362 11716
rect 16761 11713 16773 11716
rect 16807 11713 16819 11747
rect 16761 11707 16819 11713
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11744 18935 11747
rect 19058 11744 19064 11756
rect 18923 11716 19064 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 19058 11704 19064 11716
rect 19116 11704 19122 11756
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11744 22155 11747
rect 22278 11744 22284 11756
rect 22143 11716 22284 11744
rect 22143 11713 22155 11716
rect 22097 11707 22155 11713
rect 22278 11704 22284 11716
rect 22336 11704 22342 11756
rect 22738 11704 22744 11756
rect 22796 11744 22802 11756
rect 23492 11753 23520 11852
rect 25038 11840 25044 11852
rect 25096 11880 25102 11892
rect 25958 11880 25964 11892
rect 25096 11852 25964 11880
rect 25096 11840 25102 11852
rect 25958 11840 25964 11852
rect 26016 11840 26022 11892
rect 23477 11747 23535 11753
rect 22796 11716 23336 11744
rect 22796 11704 22802 11716
rect 4338 11676 4344 11688
rect 4264 11648 4344 11676
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 6454 11636 6460 11688
rect 6512 11676 6518 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 6512 11648 7481 11676
rect 6512 11636 6518 11648
rect 7469 11645 7481 11648
rect 7515 11676 7527 11679
rect 7837 11679 7895 11685
rect 7837 11676 7849 11679
rect 7515 11648 7849 11676
rect 7515 11645 7527 11648
rect 7469 11639 7527 11645
rect 7837 11645 7849 11648
rect 7883 11676 7895 11679
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 7883 11648 8217 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 8205 11645 8217 11648
rect 8251 11676 8263 11679
rect 8294 11676 8300 11688
rect 8251 11648 8300 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 8294 11636 8300 11648
rect 8352 11676 8358 11688
rect 9033 11679 9091 11685
rect 9033 11676 9045 11679
rect 8352 11648 9045 11676
rect 8352 11636 8358 11648
rect 9033 11645 9045 11648
rect 9079 11676 9091 11679
rect 9214 11676 9220 11688
rect 9079 11648 9220 11676
rect 9079 11645 9091 11648
rect 9033 11639 9091 11645
rect 9214 11636 9220 11648
rect 9272 11676 9278 11688
rect 9401 11679 9459 11685
rect 9401 11676 9413 11679
rect 9272 11648 9413 11676
rect 9272 11636 9278 11648
rect 9401 11645 9413 11648
rect 9447 11645 9459 11679
rect 9401 11639 9459 11645
rect 10870 11636 10876 11688
rect 10928 11676 10934 11688
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 10928 11648 10977 11676
rect 10928 11636 10934 11648
rect 10965 11645 10977 11648
rect 11011 11645 11023 11679
rect 12713 11679 12771 11685
rect 12713 11676 12725 11679
rect 10965 11639 11023 11645
rect 12176 11648 12725 11676
rect 1670 11608 1676 11620
rect 1631 11580 1676 11608
rect 1670 11568 1676 11580
rect 1728 11568 1734 11620
rect 3237 11611 3295 11617
rect 3237 11577 3249 11611
rect 3283 11608 3295 11611
rect 3418 11608 3424 11620
rect 3283 11580 3424 11608
rect 3283 11577 3295 11580
rect 3237 11571 3295 11577
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 3789 11611 3847 11617
rect 3789 11577 3801 11611
rect 3835 11608 3847 11611
rect 4494 11611 4552 11617
rect 4494 11608 4506 11611
rect 3835 11580 4506 11608
rect 3835 11577 3847 11580
rect 3789 11571 3847 11577
rect 4494 11577 4506 11580
rect 4540 11608 4552 11611
rect 5442 11608 5448 11620
rect 4540 11580 5448 11608
rect 4540 11577 4552 11580
rect 4494 11571 4552 11577
rect 5442 11568 5448 11580
rect 5500 11568 5506 11620
rect 7193 11611 7251 11617
rect 7193 11608 7205 11611
rect 6840 11580 7205 11608
rect 6840 11552 6868 11580
rect 7193 11577 7205 11580
rect 7239 11577 7251 11611
rect 8938 11608 8944 11620
rect 8899 11580 8944 11608
rect 7193 11571 7251 11577
rect 8938 11568 8944 11580
rect 8996 11568 9002 11620
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 11149 11611 11207 11617
rect 11149 11608 11161 11611
rect 11112 11580 11161 11608
rect 11112 11568 11118 11580
rect 11149 11577 11161 11580
rect 11195 11577 11207 11611
rect 11149 11571 11207 11577
rect 11422 11568 11428 11620
rect 11480 11608 11486 11620
rect 11701 11611 11759 11617
rect 11701 11608 11713 11611
rect 11480 11580 11713 11608
rect 11480 11568 11486 11580
rect 11701 11577 11713 11580
rect 11747 11608 11759 11611
rect 11974 11608 11980 11620
rect 11747 11580 11980 11608
rect 11747 11577 11759 11580
rect 11701 11571 11759 11577
rect 11974 11568 11980 11580
rect 12032 11568 12038 11620
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 6328 11512 6377 11540
rect 6328 11500 6334 11512
rect 6365 11509 6377 11512
rect 6411 11509 6423 11543
rect 6365 11503 6423 11509
rect 6641 11543 6699 11549
rect 6641 11509 6653 11543
rect 6687 11540 6699 11543
rect 6822 11540 6828 11552
rect 6687 11512 6828 11540
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 6972 11512 7389 11540
rect 6972 11500 6978 11512
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 7377 11503 7435 11509
rect 10321 11543 10379 11549
rect 10321 11509 10333 11543
rect 10367 11540 10379 11543
rect 10870 11540 10876 11552
rect 10367 11512 10876 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 12176 11549 12204 11648
rect 12713 11645 12725 11648
rect 12759 11645 12771 11679
rect 12713 11639 12771 11645
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13228 11648 13737 11676
rect 13228 11636 13234 11648
rect 13725 11645 13737 11648
rect 13771 11676 13783 11679
rect 13817 11679 13875 11685
rect 13817 11676 13829 11679
rect 13771 11648 13829 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 13817 11645 13829 11648
rect 13863 11676 13875 11679
rect 15746 11676 15752 11688
rect 13863 11648 15752 11676
rect 13863 11645 13875 11648
rect 13817 11639 13875 11645
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 17865 11679 17923 11685
rect 17865 11645 17877 11679
rect 17911 11676 17923 11679
rect 18690 11676 18696 11688
rect 17911 11648 18696 11676
rect 17911 11645 17923 11648
rect 17865 11639 17923 11645
rect 18690 11636 18696 11648
rect 18748 11676 18754 11688
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18748 11648 18981 11676
rect 18748 11636 18754 11648
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 20533 11679 20591 11685
rect 20533 11676 20545 11679
rect 19484 11648 20545 11676
rect 19484 11636 19490 11648
rect 20533 11645 20545 11648
rect 20579 11645 20591 11679
rect 20533 11639 20591 11645
rect 20993 11679 21051 11685
rect 20993 11645 21005 11679
rect 21039 11676 21051 11679
rect 21266 11676 21272 11688
rect 21039 11648 21272 11676
rect 21039 11645 21051 11648
rect 20993 11639 21051 11645
rect 13357 11611 13415 11617
rect 13357 11577 13369 11611
rect 13403 11608 13415 11611
rect 14084 11611 14142 11617
rect 14084 11608 14096 11611
rect 13403 11580 14096 11608
rect 13403 11577 13415 11580
rect 13357 11571 13415 11577
rect 14084 11577 14096 11580
rect 14130 11608 14142 11611
rect 14274 11608 14280 11620
rect 14130 11580 14280 11608
rect 14130 11577 14142 11580
rect 14084 11571 14142 11577
rect 14274 11568 14280 11580
rect 14332 11608 14338 11620
rect 14550 11608 14556 11620
rect 14332 11580 14556 11608
rect 14332 11568 14338 11580
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 15562 11568 15568 11620
rect 15620 11608 15626 11620
rect 15620 11580 16252 11608
rect 15620 11568 15626 11580
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11848 11512 12173 11540
rect 11848 11500 11854 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 16224 11549 16252 11580
rect 16666 11568 16672 11620
rect 16724 11608 16730 11620
rect 16945 11611 17003 11617
rect 16945 11608 16957 11611
rect 16724 11580 16957 11608
rect 16724 11568 16730 11580
rect 16945 11577 16957 11580
rect 16991 11608 17003 11611
rect 17313 11611 17371 11617
rect 17313 11608 17325 11611
rect 16991 11580 17325 11608
rect 16991 11577 17003 11580
rect 16945 11571 17003 11577
rect 17313 11577 17325 11580
rect 17359 11577 17371 11611
rect 18874 11608 18880 11620
rect 18835 11580 18880 11608
rect 17313 11571 17371 11577
rect 18874 11568 18880 11580
rect 18932 11568 18938 11620
rect 20257 11611 20315 11617
rect 20257 11608 20269 11611
rect 19720 11580 20269 11608
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12860 11512 12909 11540
rect 12860 11500 12866 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 12897 11503 12955 11509
rect 16209 11543 16267 11549
rect 16209 11509 16221 11543
rect 16255 11540 16267 11543
rect 16850 11540 16856 11552
rect 16255 11512 16856 11540
rect 16255 11509 16267 11512
rect 16209 11503 16267 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 19720 11549 19748 11580
rect 20257 11577 20269 11580
rect 20303 11608 20315 11611
rect 20346 11608 20352 11620
rect 20303 11580 20352 11608
rect 20303 11577 20315 11580
rect 20257 11571 20315 11577
rect 20346 11568 20352 11580
rect 20404 11568 20410 11620
rect 20441 11611 20499 11617
rect 20441 11577 20453 11611
rect 20487 11608 20499 11611
rect 20622 11608 20628 11620
rect 20487 11580 20628 11608
rect 20487 11577 20499 11580
rect 20441 11571 20499 11577
rect 20622 11568 20628 11580
rect 20680 11608 20686 11620
rect 21008 11608 21036 11639
rect 21266 11636 21272 11648
rect 21324 11676 21330 11688
rect 23308 11676 23336 11716
rect 23477 11713 23489 11747
rect 23523 11744 23535 11747
rect 23661 11747 23719 11753
rect 23661 11744 23673 11747
rect 23523 11716 23673 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 23661 11713 23673 11716
rect 23707 11713 23719 11747
rect 23661 11707 23719 11713
rect 25590 11676 25596 11688
rect 21324 11648 22048 11676
rect 23308 11648 25360 11676
rect 25551 11648 25596 11676
rect 21324 11636 21330 11648
rect 22020 11620 22048 11648
rect 20680 11580 21036 11608
rect 21821 11611 21879 11617
rect 20680 11568 20686 11580
rect 21821 11577 21833 11611
rect 21867 11577 21879 11611
rect 22002 11608 22008 11620
rect 21963 11580 22008 11608
rect 21821 11571 21879 11577
rect 19705 11543 19763 11549
rect 19705 11540 19717 11543
rect 19392 11512 19717 11540
rect 19392 11500 19398 11512
rect 19705 11509 19717 11512
rect 19751 11509 19763 11543
rect 19705 11503 19763 11509
rect 20162 11500 20168 11552
rect 20220 11540 20226 11552
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 20220 11512 21281 11540
rect 20220 11500 20226 11512
rect 21269 11509 21281 11512
rect 21315 11540 21327 11543
rect 21836 11540 21864 11571
rect 22002 11568 22008 11580
rect 22060 11568 22066 11620
rect 23109 11611 23167 11617
rect 23109 11577 23121 11611
rect 23155 11608 23167 11611
rect 23928 11611 23986 11617
rect 23928 11608 23940 11611
rect 23155 11580 23940 11608
rect 23155 11577 23167 11580
rect 23109 11571 23167 11577
rect 23928 11577 23940 11580
rect 23974 11608 23986 11611
rect 24762 11608 24768 11620
rect 23974 11580 24768 11608
rect 23974 11577 23986 11580
rect 23928 11571 23986 11577
rect 24762 11568 24768 11580
rect 24820 11568 24826 11620
rect 25332 11608 25360 11648
rect 25590 11636 25596 11648
rect 25648 11636 25654 11688
rect 26326 11608 26332 11620
rect 25332 11580 26332 11608
rect 26326 11568 26332 11580
rect 26384 11568 26390 11620
rect 21315 11512 21864 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 25961 11543 26019 11549
rect 25961 11540 25973 11543
rect 25556 11512 25973 11540
rect 25556 11500 25562 11512
rect 25961 11509 25973 11512
rect 26007 11509 26019 11543
rect 25961 11503 26019 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1394 11336 1400 11348
rect 1355 11308 1400 11336
rect 1394 11296 1400 11308
rect 1452 11296 1458 11348
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2314 11336 2320 11348
rect 1995 11308 2320 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2314 11296 2320 11308
rect 2372 11336 2378 11348
rect 3234 11336 3240 11348
rect 2372 11308 3240 11336
rect 2372 11296 2378 11308
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 3326 11296 3332 11348
rect 3384 11336 3390 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3384 11308 3433 11336
rect 3384 11296 3390 11308
rect 3421 11305 3433 11308
rect 3467 11336 3479 11339
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3467 11308 3801 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 4338 11296 4344 11348
rect 4396 11296 4402 11348
rect 5902 11296 5908 11348
rect 5960 11336 5966 11348
rect 5997 11339 6055 11345
rect 5997 11336 6009 11339
rect 5960 11308 6009 11336
rect 5960 11296 5966 11308
rect 5997 11305 6009 11308
rect 6043 11336 6055 11339
rect 6178 11336 6184 11348
rect 6043 11308 6184 11336
rect 6043 11305 6055 11308
rect 5997 11299 6055 11305
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7616 11308 7757 11336
rect 7616 11296 7622 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 7745 11299 7803 11305
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11882 11336 11888 11348
rect 11112 11308 11888 11336
rect 11112 11296 11118 11308
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 13170 11336 13176 11348
rect 12728 11308 13176 11336
rect 2958 11268 2964 11280
rect 2919 11240 2964 11268
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 3053 11271 3111 11277
rect 3053 11237 3065 11271
rect 3099 11268 3111 11271
rect 3344 11268 3372 11296
rect 4356 11268 4384 11296
rect 7098 11268 7104 11280
rect 3099 11240 3372 11268
rect 4080 11240 4384 11268
rect 7059 11240 7104 11268
rect 3099 11237 3111 11240
rect 3053 11231 3111 11237
rect 3234 11160 3240 11212
rect 3292 11200 3298 11212
rect 4080 11209 4108 11240
rect 7098 11228 7104 11240
rect 7156 11228 7162 11280
rect 8478 11268 8484 11280
rect 8005 11240 8484 11268
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3292 11172 4077 11200
rect 3292 11160 3298 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4332 11203 4390 11209
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 4798 11200 4804 11212
rect 4378 11172 4804 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 8005 11200 8033 11240
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 10134 11228 10140 11280
rect 10192 11268 10198 11280
rect 10290 11271 10348 11277
rect 10290 11268 10302 11271
rect 10192 11240 10302 11268
rect 10192 11228 10198 11240
rect 10290 11237 10302 11240
rect 10336 11237 10348 11271
rect 10290 11231 10348 11237
rect 10962 11228 10968 11280
rect 11020 11268 11026 11280
rect 12618 11268 12624 11280
rect 11020 11240 12624 11268
rect 11020 11228 11026 11240
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 8110 11200 8116 11212
rect 6963 11172 8033 11200
rect 8071 11172 8116 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 8110 11160 8116 11172
rect 8168 11160 8174 11212
rect 8754 11200 8760 11212
rect 8404 11172 8760 11200
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3050 11132 3056 11144
rect 3007 11104 3056 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3050 11092 3056 11104
rect 3108 11132 3114 11144
rect 3326 11132 3332 11144
rect 3108 11104 3332 11132
rect 3108 11092 3114 11104
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 6546 11132 6552 11144
rect 5552 11104 6552 11132
rect 2406 11024 2412 11076
rect 2464 11064 2470 11076
rect 2501 11067 2559 11073
rect 2501 11064 2513 11067
rect 2464 11036 2513 11064
rect 2464 11024 2470 11036
rect 2501 11033 2513 11036
rect 2547 11033 2559 11067
rect 5442 11064 5448 11076
rect 5403 11036 5448 11064
rect 2501 11027 2559 11033
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 5166 10956 5172 11008
rect 5224 10996 5230 11008
rect 5552 10996 5580 11104
rect 6546 11092 6552 11104
rect 6604 11092 6610 11144
rect 7190 11132 7196 11144
rect 7151 11104 7196 11132
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 8294 11132 8300 11144
rect 8255 11104 8300 11132
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 6638 11064 6644 11076
rect 6599 11036 6644 11064
rect 6638 11024 6644 11036
rect 6696 11024 6702 11076
rect 6454 10996 6460 11008
rect 5224 10968 5580 10996
rect 6367 10968 6460 10996
rect 5224 10956 5230 10968
rect 6454 10956 6460 10968
rect 6512 10996 6518 11008
rect 6914 10996 6920 11008
rect 6512 10968 6920 10996
rect 6512 10956 6518 10968
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8404 10996 8432 11172
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 10045 11203 10103 11209
rect 10045 11169 10057 11203
rect 10091 11200 10103 11203
rect 11330 11200 11336 11212
rect 10091 11172 11336 11200
rect 10091 11169 10103 11172
rect 10045 11163 10103 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11200 12587 11203
rect 12728 11200 12756 11308
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 15838 11336 15844 11348
rect 15799 11308 15844 11336
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 18417 11339 18475 11345
rect 18417 11305 18429 11339
rect 18463 11336 18475 11339
rect 19058 11336 19064 11348
rect 18463 11308 19064 11336
rect 18463 11305 18475 11308
rect 18417 11299 18475 11305
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 20165 11339 20223 11345
rect 20165 11336 20177 11339
rect 19628 11308 20177 11336
rect 12796 11271 12854 11277
rect 12796 11237 12808 11271
rect 12842 11268 12854 11271
rect 12986 11268 12992 11280
rect 12842 11240 12992 11268
rect 12842 11237 12854 11240
rect 12796 11231 12854 11237
rect 12986 11228 12992 11240
rect 13044 11228 13050 11280
rect 12575 11172 12756 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 13078 11160 13084 11212
rect 13136 11200 13142 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 13136 11172 15025 11200
rect 13136 11160 13142 11172
rect 15013 11169 15025 11172
rect 15059 11169 15071 11203
rect 15856 11200 15884 11296
rect 16482 11277 16488 11280
rect 16476 11268 16488 11277
rect 16443 11240 16488 11268
rect 16476 11231 16488 11240
rect 16482 11228 16488 11231
rect 16540 11228 16546 11280
rect 18690 11268 18696 11280
rect 18651 11240 18696 11268
rect 18690 11228 18696 11240
rect 18748 11268 18754 11280
rect 19628 11268 19656 11308
rect 20165 11305 20177 11308
rect 20211 11305 20223 11339
rect 20714 11336 20720 11348
rect 20675 11308 20720 11336
rect 20165 11299 20223 11305
rect 18748 11240 19656 11268
rect 18748 11228 18754 11240
rect 19702 11228 19708 11280
rect 19760 11268 19766 11280
rect 20180 11268 20208 11299
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 21453 11339 21511 11345
rect 21453 11305 21465 11339
rect 21499 11336 21511 11339
rect 21634 11336 21640 11348
rect 21499 11308 21640 11336
rect 21499 11305 21511 11308
rect 21453 11299 21511 11305
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 22278 11336 22284 11348
rect 22239 11308 22284 11336
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22388 11308 23152 11336
rect 20622 11268 20628 11280
rect 19760 11240 19805 11268
rect 20180 11240 20628 11268
rect 19760 11228 19766 11240
rect 20622 11228 20628 11240
rect 20680 11268 20686 11280
rect 21913 11271 21971 11277
rect 21913 11268 21925 11271
rect 20680 11240 21925 11268
rect 20680 11228 20686 11240
rect 21913 11237 21925 11240
rect 21959 11237 21971 11271
rect 21913 11231 21971 11237
rect 22002 11228 22008 11280
rect 22060 11268 22066 11280
rect 22388 11268 22416 11308
rect 22830 11268 22836 11280
rect 22060 11240 22416 11268
rect 22791 11240 22836 11268
rect 22060 11228 22066 11240
rect 22830 11228 22836 11240
rect 22888 11228 22894 11280
rect 23014 11268 23020 11280
rect 22975 11240 23020 11268
rect 23014 11228 23020 11240
rect 23072 11228 23078 11280
rect 23124 11268 23152 11308
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 24578 11336 24584 11348
rect 23532 11308 24584 11336
rect 23532 11296 23538 11308
rect 24578 11296 24584 11308
rect 24636 11336 24642 11348
rect 24636 11308 25176 11336
rect 24636 11296 24642 11308
rect 24673 11271 24731 11277
rect 23124 11240 24532 11268
rect 16209 11203 16267 11209
rect 16209 11200 16221 11203
rect 15856 11172 16221 11200
rect 15013 11163 15071 11169
rect 16209 11169 16221 11172
rect 16255 11169 16267 11203
rect 16209 11163 16267 11169
rect 19426 11160 19432 11212
rect 19484 11200 19490 11212
rect 19797 11203 19855 11209
rect 19797 11200 19809 11203
rect 19484 11172 19809 11200
rect 19484 11160 19490 11172
rect 19797 11169 19809 11172
rect 19843 11200 19855 11203
rect 21545 11203 21603 11209
rect 21545 11200 21557 11203
rect 19843 11172 21557 11200
rect 19843 11169 19855 11172
rect 19797 11163 19855 11169
rect 21545 11169 21557 11172
rect 21591 11169 21603 11203
rect 23474 11200 23480 11212
rect 21545 11163 21603 11169
rect 21652 11172 23480 11200
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 8536 11104 9229 11132
rect 8536 11092 8542 11104
rect 9217 11101 9229 11104
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 15470 11132 15476 11144
rect 12492 11104 12537 11132
rect 15431 11104 15476 11132
rect 12492 11092 12498 11104
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 18564 11104 19717 11132
rect 18564 11092 18570 11104
rect 19705 11101 19717 11104
rect 19751 11132 19763 11135
rect 20346 11132 20352 11144
rect 19751 11104 20352 11132
rect 19751 11101 19763 11104
rect 19705 11095 19763 11101
rect 20346 11092 20352 11104
rect 20404 11092 20410 11144
rect 21450 11132 21456 11144
rect 21363 11104 21456 11132
rect 21450 11092 21456 11104
rect 21508 11132 21514 11144
rect 21652 11132 21680 11172
rect 23474 11160 23480 11172
rect 23532 11160 23538 11212
rect 24210 11160 24216 11212
rect 24268 11200 24274 11212
rect 24397 11203 24455 11209
rect 24397 11200 24409 11203
rect 24268 11172 24409 11200
rect 24268 11160 24274 11172
rect 24397 11169 24409 11172
rect 24443 11169 24455 11203
rect 24504 11200 24532 11240
rect 24673 11237 24685 11271
rect 24719 11268 24731 11271
rect 24762 11268 24768 11280
rect 24719 11240 24768 11268
rect 24719 11237 24731 11240
rect 24673 11231 24731 11237
rect 24762 11228 24768 11240
rect 24820 11228 24826 11280
rect 25148 11268 25176 11308
rect 25314 11296 25320 11348
rect 25372 11336 25378 11348
rect 25590 11336 25596 11348
rect 25372 11308 25596 11336
rect 25372 11296 25378 11308
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 26510 11268 26516 11280
rect 25148 11240 26516 11268
rect 26510 11228 26516 11240
rect 26568 11228 26574 11280
rect 25777 11203 25835 11209
rect 25777 11200 25789 11203
rect 24504 11172 25789 11200
rect 24397 11163 24455 11169
rect 25777 11169 25789 11172
rect 25823 11169 25835 11203
rect 25777 11163 25835 11169
rect 23106 11132 23112 11144
rect 21508 11104 21680 11132
rect 22020 11104 22692 11132
rect 23067 11104 23112 11132
rect 21508 11092 21514 11104
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 8849 11067 8907 11073
rect 8849 11064 8861 11067
rect 8812 11036 8861 11064
rect 8812 11024 8818 11036
rect 8849 11033 8861 11036
rect 8895 11033 8907 11067
rect 11425 11067 11483 11073
rect 11425 11064 11437 11067
rect 8849 11027 8907 11033
rect 10980 11036 11437 11064
rect 8352 10968 8432 10996
rect 8352 10956 8358 10968
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 9861 10999 9919 11005
rect 9861 10996 9873 10999
rect 9364 10968 9873 10996
rect 9364 10956 9370 10968
rect 9861 10965 9873 10968
rect 9907 10996 9919 10999
rect 10980 10996 11008 11036
rect 11425 11033 11437 11036
rect 11471 11033 11483 11067
rect 11425 11027 11483 11033
rect 14918 11024 14924 11076
rect 14976 11024 14982 11076
rect 17218 11024 17224 11076
rect 17276 11064 17282 11076
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 17276 11036 17601 11064
rect 17276 11024 17282 11036
rect 17589 11033 17601 11036
rect 17635 11033 17647 11067
rect 17589 11027 17647 11033
rect 19150 11024 19156 11076
rect 19208 11064 19214 11076
rect 19245 11067 19303 11073
rect 19245 11064 19257 11067
rect 19208 11036 19257 11064
rect 19208 11024 19214 11036
rect 19245 11033 19257 11036
rect 19291 11033 19303 11067
rect 19245 11027 19303 11033
rect 20993 11067 21051 11073
rect 20993 11033 21005 11067
rect 21039 11064 21051 11067
rect 22020 11064 22048 11104
rect 22554 11064 22560 11076
rect 21039 11036 22048 11064
rect 22515 11036 22560 11064
rect 21039 11033 21051 11036
rect 20993 11027 21051 11033
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 22664 11064 22692 11104
rect 23106 11092 23112 11104
rect 23164 11092 23170 11144
rect 25038 11132 25044 11144
rect 24999 11104 25044 11132
rect 25038 11092 25044 11104
rect 25096 11132 25102 11144
rect 25222 11132 25228 11144
rect 25096 11104 25228 11132
rect 25096 11092 25102 11104
rect 25222 11092 25228 11104
rect 25280 11092 25286 11144
rect 24118 11064 24124 11076
rect 22664 11036 23778 11064
rect 24079 11036 24124 11064
rect 12066 10996 12072 11008
rect 9907 10968 11008 10996
rect 12027 10968 12072 10996
rect 9907 10965 9919 10968
rect 9861 10959 9919 10965
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 13262 10956 13268 11008
rect 13320 10996 13326 11008
rect 13909 10999 13967 11005
rect 13909 10996 13921 10999
rect 13320 10968 13921 10996
rect 13320 10956 13326 10968
rect 13909 10965 13921 10968
rect 13955 10965 13967 10999
rect 13909 10959 13967 10965
rect 14550 10956 14556 11008
rect 14608 10996 14614 11008
rect 14645 10999 14703 11005
rect 14645 10996 14657 10999
rect 14608 10968 14657 10996
rect 14608 10956 14614 10968
rect 14645 10965 14657 10968
rect 14691 10965 14703 10999
rect 14936 10996 14964 11024
rect 15562 10996 15568 11008
rect 14936 10968 15568 10996
rect 14645 10959 14703 10965
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 22462 10956 22468 11008
rect 22520 10996 22526 11008
rect 22664 10996 22692 11036
rect 23658 10996 23664 11008
rect 22520 10968 22692 10996
rect 23619 10968 23664 10996
rect 22520 10956 22526 10968
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 23750 10996 23778 11036
rect 24118 11024 24124 11036
rect 24176 11024 24182 11076
rect 25409 10999 25467 11005
rect 25409 10996 25421 10999
rect 23750 10968 25421 10996
rect 25409 10965 25421 10968
rect 25455 10965 25467 10999
rect 25409 10959 25467 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1857 10795 1915 10801
rect 1857 10761 1869 10795
rect 1903 10792 1915 10795
rect 2682 10792 2688 10804
rect 1903 10764 2688 10792
rect 1903 10761 1915 10764
rect 1857 10755 1915 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 3234 10792 3240 10804
rect 3195 10764 3240 10792
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5592 10764 5641 10792
rect 5592 10752 5598 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9214 10792 9220 10804
rect 9171 10764 9220 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 9916 10764 10057 10792
rect 9916 10752 9922 10764
rect 10045 10761 10057 10764
rect 10091 10761 10103 10795
rect 10045 10755 10103 10761
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2409 10659 2467 10665
rect 2409 10656 2421 10659
rect 2372 10628 2421 10656
rect 2372 10616 2378 10628
rect 2409 10625 2421 10628
rect 2455 10625 2467 10659
rect 3252 10656 3280 10752
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 3252 10628 3341 10656
rect 2409 10619 2467 10625
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 10060 10656 10088 10755
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11422 10792 11428 10804
rect 11020 10764 11428 10792
rect 11020 10752 11026 10764
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 11606 10792 11612 10804
rect 11567 10764 11612 10792
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12986 10792 12992 10804
rect 12299 10764 12992 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 14642 10792 14648 10804
rect 14599 10764 14648 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 15838 10792 15844 10804
rect 15799 10764 15844 10792
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 16390 10752 16396 10804
rect 16448 10792 16454 10804
rect 16485 10795 16543 10801
rect 16485 10792 16497 10795
rect 16448 10764 16497 10792
rect 16448 10752 16454 10764
rect 16485 10761 16497 10764
rect 16531 10761 16543 10795
rect 16485 10755 16543 10761
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 17405 10795 17463 10801
rect 17405 10792 17417 10795
rect 16632 10764 17417 10792
rect 16632 10752 16638 10764
rect 17405 10761 17417 10764
rect 17451 10761 17463 10795
rect 17405 10755 17463 10761
rect 18417 10795 18475 10801
rect 18417 10761 18429 10795
rect 18463 10792 18475 10795
rect 18506 10792 18512 10804
rect 18463 10764 18512 10792
rect 18463 10761 18475 10764
rect 18417 10755 18475 10761
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 18601 10795 18659 10801
rect 18601 10761 18613 10795
rect 18647 10792 18659 10795
rect 19058 10792 19064 10804
rect 18647 10764 19064 10792
rect 18647 10761 18659 10764
rect 18601 10755 18659 10761
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 21450 10792 21456 10804
rect 21411 10764 21456 10792
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 21729 10795 21787 10801
rect 21729 10761 21741 10795
rect 21775 10792 21787 10795
rect 22002 10792 22008 10804
rect 21775 10764 22008 10792
rect 21775 10761 21787 10764
rect 21729 10755 21787 10761
rect 10318 10724 10324 10736
rect 10279 10696 10324 10724
rect 10318 10684 10324 10696
rect 10376 10684 10382 10736
rect 11330 10724 11336 10736
rect 11243 10696 11336 10724
rect 11330 10684 11336 10696
rect 11388 10724 11394 10736
rect 12342 10724 12348 10736
rect 11388 10696 12348 10724
rect 11388 10684 11394 10696
rect 12342 10684 12348 10696
rect 12400 10724 12406 10736
rect 12713 10727 12771 10733
rect 12713 10724 12725 10727
rect 12400 10696 12725 10724
rect 12400 10684 12406 10696
rect 12713 10693 12725 10696
rect 12759 10724 12771 10727
rect 13170 10724 13176 10736
rect 12759 10696 13176 10724
rect 12759 10693 12771 10696
rect 12713 10687 12771 10693
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 14737 10727 14795 10733
rect 14737 10724 14749 10727
rect 13872 10696 14749 10724
rect 13872 10684 13878 10696
rect 14737 10693 14749 10696
rect 14783 10693 14795 10727
rect 14737 10687 14795 10693
rect 19334 10684 19340 10736
rect 19392 10724 19398 10736
rect 19521 10727 19579 10733
rect 19521 10724 19533 10727
rect 19392 10696 19533 10724
rect 19392 10684 19398 10696
rect 19521 10693 19533 10696
rect 19567 10724 19579 10727
rect 19610 10724 19616 10736
rect 19567 10696 19616 10724
rect 19567 10693 19579 10696
rect 19521 10687 19579 10693
rect 19610 10684 19616 10696
rect 19668 10684 19674 10736
rect 20162 10724 20168 10736
rect 20123 10696 20168 10724
rect 20162 10684 20168 10696
rect 20220 10684 20226 10736
rect 21177 10727 21235 10733
rect 21177 10693 21189 10727
rect 21223 10724 21235 10727
rect 21634 10724 21640 10736
rect 21223 10696 21640 10724
rect 21223 10693 21235 10696
rect 21177 10687 21235 10693
rect 21634 10684 21640 10696
rect 21692 10684 21698 10736
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 7616 10628 7880 10656
rect 10060 10628 10701 10656
rect 7616 10616 7622 10628
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 5626 10588 5632 10600
rect 1719 10560 5632 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 1946 10480 1952 10532
rect 2004 10520 2010 10532
rect 2133 10523 2191 10529
rect 2133 10520 2145 10523
rect 2004 10492 2145 10520
rect 2004 10480 2010 10492
rect 2133 10489 2145 10492
rect 2179 10520 2191 10523
rect 2222 10520 2228 10532
rect 2179 10492 2228 10520
rect 2179 10489 2191 10492
rect 2133 10483 2191 10489
rect 2222 10480 2228 10492
rect 2280 10480 2286 10532
rect 2332 10529 2360 10560
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7576 10560 7757 10588
rect 2317 10523 2375 10529
rect 2317 10489 2329 10523
rect 2363 10489 2375 10523
rect 2317 10483 2375 10489
rect 2869 10523 2927 10529
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 3574 10523 3632 10529
rect 3574 10520 3586 10523
rect 2915 10492 3586 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 3574 10489 3586 10492
rect 3620 10520 3632 10523
rect 4614 10520 4620 10532
rect 3620 10492 4620 10520
rect 3620 10489 3632 10492
rect 3574 10483 3632 10489
rect 4614 10480 4620 10492
rect 4672 10520 4678 10532
rect 6549 10523 6607 10529
rect 6549 10520 6561 10523
rect 4672 10492 6561 10520
rect 4672 10480 4678 10492
rect 6549 10489 6561 10492
rect 6595 10520 6607 10523
rect 7190 10520 7196 10532
rect 6595 10492 7196 10520
rect 6595 10489 6607 10492
rect 6549 10483 6607 10489
rect 7190 10480 7196 10492
rect 7248 10480 7254 10532
rect 7576 10464 7604 10560
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 7852 10588 7880 10628
rect 10689 10625 10701 10628
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13725 10659 13783 10665
rect 13725 10656 13737 10659
rect 13044 10628 13737 10656
rect 13044 10616 13050 10628
rect 13725 10625 13737 10628
rect 13771 10625 13783 10659
rect 13725 10619 13783 10625
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 15378 10656 15384 10668
rect 14231 10628 15384 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 8001 10591 8059 10597
rect 8001 10588 8013 10591
rect 7852 10560 8013 10588
rect 7745 10551 7803 10557
rect 8001 10557 8013 10560
rect 8047 10557 8059 10591
rect 8001 10551 8059 10557
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 13446 10588 13452 10600
rect 12492 10560 13452 10588
rect 12492 10548 12498 10560
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 14200 10588 14228 10619
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 16850 10616 16856 10668
rect 16908 10656 16914 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16908 10628 17049 10656
rect 16908 10616 16914 10628
rect 17037 10625 17049 10628
rect 17083 10656 17095 10659
rect 17862 10656 17868 10668
rect 17083 10628 17868 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 19061 10659 19119 10665
rect 19061 10625 19073 10659
rect 19107 10656 19119 10659
rect 21744 10656 21772 10755
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 22741 10795 22799 10801
rect 22741 10761 22753 10795
rect 22787 10792 22799 10795
rect 23014 10792 23020 10804
rect 22787 10764 23020 10792
rect 22787 10761 22799 10764
rect 22741 10755 22799 10761
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 23474 10792 23480 10804
rect 23435 10764 23480 10792
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 24118 10752 24124 10804
rect 24176 10792 24182 10804
rect 24673 10795 24731 10801
rect 24673 10792 24685 10795
rect 24176 10764 24685 10792
rect 24176 10752 24182 10764
rect 24673 10761 24685 10764
rect 24719 10761 24731 10795
rect 24673 10755 24731 10761
rect 23753 10727 23811 10733
rect 23753 10693 23765 10727
rect 23799 10724 23811 10727
rect 24762 10724 24768 10736
rect 23799 10696 24768 10724
rect 23799 10693 23811 10696
rect 23753 10687 23811 10693
rect 24762 10684 24768 10696
rect 24820 10684 24826 10736
rect 19107 10628 21772 10656
rect 22189 10659 22247 10665
rect 19107 10625 19119 10628
rect 19061 10619 19119 10625
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22738 10656 22744 10668
rect 22235 10628 22744 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 13648 10560 14228 10588
rect 10873 10523 10931 10529
rect 10873 10489 10885 10523
rect 10919 10520 10931 10523
rect 10962 10520 10968 10532
rect 10919 10492 10968 10520
rect 10919 10489 10931 10492
rect 10873 10483 10931 10489
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 12066 10480 12072 10532
rect 12124 10520 12130 10532
rect 13170 10529 13176 10532
rect 13155 10523 13176 10529
rect 13155 10520 13167 10523
rect 12124 10492 13167 10520
rect 12124 10480 12130 10492
rect 13155 10489 13167 10492
rect 13228 10520 13234 10532
rect 13648 10529 13676 10560
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 14608 10560 15301 10588
rect 14608 10548 14614 10560
rect 15289 10557 15301 10560
rect 15335 10588 15347 10591
rect 16666 10588 16672 10600
rect 15335 10560 16672 10588
rect 15335 10557 15347 10560
rect 15289 10551 15347 10557
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 19978 10548 19984 10600
rect 20036 10588 20042 10600
rect 22204 10588 22232 10619
rect 22738 10616 22744 10628
rect 22796 10616 22802 10668
rect 22830 10616 22836 10668
rect 22888 10656 22894 10668
rect 23017 10659 23075 10665
rect 23017 10656 23029 10659
rect 22888 10628 23029 10656
rect 22888 10616 22894 10628
rect 23017 10625 23029 10628
rect 23063 10625 23075 10659
rect 23198 10656 23204 10668
rect 23017 10619 23075 10625
rect 23124 10628 23204 10656
rect 20036 10560 22232 10588
rect 20036 10548 20042 10560
rect 13633 10523 13691 10529
rect 13228 10492 13303 10520
rect 13155 10483 13176 10489
rect 13170 10480 13176 10483
rect 13228 10480 13234 10492
rect 13633 10489 13645 10523
rect 13679 10489 13691 10523
rect 13633 10483 13691 10489
rect 14826 10480 14832 10532
rect 14884 10520 14890 10532
rect 15013 10523 15071 10529
rect 15013 10520 15025 10523
rect 14884 10492 15025 10520
rect 14884 10480 14890 10492
rect 15013 10489 15025 10492
rect 15059 10489 15071 10523
rect 15013 10483 15071 10489
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 16209 10523 16267 10529
rect 16209 10520 16221 10523
rect 15620 10492 16221 10520
rect 15620 10480 15626 10492
rect 16209 10489 16221 10492
rect 16255 10489 16267 10523
rect 16209 10483 16267 10489
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10452 4767 10455
rect 4798 10452 4804 10464
rect 4755 10424 4804 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 4798 10412 4804 10424
rect 4856 10452 4862 10464
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 4856 10424 5273 10452
rect 4856 10412 4862 10424
rect 5261 10421 5273 10424
rect 5307 10421 5319 10455
rect 5261 10415 5319 10421
rect 5902 10412 5908 10464
rect 5960 10452 5966 10464
rect 5997 10455 6055 10461
rect 5997 10452 6009 10455
rect 5960 10424 6009 10452
rect 5960 10412 5966 10424
rect 5997 10421 6009 10424
rect 6043 10421 6055 10455
rect 7006 10452 7012 10464
rect 6967 10424 7012 10452
rect 5997 10415 6055 10421
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7558 10452 7564 10464
rect 7519 10424 7564 10452
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 9769 10455 9827 10461
rect 9769 10421 9781 10455
rect 9815 10452 9827 10455
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 9815 10424 10793 10452
rect 9815 10421 9827 10424
rect 9769 10415 9827 10421
rect 10781 10421 10793 10424
rect 10827 10452 10839 10455
rect 11330 10452 11336 10464
rect 10827 10424 11336 10452
rect 10827 10421 10839 10424
rect 10781 10415 10839 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 14642 10412 14648 10464
rect 14700 10452 14706 10464
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 14700 10424 15209 10452
rect 14700 10412 14706 10424
rect 15197 10421 15209 10424
rect 15243 10421 15255 10455
rect 16224 10452 16252 10483
rect 16390 10480 16396 10532
rect 16448 10520 16454 10532
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 16448 10492 16773 10520
rect 16448 10480 16454 10492
rect 16761 10489 16773 10492
rect 16807 10489 16819 10523
rect 16761 10483 16819 10489
rect 17865 10523 17923 10529
rect 17865 10489 17877 10523
rect 17911 10520 17923 10523
rect 18966 10520 18972 10532
rect 17911 10492 18972 10520
rect 17911 10489 17923 10492
rect 17865 10483 17923 10489
rect 18966 10480 18972 10492
rect 19024 10520 19030 10532
rect 19153 10523 19211 10529
rect 19153 10520 19165 10523
rect 19024 10492 19165 10520
rect 19024 10480 19030 10492
rect 19153 10489 19165 10492
rect 19199 10489 19211 10523
rect 19153 10483 19211 10489
rect 20070 10480 20076 10532
rect 20128 10520 20134 10532
rect 20441 10523 20499 10529
rect 20441 10520 20453 10523
rect 20128 10492 20453 10520
rect 20128 10480 20134 10492
rect 20441 10489 20453 10492
rect 20487 10489 20499 10523
rect 20441 10483 20499 10489
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 22002 10520 22008 10532
rect 20772 10492 22008 10520
rect 20772 10480 20778 10492
rect 22002 10480 22008 10492
rect 22060 10520 22066 10532
rect 22281 10523 22339 10529
rect 22281 10520 22293 10523
rect 22060 10492 22293 10520
rect 22060 10480 22066 10492
rect 22281 10489 22293 10492
rect 22327 10489 22339 10523
rect 22281 10483 22339 10489
rect 22462 10480 22468 10532
rect 22520 10480 22526 10532
rect 22830 10480 22836 10532
rect 22888 10520 22894 10532
rect 23124 10520 23152 10628
rect 23198 10616 23204 10628
rect 23256 10616 23262 10668
rect 23934 10616 23940 10668
rect 23992 10656 23998 10668
rect 23992 10628 24440 10656
rect 23992 10616 23998 10628
rect 23658 10548 23664 10600
rect 23716 10588 23722 10600
rect 24210 10588 24216 10600
rect 23716 10560 24216 10588
rect 23716 10548 23722 10560
rect 24210 10548 24216 10560
rect 24268 10588 24274 10600
rect 24305 10591 24363 10597
rect 24305 10588 24317 10591
rect 24268 10560 24317 10588
rect 24268 10548 24274 10560
rect 24305 10557 24317 10560
rect 24351 10557 24363 10591
rect 24305 10551 24363 10557
rect 22888 10492 23152 10520
rect 22888 10480 22894 10492
rect 23198 10480 23204 10532
rect 23256 10520 23262 10532
rect 23256 10492 23520 10520
rect 23256 10480 23262 10492
rect 16945 10455 17003 10461
rect 16945 10452 16957 10455
rect 16224 10424 16957 10452
rect 15197 10415 15255 10421
rect 16945 10421 16957 10424
rect 16991 10421 17003 10455
rect 16945 10415 17003 10421
rect 19061 10455 19119 10461
rect 19061 10421 19073 10455
rect 19107 10452 19119 10455
rect 19242 10452 19248 10464
rect 19107 10424 19248 10452
rect 19107 10421 19119 10424
rect 19061 10415 19119 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 19981 10455 20039 10461
rect 19981 10421 19993 10455
rect 20027 10452 20039 10455
rect 20625 10455 20683 10461
rect 20625 10452 20637 10455
rect 20027 10424 20637 10452
rect 20027 10421 20039 10424
rect 19981 10415 20039 10421
rect 20625 10421 20637 10424
rect 20671 10452 20683 10455
rect 22094 10452 22100 10464
rect 20671 10424 22100 10452
rect 20671 10421 20683 10424
rect 20625 10415 20683 10421
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 22189 10455 22247 10461
rect 22189 10421 22201 10455
rect 22235 10452 22247 10455
rect 22480 10452 22508 10480
rect 22235 10424 22508 10452
rect 23492 10452 23520 10492
rect 23934 10480 23940 10532
rect 23992 10520 23998 10532
rect 24029 10523 24087 10529
rect 24029 10520 24041 10523
rect 23992 10492 24041 10520
rect 23992 10480 23998 10492
rect 24029 10489 24041 10492
rect 24075 10489 24087 10523
rect 24412 10520 24440 10628
rect 24670 10616 24676 10668
rect 24728 10656 24734 10668
rect 25041 10659 25099 10665
rect 25041 10656 25053 10659
rect 24728 10628 25053 10656
rect 24728 10616 24734 10628
rect 25041 10625 25053 10628
rect 25087 10625 25099 10659
rect 25041 10619 25099 10625
rect 25501 10659 25559 10665
rect 25501 10625 25513 10659
rect 25547 10656 25559 10659
rect 25774 10656 25780 10668
rect 25547 10628 25780 10656
rect 25547 10625 25559 10628
rect 25501 10619 25559 10625
rect 25774 10616 25780 10628
rect 25832 10616 25838 10668
rect 25222 10588 25228 10600
rect 25183 10560 25228 10588
rect 25222 10548 25228 10560
rect 25280 10588 25286 10600
rect 25961 10591 26019 10597
rect 25961 10588 25973 10591
rect 25280 10560 25973 10588
rect 25280 10548 25286 10560
rect 25961 10557 25973 10560
rect 26007 10557 26019 10591
rect 25961 10551 26019 10557
rect 26234 10520 26240 10532
rect 24412 10492 26240 10520
rect 24029 10483 24087 10489
rect 26234 10480 26240 10492
rect 26292 10480 26298 10532
rect 24213 10455 24271 10461
rect 24213 10452 24225 10455
rect 23492 10424 24225 10452
rect 22235 10421 22247 10424
rect 22189 10415 22247 10421
rect 24213 10421 24225 10424
rect 24259 10421 24271 10455
rect 24213 10415 24271 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 2314 10208 2320 10220
rect 2372 10248 2378 10260
rect 2498 10248 2504 10260
rect 2372 10220 2504 10248
rect 2372 10208 2378 10220
rect 2498 10208 2504 10220
rect 2556 10248 2562 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 2556 10220 3617 10248
rect 2556 10208 2562 10220
rect 2958 10180 2964 10192
rect 2919 10152 2964 10180
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 3068 10189 3096 10220
rect 3605 10217 3617 10220
rect 3651 10248 3663 10251
rect 4062 10248 4068 10260
rect 3651 10220 4068 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4338 10248 4344 10260
rect 4299 10220 4344 10248
rect 4338 10208 4344 10220
rect 4396 10208 4402 10260
rect 5258 10248 5264 10260
rect 5219 10220 5264 10248
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 5684 10220 7052 10248
rect 5684 10208 5690 10220
rect 3053 10183 3111 10189
rect 3053 10149 3065 10183
rect 3099 10180 3111 10183
rect 5077 10183 5135 10189
rect 3099 10152 3133 10180
rect 3099 10149 3111 10152
rect 3053 10143 3111 10149
rect 5077 10149 5089 10183
rect 5123 10180 5135 10183
rect 5166 10180 5172 10192
rect 5123 10152 5172 10180
rect 5123 10149 5135 10152
rect 5077 10143 5135 10149
rect 5166 10140 5172 10152
rect 5224 10140 5230 10192
rect 6181 10183 6239 10189
rect 6181 10149 6193 10183
rect 6227 10180 6239 10183
rect 6518 10183 6576 10189
rect 6518 10180 6530 10183
rect 6227 10152 6530 10180
rect 6227 10149 6239 10152
rect 6181 10143 6239 10149
rect 6518 10149 6530 10152
rect 6564 10180 6576 10183
rect 6914 10180 6920 10192
rect 6564 10152 6920 10180
rect 6564 10149 6576 10152
rect 6518 10143 6576 10149
rect 6914 10140 6920 10152
rect 6972 10140 6978 10192
rect 7024 10180 7052 10220
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7248 10220 7665 10248
rect 7248 10208 7254 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 7653 10211 7711 10217
rect 8849 10251 8907 10257
rect 8849 10217 8861 10251
rect 8895 10248 8907 10251
rect 9306 10248 9312 10260
rect 8895 10220 9312 10248
rect 8895 10217 8907 10220
rect 8849 10211 8907 10217
rect 9306 10208 9312 10220
rect 9364 10248 9370 10260
rect 10962 10248 10968 10260
rect 9364 10220 10968 10248
rect 9364 10208 9370 10220
rect 7024 10152 7696 10180
rect 4614 10072 4620 10124
rect 4672 10112 4678 10124
rect 5353 10115 5411 10121
rect 5353 10112 5365 10115
rect 4672 10084 5365 10112
rect 4672 10072 4678 10084
rect 5353 10081 5365 10084
rect 5399 10081 5411 10115
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 5353 10075 5411 10081
rect 5460 10084 6285 10112
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2682 10004 2688 10056
rect 2740 10044 2746 10056
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 2740 10016 2973 10044
rect 2740 10004 2746 10016
rect 2961 10013 2973 10016
rect 3007 10044 3019 10047
rect 3007 10016 4292 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 2501 9979 2559 9985
rect 2501 9945 2513 9979
rect 2547 9976 2559 9979
rect 3418 9976 3424 9988
rect 2547 9948 3424 9976
rect 2547 9945 2559 9948
rect 2501 9939 2559 9945
rect 3418 9936 3424 9948
rect 3476 9936 3482 9988
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 4154 9908 4160 9920
rect 3108 9880 4160 9908
rect 3108 9868 3114 9880
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4264 9908 4292 10016
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 5166 10044 5172 10056
rect 4396 10016 5172 10044
rect 4396 10004 4402 10016
rect 5166 10004 5172 10016
rect 5224 10044 5230 10056
rect 5460 10044 5488 10084
rect 6273 10081 6285 10084
rect 6319 10112 6331 10115
rect 7558 10112 7564 10124
rect 6319 10084 7564 10112
rect 6319 10081 6331 10084
rect 6273 10075 6331 10081
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 5718 10044 5724 10056
rect 5224 10016 5488 10044
rect 5679 10016 5724 10044
rect 5224 10004 5230 10016
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 5902 10004 5908 10056
rect 5960 10044 5966 10056
rect 6086 10044 6092 10056
rect 5960 10016 6092 10044
rect 5960 10004 5966 10016
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 7668 10044 7696 10152
rect 10134 10140 10140 10192
rect 10192 10180 10198 10192
rect 10336 10189 10364 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 12621 10251 12679 10257
rect 12621 10217 12633 10251
rect 12667 10248 12679 10251
rect 13170 10248 13176 10260
rect 12667 10220 13176 10248
rect 12667 10217 12679 10220
rect 12621 10211 12679 10217
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 16390 10248 16396 10260
rect 16351 10220 16396 10248
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 16850 10248 16856 10260
rect 16811 10220 16856 10248
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 18322 10248 18328 10260
rect 18283 10220 18328 10248
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 19518 10248 19524 10260
rect 19479 10220 19524 10248
rect 19518 10208 19524 10220
rect 19576 10248 19582 10260
rect 20625 10251 20683 10257
rect 20625 10248 20637 10251
rect 19576 10220 20637 10248
rect 19576 10208 19582 10220
rect 20625 10217 20637 10220
rect 20671 10217 20683 10251
rect 20625 10211 20683 10217
rect 10229 10183 10287 10189
rect 10229 10180 10241 10183
rect 10192 10152 10241 10180
rect 10192 10140 10198 10152
rect 10229 10149 10241 10152
rect 10275 10149 10287 10183
rect 10229 10143 10287 10149
rect 10321 10183 10379 10189
rect 10321 10149 10333 10183
rect 10367 10149 10379 10183
rect 10321 10143 10379 10149
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8352 10084 9137 10112
rect 8352 10072 8358 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 10244 10112 10272 10143
rect 12342 10140 12348 10192
rect 12400 10180 12406 10192
rect 12713 10183 12771 10189
rect 12713 10180 12725 10183
rect 12400 10152 12725 10180
rect 12400 10140 12406 10152
rect 12713 10149 12725 10152
rect 12759 10180 12771 10183
rect 13262 10180 13268 10192
rect 12759 10152 13268 10180
rect 12759 10149 12771 10152
rect 12713 10143 12771 10149
rect 13262 10140 13268 10152
rect 13320 10140 13326 10192
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 14185 10183 14243 10189
rect 14185 10180 14197 10183
rect 13872 10152 14197 10180
rect 13872 10140 13878 10152
rect 14185 10149 14197 10152
rect 14231 10180 14243 10183
rect 15562 10180 15568 10192
rect 14231 10152 15568 10180
rect 14231 10149 14243 10152
rect 14185 10143 14243 10149
rect 15562 10140 15568 10152
rect 15620 10140 15626 10192
rect 15746 10140 15752 10192
rect 15804 10180 15810 10192
rect 15933 10183 15991 10189
rect 15933 10180 15945 10183
rect 15804 10152 15945 10180
rect 15804 10140 15810 10152
rect 15933 10149 15945 10152
rect 15979 10149 15991 10183
rect 17494 10180 17500 10192
rect 17455 10152 17500 10180
rect 15933 10143 15991 10149
rect 17494 10140 17500 10152
rect 17552 10140 17558 10192
rect 17954 10180 17960 10192
rect 17915 10152 17960 10180
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 19058 10180 19064 10192
rect 19019 10152 19064 10180
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 20070 10180 20076 10192
rect 20031 10152 20076 10180
rect 20070 10140 20076 10152
rect 20128 10140 20134 10192
rect 20640 10180 20668 10211
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 22060 10220 22293 10248
rect 22060 10208 22066 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22281 10211 22339 10217
rect 22649 10251 22707 10257
rect 22649 10217 22661 10251
rect 22695 10248 22707 10251
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 22695 10220 22937 10248
rect 22695 10217 22707 10220
rect 22649 10211 22707 10217
rect 22925 10217 22937 10220
rect 22971 10248 22983 10251
rect 23106 10248 23112 10260
rect 22971 10220 23112 10248
rect 22971 10217 22983 10220
rect 22925 10211 22983 10217
rect 23106 10208 23112 10220
rect 23164 10208 23170 10260
rect 23934 10208 23940 10260
rect 23992 10248 23998 10260
rect 25317 10251 25375 10257
rect 25317 10248 25329 10251
rect 23992 10220 25329 10248
rect 23992 10208 23998 10220
rect 25317 10217 25329 10220
rect 25363 10217 25375 10251
rect 25317 10211 25375 10217
rect 25406 10208 25412 10260
rect 25464 10248 25470 10260
rect 25685 10251 25743 10257
rect 25685 10248 25697 10251
rect 25464 10220 25697 10248
rect 25464 10208 25470 10220
rect 25685 10217 25697 10220
rect 25731 10217 25743 10251
rect 25685 10211 25743 10217
rect 20714 10180 20720 10192
rect 20627 10152 20720 10180
rect 20714 10140 20720 10152
rect 20772 10180 20778 10192
rect 21146 10183 21204 10189
rect 21146 10180 21158 10183
rect 20772 10152 21158 10180
rect 20772 10140 20778 10152
rect 21146 10149 21158 10152
rect 21192 10149 21204 10183
rect 21146 10143 21204 10149
rect 21358 10140 21364 10192
rect 21416 10180 21422 10192
rect 22462 10180 22468 10192
rect 21416 10152 22468 10180
rect 21416 10140 21422 10152
rect 22462 10140 22468 10152
rect 22520 10140 22526 10192
rect 10502 10112 10508 10124
rect 10244 10084 10508 10112
rect 9125 10075 9183 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10612 10084 12572 10112
rect 10226 10044 10232 10056
rect 7668 10016 10088 10044
rect 10187 10016 10232 10044
rect 4801 9979 4859 9985
rect 4801 9945 4813 9979
rect 4847 9976 4859 9979
rect 4890 9976 4896 9988
rect 4847 9948 4896 9976
rect 4847 9945 4859 9948
rect 4801 9939 4859 9945
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 9272 9948 9628 9976
rect 9272 9936 9278 9948
rect 7190 9908 7196 9920
rect 4264 9880 7196 9908
rect 7190 9868 7196 9880
rect 7248 9908 7254 9920
rect 7742 9908 7748 9920
rect 7248 9880 7748 9908
rect 7248 9868 7254 9880
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 8481 9911 8539 9917
rect 8481 9877 8493 9911
rect 8527 9908 8539 9911
rect 9398 9908 9404 9920
rect 8527 9880 9404 9908
rect 8527 9877 8539 9880
rect 8481 9871 8539 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 9600 9908 9628 9948
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 9769 9979 9827 9985
rect 9769 9976 9781 9979
rect 9732 9948 9781 9976
rect 9732 9936 9738 9948
rect 9769 9945 9781 9948
rect 9815 9945 9827 9979
rect 10060 9976 10088 10016
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10410 10004 10416 10056
rect 10468 10044 10474 10056
rect 10612 10044 10640 10084
rect 10468 10016 10640 10044
rect 10468 10004 10474 10016
rect 10686 10004 10692 10056
rect 10744 10044 10750 10056
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 10744 10016 11529 10044
rect 10744 10004 10750 10016
rect 11517 10013 11529 10016
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 11054 9976 11060 9988
rect 10060 9948 11060 9976
rect 9769 9939 9827 9945
rect 11054 9936 11060 9948
rect 11112 9936 11118 9988
rect 11146 9936 11152 9988
rect 11204 9976 11210 9988
rect 12161 9979 12219 9985
rect 12161 9976 12173 9979
rect 11204 9948 12173 9976
rect 11204 9936 11210 9948
rect 12161 9945 12173 9948
rect 12207 9945 12219 9979
rect 12161 9939 12219 9945
rect 10410 9908 10416 9920
rect 9600 9880 10416 9908
rect 10410 9868 10416 9880
rect 10468 9868 10474 9920
rect 10594 9868 10600 9920
rect 10652 9908 10658 9920
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 10652 9880 10793 9908
rect 10652 9868 10658 9880
rect 10781 9877 10793 9880
rect 10827 9877 10839 9911
rect 10781 9871 10839 9877
rect 11241 9911 11299 9917
rect 11241 9877 11253 9911
rect 11287 9908 11299 9911
rect 11422 9908 11428 9920
rect 11287 9880 11428 9908
rect 11287 9877 11299 9880
rect 11241 9871 11299 9877
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 11882 9908 11888 9920
rect 11843 9880 11888 9908
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12544 9908 12572 10084
rect 12986 10072 12992 10124
rect 13044 10112 13050 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 13044 10084 13185 10112
rect 13044 10072 13050 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 13541 10115 13599 10121
rect 13541 10081 13553 10115
rect 13587 10112 13599 10115
rect 13587 10084 14320 10112
rect 13587 10081 13599 10084
rect 13541 10075 13599 10081
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 13078 10044 13084 10056
rect 12667 10016 13084 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 14182 10044 14188 10056
rect 14143 10016 14188 10044
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14292 10053 14320 10084
rect 15378 10072 15384 10124
rect 15436 10112 15442 10124
rect 16025 10115 16083 10121
rect 16025 10112 16037 10115
rect 15436 10084 16037 10112
rect 15436 10072 15442 10084
rect 16025 10081 16037 10084
rect 16071 10112 16083 10115
rect 16482 10112 16488 10124
rect 16071 10084 16488 10112
rect 16071 10081 16083 10084
rect 16025 10075 16083 10081
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 23652 10115 23710 10121
rect 23652 10081 23664 10115
rect 23698 10112 23710 10115
rect 23934 10112 23940 10124
rect 23698 10084 23940 10112
rect 23698 10081 23710 10084
rect 23652 10075 23710 10081
rect 23934 10072 23940 10084
rect 23992 10072 23998 10124
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 14550 10044 14556 10056
rect 14323 10016 14556 10044
rect 14323 10013 14335 10016
rect 14277 10007 14335 10013
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10013 15991 10047
rect 17402 10044 17408 10056
rect 17363 10016 17408 10044
rect 15933 10007 15991 10013
rect 13722 9976 13728 9988
rect 13683 9948 13728 9976
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 14090 9936 14096 9988
rect 14148 9976 14154 9988
rect 15013 9979 15071 9985
rect 15013 9976 15025 9979
rect 14148 9948 15025 9976
rect 14148 9936 14154 9948
rect 15013 9945 15025 9948
rect 15059 9976 15071 9979
rect 15470 9976 15476 9988
rect 15059 9948 15148 9976
rect 15431 9948 15476 9976
rect 15059 9945 15071 9948
rect 15013 9939 15071 9945
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 12544 9880 14657 9908
rect 14645 9877 14657 9880
rect 14691 9908 14703 9911
rect 14826 9908 14832 9920
rect 14691 9880 14832 9908
rect 14691 9877 14703 9880
rect 14645 9871 14703 9877
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 15120 9908 15148 9948
rect 15470 9936 15476 9948
rect 15528 9936 15534 9988
rect 15948 9976 15976 10007
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 17586 10044 17592 10056
rect 17547 10016 17592 10044
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 19061 10047 19119 10053
rect 19061 10013 19073 10047
rect 19107 10013 19119 10047
rect 19061 10007 19119 10013
rect 18598 9976 18604 9988
rect 15948 9948 17080 9976
rect 18559 9948 18604 9976
rect 17052 9920 17080 9948
rect 18598 9936 18604 9948
rect 18656 9936 18662 9988
rect 19076 9976 19104 10007
rect 19150 10004 19156 10056
rect 19208 10044 19214 10056
rect 20898 10044 20904 10056
rect 19208 10016 19253 10044
rect 20859 10016 20904 10044
rect 19208 10004 19214 10016
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 22738 10004 22744 10056
rect 22796 10044 22802 10056
rect 23385 10047 23443 10053
rect 23385 10044 23397 10047
rect 22796 10016 23397 10044
rect 22796 10004 22802 10016
rect 23385 10013 23397 10016
rect 23431 10013 23443 10047
rect 23385 10007 23443 10013
rect 19242 9976 19248 9988
rect 19076 9948 19248 9976
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 23014 9936 23020 9988
rect 23072 9976 23078 9988
rect 23072 9948 23428 9976
rect 23072 9936 23078 9948
rect 15562 9908 15568 9920
rect 15120 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 17034 9908 17040 9920
rect 16995 9880 17040 9908
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 22649 9911 22707 9917
rect 22649 9908 22661 9911
rect 22060 9880 22661 9908
rect 22060 9868 22066 9880
rect 22649 9877 22661 9880
rect 22695 9877 22707 9911
rect 23198 9908 23204 9920
rect 23159 9880 23204 9908
rect 22649 9871 22707 9877
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 23400 9908 23428 9948
rect 24670 9936 24676 9988
rect 24728 9976 24734 9988
rect 24765 9979 24823 9985
rect 24765 9976 24777 9979
rect 24728 9948 24777 9976
rect 24728 9936 24734 9948
rect 24765 9945 24777 9948
rect 24811 9945 24823 9979
rect 24765 9939 24823 9945
rect 25406 9936 25412 9988
rect 25464 9976 25470 9988
rect 25958 9976 25964 9988
rect 25464 9948 25964 9976
rect 25464 9936 25470 9948
rect 25958 9936 25964 9948
rect 26016 9936 26022 9988
rect 24946 9908 24952 9920
rect 23400 9880 24952 9908
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 25222 9868 25228 9920
rect 25280 9908 25286 9920
rect 26053 9911 26111 9917
rect 26053 9908 26065 9911
rect 25280 9880 26065 9908
rect 25280 9868 25286 9880
rect 26053 9877 26065 9880
rect 26099 9877 26111 9911
rect 26053 9871 26111 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2682 9664 2688 9716
rect 2740 9664 2746 9716
rect 4614 9704 4620 9716
rect 4575 9676 4620 9704
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 6270 9664 6276 9716
rect 6328 9704 6334 9716
rect 6917 9707 6975 9713
rect 6917 9704 6929 9707
rect 6328 9676 6929 9704
rect 6328 9664 6334 9676
rect 6917 9673 6929 9676
rect 6963 9673 6975 9707
rect 6917 9667 6975 9673
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7837 9707 7895 9713
rect 7837 9704 7849 9707
rect 7616 9676 7849 9704
rect 7616 9664 7622 9676
rect 7837 9673 7849 9676
rect 7883 9673 7895 9707
rect 7837 9667 7895 9673
rect 10594 9664 10600 9716
rect 10652 9704 10658 9716
rect 10652 9676 11008 9704
rect 10652 9664 10658 9676
rect 2130 9636 2136 9648
rect 2091 9608 2136 9636
rect 2130 9596 2136 9608
rect 2188 9596 2194 9648
rect 2700 9636 2728 9664
rect 2424 9608 2728 9636
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2424 9568 2452 9608
rect 3142 9596 3148 9648
rect 3200 9636 3206 9648
rect 3697 9639 3755 9645
rect 3697 9636 3709 9639
rect 3200 9608 3709 9636
rect 3200 9596 3206 9608
rect 3697 9605 3709 9608
rect 3743 9605 3755 9639
rect 3697 9599 3755 9605
rect 4706 9596 4712 9648
rect 4764 9636 4770 9648
rect 4890 9636 4896 9648
rect 4764 9608 4896 9636
rect 4764 9596 4770 9608
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 5258 9636 5264 9648
rect 5219 9608 5264 9636
rect 5258 9596 5264 9608
rect 5316 9596 5322 9648
rect 2590 9568 2596 9580
rect 1995 9540 2452 9568
rect 2503 9540 2596 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2590 9528 2596 9540
rect 2648 9568 2654 9580
rect 3786 9568 3792 9580
rect 2648 9540 3792 9568
rect 2648 9528 2654 9540
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 4212 9540 4261 9568
rect 4212 9528 4218 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 4338 9528 4344 9580
rect 4396 9568 4402 9580
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 4396 9540 5733 9568
rect 4396 9528 4402 9540
rect 5721 9537 5733 9540
rect 5767 9568 5779 9571
rect 6178 9568 6184 9580
rect 5767 9540 6184 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 2498 9460 2504 9512
rect 2556 9500 2562 9512
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2556 9472 2697 9500
rect 2556 9460 2562 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3936 9472 3985 9500
rect 3936 9460 3942 9472
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 5626 9500 5632 9512
rect 5224 9472 5632 9500
rect 5224 9460 5230 9472
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 6288 9500 6316 9664
rect 8481 9639 8539 9645
rect 8481 9605 8493 9639
rect 8527 9636 8539 9639
rect 8938 9636 8944 9648
rect 8527 9608 8944 9636
rect 8527 9605 8539 9608
rect 8481 9599 8539 9605
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 10870 9636 10876 9648
rect 10831 9608 10876 9636
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8570 9568 8576 9580
rect 8343 9540 8576 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8570 9528 8576 9540
rect 8628 9568 8634 9580
rect 9033 9571 9091 9577
rect 8628 9540 8984 9568
rect 8628 9528 8634 9540
rect 5736 9472 6316 9500
rect 6365 9503 6423 9509
rect 5736 9441 5764 9472
rect 6365 9469 6377 9503
rect 6411 9500 6423 9503
rect 7282 9500 7288 9512
rect 6411 9472 7288 9500
rect 6411 9469 6423 9472
rect 6365 9463 6423 9469
rect 7282 9460 7288 9472
rect 7340 9500 7346 9512
rect 7340 9472 7420 9500
rect 7340 9460 7346 9472
rect 5721 9435 5779 9441
rect 5721 9401 5733 9435
rect 5767 9401 5779 9435
rect 5721 9395 5779 9401
rect 5813 9435 5871 9441
rect 5813 9401 5825 9435
rect 5859 9432 5871 9435
rect 7006 9432 7012 9444
rect 5859 9404 7012 9432
rect 5859 9401 5871 9404
rect 5813 9395 5871 9401
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 2593 9367 2651 9373
rect 2593 9364 2605 9367
rect 2280 9336 2605 9364
rect 2280 9324 2286 9336
rect 2593 9333 2605 9336
rect 2639 9333 2651 9367
rect 3050 9364 3056 9376
rect 3011 9336 3056 9364
rect 2593 9327 2651 9333
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3513 9367 3571 9373
rect 3513 9333 3525 9367
rect 3559 9364 3571 9367
rect 4154 9364 4160 9376
rect 3559 9336 4160 9364
rect 3559 9333 3571 9336
rect 3513 9327 3571 9333
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5828 9364 5856 9395
rect 7006 9392 7012 9404
rect 7064 9392 7070 9444
rect 7392 9441 7420 9472
rect 7193 9435 7251 9441
rect 7193 9401 7205 9435
rect 7239 9401 7251 9435
rect 7193 9395 7251 9401
rect 7377 9435 7435 9441
rect 7377 9401 7389 9435
rect 7423 9401 7435 9435
rect 7377 9395 7435 9401
rect 7469 9435 7527 9441
rect 7469 9401 7481 9435
rect 7515 9432 7527 9435
rect 7558 9432 7564 9444
rect 7515 9404 7564 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 6270 9364 6276 9376
rect 5123 9336 5856 9364
rect 6231 9336 6276 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 6270 9324 6276 9336
rect 6328 9364 6334 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 6328 9336 6377 9364
rect 6328 9324 6334 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6546 9364 6552 9376
rect 6507 9336 6552 9364
rect 6365 9327 6423 9333
rect 6546 9324 6552 9336
rect 6604 9364 6610 9376
rect 7208 9364 7236 9395
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 8956 9441 8984 9540
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9306 9568 9312 9580
rect 9079 9540 9312 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10042 9568 10048 9580
rect 9732 9540 10048 9568
rect 9732 9528 9738 9540
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 10134 9500 10140 9512
rect 10095 9472 10140 9500
rect 10134 9460 10140 9472
rect 10192 9500 10198 9512
rect 10502 9500 10508 9512
rect 10192 9472 10508 9500
rect 10192 9460 10198 9472
rect 10502 9460 10508 9472
rect 10560 9460 10566 9512
rect 10980 9500 11008 9676
rect 11882 9664 11888 9716
rect 11940 9704 11946 9716
rect 11940 9676 12480 9704
rect 11940 9664 11946 9676
rect 11974 9596 11980 9648
rect 12032 9636 12038 9648
rect 12069 9639 12127 9645
rect 12069 9636 12081 9639
rect 12032 9608 12081 9636
rect 12032 9596 12038 9608
rect 12069 9605 12081 9608
rect 12115 9636 12127 9639
rect 12342 9636 12348 9648
rect 12115 9608 12348 9636
rect 12115 9605 12127 9608
rect 12069 9599 12127 9605
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 11422 9568 11428 9580
rect 11383 9540 11428 9568
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 12452 9568 12480 9676
rect 13446 9664 13452 9716
rect 13504 9704 13510 9716
rect 16850 9704 16856 9716
rect 13504 9676 13768 9704
rect 16763 9676 16856 9704
rect 13504 9664 13510 9676
rect 13740 9636 13768 9676
rect 16850 9664 16856 9676
rect 16908 9704 16914 9716
rect 17497 9707 17555 9713
rect 17497 9704 17509 9707
rect 16908 9676 17509 9704
rect 16908 9664 16914 9676
rect 17497 9673 17509 9676
rect 17543 9704 17555 9707
rect 17586 9704 17592 9716
rect 17543 9676 17592 9704
rect 17543 9673 17555 9676
rect 17497 9667 17555 9673
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 18325 9707 18383 9713
rect 18325 9673 18337 9707
rect 18371 9704 18383 9707
rect 19150 9704 19156 9716
rect 18371 9676 19156 9704
rect 18371 9673 18383 9676
rect 18325 9667 18383 9673
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 20530 9664 20536 9716
rect 20588 9664 20594 9716
rect 20898 9704 20904 9716
rect 20859 9676 20904 9704
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 21266 9664 21272 9716
rect 21324 9704 21330 9716
rect 21450 9704 21456 9716
rect 21324 9676 21456 9704
rect 21324 9664 21330 9676
rect 21450 9664 21456 9676
rect 21508 9664 21514 9716
rect 22278 9664 22284 9716
rect 22336 9704 22342 9716
rect 23658 9704 23664 9716
rect 22336 9676 23664 9704
rect 22336 9664 22342 9676
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 24210 9664 24216 9716
rect 24268 9704 24274 9716
rect 24489 9707 24547 9713
rect 24489 9704 24501 9707
rect 24268 9676 24501 9704
rect 24268 9664 24274 9676
rect 24489 9673 24501 9676
rect 24535 9673 24547 9707
rect 24489 9667 24547 9673
rect 13817 9639 13875 9645
rect 13817 9636 13829 9639
rect 13740 9608 13829 9636
rect 13817 9605 13829 9608
rect 13863 9605 13875 9639
rect 13817 9599 13875 9605
rect 14458 9596 14464 9648
rect 14516 9636 14522 9648
rect 14737 9639 14795 9645
rect 14737 9636 14749 9639
rect 14516 9608 14749 9636
rect 14516 9596 14522 9608
rect 14737 9605 14749 9608
rect 14783 9605 14795 9639
rect 14737 9599 14795 9605
rect 16758 9596 16764 9648
rect 16816 9636 16822 9648
rect 17310 9636 17316 9648
rect 16816 9608 17316 9636
rect 16816 9596 16822 9608
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 17770 9636 17776 9648
rect 17731 9608 17776 9636
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 20070 9596 20076 9648
rect 20128 9636 20134 9648
rect 20548 9636 20576 9664
rect 20128 9608 20576 9636
rect 20916 9636 20944 9664
rect 22649 9639 22707 9645
rect 22649 9636 22661 9639
rect 20916 9608 21496 9636
rect 20128 9596 20134 9608
rect 14274 9568 14280 9580
rect 12452 9540 12664 9568
rect 14235 9540 14280 9568
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10980 9472 11161 9500
rect 11149 9469 11161 9472
rect 11195 9500 11207 9503
rect 12342 9500 12348 9512
rect 11195 9472 12348 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 12636 9509 12664 9540
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9469 12679 9503
rect 12621 9463 12679 9469
rect 13170 9460 13176 9512
rect 13228 9500 13234 9512
rect 13633 9503 13691 9509
rect 13633 9500 13645 9503
rect 13228 9472 13645 9500
rect 13228 9460 13234 9472
rect 13633 9469 13645 9472
rect 13679 9500 13691 9503
rect 13814 9500 13820 9512
rect 13679 9472 13820 9500
rect 13679 9469 13691 9472
rect 13633 9463 13691 9469
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 14476 9500 14504 9596
rect 20898 9528 20904 9580
rect 20956 9568 20962 9580
rect 21174 9568 21180 9580
rect 20956 9540 21180 9568
rect 20956 9528 20962 9540
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 21468 9568 21496 9608
rect 21836 9608 22661 9636
rect 21836 9568 21864 9608
rect 22649 9605 22661 9608
rect 22695 9636 22707 9639
rect 22738 9636 22744 9648
rect 22695 9608 22744 9636
rect 22695 9605 22707 9608
rect 22649 9599 22707 9605
rect 22738 9596 22744 9608
rect 22796 9596 22802 9648
rect 23934 9596 23940 9648
rect 23992 9636 23998 9648
rect 25041 9639 25099 9645
rect 25041 9636 25053 9639
rect 23992 9608 25053 9636
rect 23992 9596 23998 9608
rect 25041 9605 25053 9608
rect 25087 9605 25099 9639
rect 25041 9599 25099 9605
rect 21468 9540 21864 9568
rect 21913 9571 21971 9577
rect 21913 9537 21925 9571
rect 21959 9568 21971 9571
rect 23109 9571 23167 9577
rect 21959 9540 22416 9568
rect 21959 9537 21971 9540
rect 21913 9531 21971 9537
rect 14292 9472 14504 9500
rect 15381 9503 15439 9509
rect 8757 9435 8815 9441
rect 8757 9401 8769 9435
rect 8803 9401 8815 9435
rect 8757 9395 8815 9401
rect 8941 9435 8999 9441
rect 8941 9401 8953 9435
rect 8987 9401 8999 9435
rect 8941 9395 8999 9401
rect 9769 9435 9827 9441
rect 9769 9401 9781 9435
rect 9815 9432 9827 9435
rect 10226 9432 10232 9444
rect 9815 9404 10232 9432
rect 9815 9401 9827 9404
rect 9769 9395 9827 9401
rect 6604 9336 7236 9364
rect 8772 9364 8800 9395
rect 10226 9392 10232 9404
rect 10284 9432 10290 9444
rect 10686 9432 10692 9444
rect 10284 9404 10692 9432
rect 10284 9392 10290 9404
rect 10686 9392 10692 9404
rect 10744 9432 10750 9444
rect 14292 9441 14320 9472
rect 15381 9469 15393 9503
rect 15427 9500 15439 9503
rect 15470 9500 15476 9512
rect 15427 9472 15476 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 15562 9460 15568 9512
rect 15620 9500 15626 9512
rect 15729 9503 15787 9509
rect 15729 9500 15741 9503
rect 15620 9472 15741 9500
rect 15620 9460 15626 9472
rect 15729 9469 15741 9472
rect 15775 9469 15787 9503
rect 18785 9503 18843 9509
rect 18785 9500 18797 9503
rect 15729 9463 15787 9469
rect 18616 9472 18797 9500
rect 14277 9435 14335 9441
rect 10744 9404 14228 9432
rect 10744 9392 10750 9404
rect 9398 9364 9404 9376
rect 8772 9336 9404 9364
rect 6604 9324 6610 9336
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 10008 9336 10609 9364
rect 10008 9324 10014 9336
rect 10597 9333 10609 9336
rect 10643 9364 10655 9367
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 10643 9336 11345 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 11333 9333 11345 9336
rect 11379 9364 11391 9367
rect 11606 9364 11612 9376
rect 11379 9336 11612 9364
rect 11379 9333 11391 9336
rect 11333 9327 11391 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 13078 9364 13084 9376
rect 12851 9336 13084 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 13262 9364 13268 9376
rect 13223 9336 13268 9364
rect 13262 9324 13268 9336
rect 13320 9364 13326 9376
rect 13722 9364 13728 9376
rect 13320 9336 13728 9364
rect 13320 9324 13326 9336
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14200 9364 14228 9404
rect 14277 9401 14289 9435
rect 14323 9401 14335 9435
rect 14277 9395 14335 9401
rect 14369 9435 14427 9441
rect 14369 9401 14381 9435
rect 14415 9432 14427 9435
rect 14550 9432 14556 9444
rect 14415 9404 14556 9432
rect 14415 9401 14427 9404
rect 14369 9395 14427 9401
rect 14550 9392 14556 9404
rect 14608 9392 14614 9444
rect 15488 9432 15516 9460
rect 15838 9432 15844 9444
rect 15488 9404 15844 9432
rect 15838 9392 15844 9404
rect 15896 9392 15902 9444
rect 16114 9364 16120 9376
rect 14200 9336 16120 9364
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 18322 9324 18328 9376
rect 18380 9364 18386 9376
rect 18616 9373 18644 9472
rect 18785 9469 18797 9472
rect 18831 9469 18843 9503
rect 18785 9463 18843 9469
rect 19052 9503 19110 9509
rect 19052 9469 19064 9503
rect 19098 9500 19110 9503
rect 19518 9500 19524 9512
rect 19098 9472 19524 9500
rect 19098 9469 19110 9472
rect 19052 9463 19110 9469
rect 19518 9460 19524 9472
rect 19576 9500 19582 9512
rect 20622 9500 20628 9512
rect 19576 9472 20628 9500
rect 19576 9460 19582 9472
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 22388 9509 22416 9540
rect 23109 9537 23121 9571
rect 23155 9568 23167 9571
rect 23290 9568 23296 9580
rect 23155 9540 23296 9568
rect 23155 9537 23167 9540
rect 23109 9531 23167 9537
rect 23290 9528 23296 9540
rect 23348 9568 23354 9580
rect 23348 9540 24256 9568
rect 23348 9528 23354 9540
rect 21637 9503 21695 9509
rect 21637 9469 21649 9503
rect 21683 9500 21695 9503
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 21683 9472 22109 9500
rect 21683 9469 21695 9472
rect 21637 9463 21695 9469
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 22373 9503 22431 9509
rect 22373 9469 22385 9503
rect 22419 9500 22431 9503
rect 23198 9500 23204 9512
rect 22419 9472 23204 9500
rect 22419 9469 22431 9472
rect 22373 9463 22431 9469
rect 23198 9460 23204 9472
rect 23256 9460 23262 9512
rect 23477 9503 23535 9509
rect 23477 9469 23489 9503
rect 23523 9500 23535 9503
rect 23566 9500 23572 9512
rect 23523 9472 23572 9500
rect 23523 9469 23535 9472
rect 23477 9463 23535 9469
rect 23566 9460 23572 9472
rect 23624 9500 23630 9512
rect 24029 9503 24087 9509
rect 24029 9500 24041 9503
rect 23624 9472 24041 9500
rect 23624 9460 23630 9472
rect 24029 9469 24041 9472
rect 24075 9469 24087 9503
rect 24029 9463 24087 9469
rect 20346 9392 20352 9444
rect 20404 9432 20410 9444
rect 24228 9441 24256 9540
rect 24302 9528 24308 9580
rect 24360 9568 24366 9580
rect 24670 9568 24676 9580
rect 24360 9540 24676 9568
rect 24360 9528 24366 9540
rect 24670 9528 24676 9540
rect 24728 9528 24734 9580
rect 25958 9568 25964 9580
rect 25919 9540 25964 9568
rect 25958 9528 25964 9540
rect 26016 9528 26022 9580
rect 25222 9500 25228 9512
rect 25183 9472 25228 9500
rect 25222 9460 25228 9472
rect 25280 9460 25286 9512
rect 21821 9435 21879 9441
rect 20404 9404 21496 9432
rect 20404 9392 20410 9404
rect 18601 9367 18659 9373
rect 18601 9364 18613 9367
rect 18380 9336 18613 9364
rect 18380 9324 18386 9336
rect 18601 9333 18613 9336
rect 18647 9333 18659 9367
rect 18601 9327 18659 9333
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 20165 9367 20223 9373
rect 20165 9364 20177 9367
rect 19024 9336 20177 9364
rect 19024 9324 19030 9336
rect 20165 9333 20177 9336
rect 20211 9333 20223 9367
rect 20165 9327 20223 9333
rect 21174 9324 21180 9376
rect 21232 9364 21238 9376
rect 21343 9367 21401 9373
rect 21343 9364 21355 9367
rect 21232 9336 21355 9364
rect 21232 9324 21238 9336
rect 21343 9333 21355 9336
rect 21389 9333 21401 9367
rect 21468 9364 21496 9404
rect 21821 9401 21833 9435
rect 21867 9432 21879 9435
rect 23735 9435 23793 9441
rect 23735 9432 23747 9435
rect 21867 9404 23747 9432
rect 21867 9401 21879 9404
rect 21821 9395 21879 9401
rect 23735 9401 23747 9404
rect 23781 9401 23793 9435
rect 23735 9395 23793 9401
rect 24213 9435 24271 9441
rect 24213 9401 24225 9435
rect 24259 9401 24271 9435
rect 24213 9395 24271 9401
rect 24305 9435 24363 9441
rect 24305 9401 24317 9435
rect 24351 9401 24363 9435
rect 25498 9432 25504 9444
rect 25459 9404 25504 9432
rect 24305 9395 24363 9401
rect 21836 9364 21864 9395
rect 21468 9336 21864 9364
rect 22097 9367 22155 9373
rect 21343 9327 21401 9333
rect 22097 9333 22109 9367
rect 22143 9364 22155 9367
rect 23106 9364 23112 9376
rect 22143 9336 23112 9364
rect 22143 9333 22155 9336
rect 22097 9327 22155 9333
rect 23106 9324 23112 9336
rect 23164 9324 23170 9376
rect 23566 9324 23572 9376
rect 23624 9364 23630 9376
rect 24320 9364 24348 9395
rect 25498 9392 25504 9404
rect 25556 9392 25562 9444
rect 24489 9367 24547 9373
rect 24489 9364 24501 9367
rect 23624 9336 24501 9364
rect 23624 9324 23630 9336
rect 24489 9333 24501 9336
rect 24535 9364 24547 9367
rect 24673 9367 24731 9373
rect 24673 9364 24685 9367
rect 24535 9336 24685 9364
rect 24535 9333 24547 9336
rect 24489 9327 24547 9333
rect 24673 9333 24685 9336
rect 24719 9333 24731 9367
rect 26326 9364 26332 9376
rect 26287 9336 26332 9364
rect 24673 9327 24731 9333
rect 26326 9324 26332 9336
rect 26384 9324 26390 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2133 9163 2191 9169
rect 2133 9129 2145 9163
rect 2179 9160 2191 9163
rect 2590 9160 2596 9172
rect 2179 9132 2596 9160
rect 2179 9129 2191 9132
rect 2133 9123 2191 9129
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 3697 9163 3755 9169
rect 3697 9129 3709 9163
rect 3743 9160 3755 9163
rect 3878 9160 3884 9172
rect 3743 9132 3884 9160
rect 3743 9129 3755 9132
rect 3697 9123 3755 9129
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4617 9163 4675 9169
rect 4212 9132 4559 9160
rect 4212 9120 4218 9132
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 2038 9092 2044 9104
rect 1636 9064 2044 9092
rect 1636 9052 1642 9064
rect 2038 9052 2044 9064
rect 2096 9052 2102 9104
rect 2961 9095 3019 9101
rect 2961 9092 2973 9095
rect 2792 9064 2973 9092
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 2038 8956 2044 8968
rect 1443 8928 2044 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 2792 8956 2820 9064
rect 2961 9061 2973 9064
rect 3007 9061 3019 9095
rect 4430 9092 4436 9104
rect 4391 9064 4436 9092
rect 2961 9055 3019 9061
rect 4430 9052 4436 9064
rect 4488 9052 4494 9104
rect 4531 9092 4559 9132
rect 4617 9129 4629 9163
rect 4663 9160 4675 9163
rect 4982 9160 4988 9172
rect 4663 9132 4988 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 6178 9160 6184 9172
rect 5592 9132 6184 9160
rect 5592 9120 5598 9132
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 9364 9132 9873 9160
rect 9364 9120 9370 9132
rect 9861 9129 9873 9132
rect 9907 9129 9919 9163
rect 9861 9123 9919 9129
rect 10321 9163 10379 9169
rect 10321 9129 10333 9163
rect 10367 9160 10379 9163
rect 10367 9132 11100 9160
rect 10367 9129 10379 9132
rect 10321 9123 10379 9129
rect 6822 9092 6828 9104
rect 4531 9064 6828 9092
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 10870 9052 10876 9104
rect 10928 9092 10934 9104
rect 11072 9101 11100 9132
rect 11606 9120 11612 9172
rect 11664 9160 11670 9172
rect 11790 9160 11796 9172
rect 11664 9132 11796 9160
rect 11664 9120 11670 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 13357 9163 13415 9169
rect 13357 9129 13369 9163
rect 13403 9160 13415 9163
rect 13538 9160 13544 9172
rect 13403 9132 13544 9160
rect 13403 9129 13415 9132
rect 13357 9123 13415 9129
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 16574 9120 16580 9172
rect 16632 9160 16638 9172
rect 16945 9163 17003 9169
rect 16945 9160 16957 9163
rect 16632 9132 16957 9160
rect 16632 9120 16638 9132
rect 16945 9129 16957 9132
rect 16991 9129 17003 9163
rect 16945 9123 17003 9129
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17497 9163 17555 9169
rect 17497 9160 17509 9163
rect 17184 9132 17509 9160
rect 17184 9120 17190 9132
rect 17497 9129 17509 9132
rect 17543 9129 17555 9163
rect 18414 9160 18420 9172
rect 18375 9132 18420 9160
rect 17497 9123 17555 9129
rect 18414 9120 18420 9132
rect 18472 9120 18478 9172
rect 18782 9120 18788 9172
rect 18840 9120 18846 9172
rect 18966 9120 18972 9172
rect 19024 9160 19030 9172
rect 19518 9160 19524 9172
rect 19024 9132 19196 9160
rect 19479 9132 19524 9160
rect 19024 9120 19030 9132
rect 10965 9095 11023 9101
rect 10965 9092 10977 9095
rect 10928 9064 10977 9092
rect 10928 9052 10934 9064
rect 10965 9061 10977 9064
rect 11011 9061 11023 9095
rect 10965 9055 11023 9061
rect 11057 9095 11115 9101
rect 11057 9061 11069 9095
rect 11103 9092 11115 9095
rect 11330 9092 11336 9104
rect 11103 9064 11336 9092
rect 11103 9061 11115 9064
rect 11057 9055 11115 9061
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 12434 9092 12440 9104
rect 11992 9064 12440 9092
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 9024 3111 9027
rect 5077 9027 5135 9033
rect 5077 9024 5089 9027
rect 3099 8996 5089 9024
rect 3099 8993 3111 8996
rect 3053 8987 3111 8993
rect 5077 8993 5089 8996
rect 5123 9024 5135 9027
rect 5442 9024 5448 9036
rect 5123 8996 5448 9024
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5896 9027 5954 9033
rect 5896 9024 5908 9027
rect 5552 8996 5908 9024
rect 2740 8928 2820 8956
rect 2869 8959 2927 8965
rect 2740 8916 2746 8928
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 5552 8956 5580 8996
rect 5896 8993 5908 8996
rect 5942 9024 5954 9027
rect 6454 9024 6460 9036
rect 5942 8996 6460 9024
rect 5942 8993 5954 8996
rect 5896 8987 5954 8993
rect 6454 8984 6460 8996
rect 6512 9024 6518 9036
rect 7558 9024 7564 9036
rect 6512 8996 7564 9024
rect 6512 8984 6518 8996
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 8478 9024 8484 9036
rect 8439 8996 8484 9024
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 11992 9033 12020 9064
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 15832 9095 15890 9101
rect 15832 9061 15844 9095
rect 15878 9092 15890 9095
rect 16298 9092 16304 9104
rect 15878 9064 16304 9092
rect 15878 9061 15890 9064
rect 15832 9055 15890 9061
rect 16298 9052 16304 9064
rect 16356 9092 16362 9104
rect 16850 9092 16856 9104
rect 16356 9064 16856 9092
rect 16356 9052 16362 9064
rect 16850 9052 16856 9064
rect 16908 9052 16914 9104
rect 18800 9092 18828 9120
rect 19168 9101 19196 9132
rect 19518 9120 19524 9132
rect 19576 9120 19582 9172
rect 20346 9160 20352 9172
rect 20307 9132 20352 9160
rect 20346 9120 20352 9132
rect 20404 9120 20410 9172
rect 21174 9120 21180 9172
rect 21232 9160 21238 9172
rect 21821 9163 21879 9169
rect 21821 9160 21833 9163
rect 21232 9132 21833 9160
rect 21232 9120 21238 9132
rect 21821 9129 21833 9132
rect 21867 9129 21879 9163
rect 21821 9123 21879 9129
rect 22002 9120 22008 9172
rect 22060 9160 22066 9172
rect 22830 9160 22836 9172
rect 22060 9132 22836 9160
rect 22060 9120 22066 9132
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 24581 9163 24639 9169
rect 24581 9160 24593 9163
rect 23532 9132 24593 9160
rect 23532 9120 23538 9132
rect 24581 9129 24593 9132
rect 24627 9129 24639 9163
rect 24581 9123 24639 9129
rect 25317 9163 25375 9169
rect 25317 9129 25329 9163
rect 25363 9160 25375 9163
rect 25866 9160 25872 9172
rect 25363 9132 25872 9160
rect 25363 9129 25375 9132
rect 25317 9123 25375 9129
rect 25866 9120 25872 9132
rect 25924 9120 25930 9172
rect 25958 9120 25964 9172
rect 26016 9160 26022 9172
rect 26142 9160 26148 9172
rect 26016 9132 26148 9160
rect 26016 9120 26022 9132
rect 26142 9120 26148 9132
rect 26200 9120 26206 9172
rect 19061 9095 19119 9101
rect 19061 9092 19073 9095
rect 18800 9064 19073 9092
rect 19061 9061 19073 9064
rect 19107 9061 19119 9095
rect 19061 9055 19119 9061
rect 19153 9095 19211 9101
rect 19153 9061 19165 9095
rect 19199 9061 19211 9095
rect 20714 9092 20720 9104
rect 20675 9064 20720 9092
rect 19153 9055 19211 9061
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 21450 9092 21456 9104
rect 21411 9064 21456 9092
rect 21450 9052 21456 9064
rect 21508 9052 21514 9104
rect 21545 9095 21603 9101
rect 21545 9061 21557 9095
rect 21591 9092 21603 9095
rect 21634 9092 21640 9104
rect 21591 9064 21640 9092
rect 21591 9061 21603 9064
rect 21545 9055 21603 9061
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 12233 9027 12291 9033
rect 12233 9024 12245 9027
rect 12124 8996 12245 9024
rect 12124 8984 12130 8996
rect 12233 8993 12245 8996
rect 12279 9024 12291 9027
rect 15013 9027 15071 9033
rect 15013 9024 15025 9027
rect 12279 8996 15025 9024
rect 12279 8993 12291 8996
rect 12233 8987 12291 8993
rect 15013 8993 15025 8996
rect 15059 9024 15071 9027
rect 15378 9024 15384 9036
rect 15059 8996 15384 9024
rect 15059 8993 15071 8996
rect 15013 8987 15071 8993
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 15562 9024 15568 9036
rect 15475 8996 15568 9024
rect 15562 8984 15568 8996
rect 15620 9024 15626 9036
rect 18322 9024 18328 9036
rect 15620 8996 18328 9024
rect 15620 8984 15626 8996
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 18877 9027 18935 9033
rect 18877 9024 18889 9027
rect 18840 8996 18889 9024
rect 18840 8984 18846 8996
rect 18877 8993 18889 8996
rect 18923 8993 18935 9027
rect 18877 8987 18935 8993
rect 21174 8984 21180 9036
rect 21232 9024 21238 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 21232 8996 21281 9024
rect 21232 8984 21238 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 21269 8987 21327 8993
rect 4755 8928 5580 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 2130 8848 2136 8900
rect 2188 8888 2194 8900
rect 2774 8888 2780 8900
rect 2188 8860 2780 8888
rect 2188 8848 2194 8860
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 2884 8888 2912 8919
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 5684 8928 5729 8956
rect 5684 8916 5690 8928
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 8996 8928 9413 8956
rect 8996 8916 9002 8928
rect 9401 8925 9413 8928
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 11054 8956 11060 8968
rect 11011 8928 11060 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 21560 8956 21588 9055
rect 21634 9052 21640 9064
rect 21692 9092 21698 9104
rect 22094 9092 22100 9104
rect 21692 9064 22100 9092
rect 21692 9052 21698 9064
rect 22094 9052 22100 9064
rect 22152 9052 22158 9104
rect 22557 9095 22615 9101
rect 22557 9061 22569 9095
rect 22603 9092 22615 9095
rect 25682 9092 25688 9104
rect 22603 9064 22876 9092
rect 25643 9064 25688 9092
rect 22603 9061 22615 9064
rect 22557 9055 22615 9061
rect 22649 9027 22707 9033
rect 22649 8993 22661 9027
rect 22695 9024 22707 9027
rect 22738 9024 22744 9036
rect 22695 8996 22744 9024
rect 22695 8993 22707 8996
rect 22649 8987 22707 8993
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 22848 9024 22876 9064
rect 25682 9052 25688 9064
rect 25740 9052 25746 9104
rect 22916 9027 22974 9033
rect 22916 9024 22928 9027
rect 22848 8996 22928 9024
rect 22916 8993 22928 8996
rect 22962 9024 22974 9027
rect 23290 9024 23296 9036
rect 22962 8996 23296 9024
rect 22962 8993 22974 8996
rect 22916 8987 22974 8993
rect 23290 8984 23296 8996
rect 23348 8984 23354 9036
rect 25133 9027 25191 9033
rect 25133 8993 25145 9027
rect 25179 9024 25191 9027
rect 25498 9024 25504 9036
rect 25179 8996 25504 9024
rect 25179 8993 25191 8996
rect 25133 8987 25191 8993
rect 25498 8984 25504 8996
rect 25556 9024 25562 9036
rect 26142 9024 26148 9036
rect 25556 8996 26148 9024
rect 25556 8984 25562 8996
rect 26142 8984 26148 8996
rect 26200 8984 26206 9036
rect 17276 8928 21588 8956
rect 17276 8916 17282 8928
rect 24854 8916 24860 8968
rect 24912 8956 24918 8968
rect 26053 8959 26111 8965
rect 26053 8956 26065 8959
rect 24912 8928 26065 8956
rect 24912 8916 24918 8928
rect 26053 8925 26065 8928
rect 26099 8925 26111 8959
rect 26053 8919 26111 8925
rect 3142 8888 3148 8900
rect 2884 8860 3148 8888
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 4157 8891 4215 8897
rect 4157 8857 4169 8891
rect 4203 8888 4215 8891
rect 4338 8888 4344 8900
rect 4203 8860 4344 8888
rect 4203 8857 4215 8860
rect 4157 8851 4215 8857
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 2280 8792 2513 8820
rect 2280 8780 2286 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 4706 8820 4712 8832
rect 3108 8792 4712 8820
rect 3108 8780 3114 8792
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 5534 8820 5540 8832
rect 5495 8792 5540 8820
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 5644 8820 5672 8916
rect 8665 8891 8723 8897
rect 8665 8857 8677 8891
rect 8711 8888 8723 8891
rect 9306 8888 9312 8900
rect 8711 8860 9312 8888
rect 8711 8857 8723 8860
rect 8665 8851 8723 8857
rect 9306 8848 9312 8860
rect 9364 8848 9370 8900
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 10505 8891 10563 8897
rect 10505 8888 10517 8891
rect 9732 8860 10517 8888
rect 9732 8848 9738 8860
rect 10505 8857 10517 8860
rect 10551 8857 10563 8891
rect 10505 8851 10563 8857
rect 14369 8891 14427 8897
rect 14369 8857 14381 8891
rect 14415 8888 14427 8891
rect 14550 8888 14556 8900
rect 14415 8860 14556 8888
rect 14415 8857 14427 8860
rect 14369 8851 14427 8857
rect 14550 8848 14556 8860
rect 14608 8888 14614 8900
rect 20990 8888 20996 8900
rect 14608 8860 14872 8888
rect 20951 8860 20996 8888
rect 14608 8848 14614 8860
rect 6362 8820 6368 8832
rect 5644 8792 6368 8820
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 7006 8820 7012 8832
rect 6967 8792 7012 8820
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 7926 8820 7932 8832
rect 7887 8792 7932 8820
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 8294 8820 8300 8832
rect 8255 8792 8300 8820
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 8812 8792 9045 8820
rect 8812 8780 8818 8792
rect 9033 8789 9045 8792
rect 9079 8789 9091 8823
rect 9033 8783 9091 8789
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 11388 8792 11437 8820
rect 11388 8780 11394 8792
rect 11425 8789 11437 8792
rect 11471 8789 11483 8823
rect 11790 8820 11796 8832
rect 11751 8792 11796 8820
rect 11425 8783 11483 8789
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 14001 8823 14059 8829
rect 14001 8820 14013 8823
rect 12400 8792 14013 8820
rect 12400 8780 12406 8792
rect 14001 8789 14013 8792
rect 14047 8820 14059 8823
rect 14274 8820 14280 8832
rect 14047 8792 14280 8820
rect 14047 8789 14059 8792
rect 14001 8783 14059 8789
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 14642 8820 14648 8832
rect 14603 8792 14648 8820
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14844 8820 14872 8860
rect 20990 8848 20996 8860
rect 21048 8848 21054 8900
rect 24949 8891 25007 8897
rect 24949 8888 24961 8891
rect 23584 8860 24961 8888
rect 15930 8820 15936 8832
rect 14844 8792 15936 8820
rect 15930 8780 15936 8792
rect 15988 8780 15994 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 17957 8823 18015 8829
rect 17957 8820 17969 8823
rect 17644 8792 17969 8820
rect 17644 8780 17650 8792
rect 17957 8789 17969 8792
rect 18003 8789 18015 8823
rect 17957 8783 18015 8789
rect 18601 8823 18659 8829
rect 18601 8789 18613 8823
rect 18647 8820 18659 8823
rect 19242 8820 19248 8832
rect 18647 8792 19248 8820
rect 18647 8789 18659 8792
rect 18601 8783 18659 8789
rect 19242 8780 19248 8792
rect 19300 8780 19306 8832
rect 19981 8823 20039 8829
rect 19981 8789 19993 8823
rect 20027 8820 20039 8823
rect 21358 8820 21364 8832
rect 20027 8792 21364 8820
rect 20027 8789 20039 8792
rect 19981 8783 20039 8789
rect 21358 8780 21364 8792
rect 21416 8780 21422 8832
rect 21818 8820 21824 8832
rect 21779 8792 21824 8820
rect 21818 8780 21824 8792
rect 21876 8780 21882 8832
rect 22002 8820 22008 8832
rect 21963 8792 22008 8820
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 22554 8780 22560 8832
rect 22612 8820 22618 8832
rect 23584 8820 23612 8860
rect 24949 8857 24961 8860
rect 24995 8857 25007 8891
rect 24949 8851 25007 8857
rect 22612 8792 23612 8820
rect 22612 8780 22618 8792
rect 23934 8780 23940 8832
rect 23992 8820 23998 8832
rect 24029 8823 24087 8829
rect 24029 8820 24041 8823
rect 23992 8792 24041 8820
rect 23992 8780 23998 8792
rect 24029 8789 24041 8792
rect 24075 8789 24087 8823
rect 24029 8783 24087 8789
rect 25590 8780 25596 8832
rect 25648 8820 25654 8832
rect 25866 8820 25872 8832
rect 25648 8792 25872 8820
rect 25648 8780 25654 8792
rect 25866 8780 25872 8792
rect 25924 8780 25930 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2406 8616 2412 8628
rect 2367 8588 2412 8616
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 4246 8616 4252 8628
rect 3835 8588 4252 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 4430 8576 4436 8628
rect 4488 8616 4494 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 4488 8588 5273 8616
rect 4488 8576 4494 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 5261 8579 5319 8585
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 6730 8616 6736 8628
rect 5675 8588 6736 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 6914 8616 6920 8628
rect 6875 8588 6920 8616
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11333 8619 11391 8625
rect 11333 8616 11345 8619
rect 11112 8588 11345 8616
rect 11112 8576 11118 8588
rect 11333 8585 11345 8588
rect 11379 8585 11391 8619
rect 12434 8616 12440 8628
rect 11333 8579 11391 8585
rect 12176 8588 12440 8616
rect 2225 8551 2283 8557
rect 2225 8517 2237 8551
rect 2271 8548 2283 8551
rect 3142 8548 3148 8560
rect 2271 8520 3148 8548
rect 2271 8517 2283 8520
rect 2225 8511 2283 8517
rect 3142 8508 3148 8520
rect 3200 8508 3206 8560
rect 3973 8551 4031 8557
rect 3973 8517 3985 8551
rect 4019 8548 4031 8551
rect 4062 8548 4068 8560
rect 4019 8520 4068 8548
rect 4019 8517 4031 8520
rect 3973 8511 4031 8517
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 4982 8548 4988 8560
rect 4943 8520 4988 8548
rect 4982 8508 4988 8520
rect 5040 8508 5046 8560
rect 6089 8551 6147 8557
rect 6089 8517 6101 8551
rect 6135 8548 6147 8551
rect 6362 8548 6368 8560
rect 6135 8520 6368 8548
rect 6135 8517 6147 8520
rect 6089 8511 6147 8517
rect 6362 8508 6368 8520
rect 6420 8548 6426 8560
rect 8110 8548 8116 8560
rect 6420 8520 8116 8548
rect 6420 8508 6426 8520
rect 8110 8508 8116 8520
rect 8168 8548 8174 8560
rect 8849 8551 8907 8557
rect 8849 8548 8861 8551
rect 8168 8520 8861 8548
rect 8168 8508 8174 8520
rect 8849 8517 8861 8520
rect 8895 8548 8907 8551
rect 8895 8520 9076 8548
rect 8895 8517 8907 8520
rect 8849 8511 8907 8517
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2590 8480 2596 8492
rect 1903 8452 2596 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 2866 8480 2872 8492
rect 2827 8452 2872 8480
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 4614 8480 4620 8492
rect 3467 8452 4620 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 8662 8480 8668 8492
rect 7331 8452 8668 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 9048 8489 9076 8520
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 10100 8452 11161 8480
rect 10100 8440 10106 8452
rect 11149 8449 11161 8452
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 4246 8412 4252 8424
rect 2884 8384 3188 8412
rect 4207 8384 4252 8412
rect 2884 8353 2912 8384
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8313 2927 8347
rect 2869 8307 2927 8313
rect 2961 8347 3019 8353
rect 2961 8313 2973 8347
rect 3007 8344 3019 8347
rect 3050 8344 3056 8356
rect 3007 8316 3056 8344
rect 3007 8313 3019 8316
rect 2961 8307 3019 8313
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 3160 8344 3188 8384
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 5442 8412 5448 8424
rect 5403 8384 5448 8412
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7374 8412 7380 8424
rect 6687 8384 7380 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7374 8372 7380 8384
rect 7432 8412 7438 8424
rect 7469 8415 7527 8421
rect 7469 8412 7481 8415
rect 7432 8384 7481 8412
rect 7432 8372 7438 8384
rect 7469 8381 7481 8384
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 11057 8415 11115 8421
rect 11057 8412 11069 8415
rect 10928 8384 11069 8412
rect 10928 8372 10934 8384
rect 11057 8381 11069 8384
rect 11103 8412 11115 8415
rect 11974 8412 11980 8424
rect 11103 8384 11980 8412
rect 11103 8381 11115 8384
rect 11057 8375 11115 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 3878 8344 3884 8356
rect 3160 8316 3884 8344
rect 3878 8304 3884 8316
rect 3936 8304 3942 8356
rect 4338 8304 4344 8356
rect 4396 8344 4402 8356
rect 4525 8347 4583 8353
rect 4525 8344 4537 8347
rect 4396 8316 4537 8344
rect 4396 8304 4402 8316
rect 4525 8313 4537 8316
rect 4571 8313 4583 8347
rect 4525 8307 4583 8313
rect 4614 8304 4620 8356
rect 4672 8304 4678 8356
rect 7558 8344 7564 8356
rect 7392 8316 7564 8344
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 3786 8276 3792 8288
rect 2648 8248 3792 8276
rect 2648 8236 2654 8248
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4632 8276 4660 8304
rect 7392 8285 7420 8316
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 8018 8344 8024 8356
rect 7975 8316 8024 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8478 8344 8484 8356
rect 8439 8316 8484 8344
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 9214 8304 9220 8356
rect 9272 8353 9278 8356
rect 9272 8347 9336 8353
rect 9272 8313 9290 8347
rect 9324 8313 9336 8347
rect 9272 8307 9336 8313
rect 9272 8304 9278 8307
rect 9398 8304 9404 8356
rect 9456 8344 9462 8356
rect 9674 8344 9680 8356
rect 9456 8316 9680 8344
rect 9456 8304 9462 8316
rect 9674 8304 9680 8316
rect 9732 8304 9738 8356
rect 12176 8353 12204 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 14366 8616 14372 8628
rect 14327 8588 14372 8616
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 15562 8616 15568 8628
rect 15523 8588 15568 8616
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 17034 8616 17040 8628
rect 16995 8588 17040 8616
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 18966 8616 18972 8628
rect 17911 8588 18972 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 19058 8576 19064 8628
rect 19116 8616 19122 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19116 8588 20085 8616
rect 19116 8576 19122 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 21266 8616 21272 8628
rect 21227 8588 21272 8616
rect 20073 8579 20131 8585
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 21358 8576 21364 8628
rect 21416 8616 21422 8628
rect 23106 8616 23112 8628
rect 21416 8588 23112 8616
rect 21416 8576 21422 8588
rect 23106 8576 23112 8588
rect 23164 8616 23170 8628
rect 23753 8619 23811 8625
rect 23753 8616 23765 8619
rect 23164 8588 23765 8616
rect 23164 8576 23170 8588
rect 23753 8585 23765 8588
rect 23799 8585 23811 8619
rect 24670 8616 24676 8628
rect 24631 8588 24676 8616
rect 23753 8579 23811 8585
rect 24670 8576 24676 8588
rect 24728 8576 24734 8628
rect 25869 8619 25927 8625
rect 25869 8585 25881 8619
rect 25915 8616 25927 8619
rect 25958 8616 25964 8628
rect 25915 8588 25964 8616
rect 25915 8585 25927 8588
rect 25869 8579 25927 8585
rect 12452 8489 12480 8576
rect 13814 8548 13820 8560
rect 13727 8520 13820 8548
rect 13814 8508 13820 8520
rect 13872 8548 13878 8560
rect 14550 8548 14556 8560
rect 13872 8520 14556 8548
rect 13872 8508 13878 8520
rect 14550 8508 14556 8520
rect 14608 8508 14614 8560
rect 16666 8548 16672 8560
rect 16627 8520 16672 8548
rect 16666 8508 16672 8520
rect 16724 8508 16730 8560
rect 17402 8548 17408 8560
rect 17363 8520 17408 8548
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 20809 8551 20867 8557
rect 20809 8517 20821 8551
rect 20855 8548 20867 8551
rect 20993 8551 21051 8557
rect 20993 8548 21005 8551
rect 20855 8520 21005 8548
rect 20855 8517 20867 8520
rect 20809 8511 20867 8517
rect 20993 8517 21005 8520
rect 21039 8548 21051 8551
rect 21450 8548 21456 8560
rect 21039 8520 21456 8548
rect 21039 8517 21051 8520
rect 20993 8511 21051 8517
rect 21450 8508 21456 8520
rect 21508 8508 21514 8560
rect 23477 8551 23535 8557
rect 23477 8517 23489 8551
rect 23523 8548 23535 8551
rect 23842 8548 23848 8560
rect 23523 8520 23848 8548
rect 23523 8517 23535 8520
rect 23477 8511 23535 8517
rect 23842 8508 23848 8520
rect 23900 8508 23906 8560
rect 25038 8548 25044 8560
rect 24999 8520 25044 8548
rect 25038 8508 25044 8520
rect 25096 8508 25102 8560
rect 25222 8508 25228 8560
rect 25280 8508 25286 8560
rect 25409 8551 25467 8557
rect 25409 8517 25421 8551
rect 25455 8548 25467 8551
rect 25590 8548 25596 8560
rect 25455 8520 25596 8548
rect 25455 8517 25467 8520
rect 25409 8511 25467 8517
rect 25590 8508 25596 8520
rect 25648 8508 25654 8560
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 16298 8480 16304 8492
rect 15243 8452 16304 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 12452 8412 12480 8443
rect 16298 8440 16304 8452
rect 16356 8440 16362 8492
rect 12986 8412 12992 8424
rect 12452 8384 12992 8412
rect 12986 8372 12992 8384
rect 13044 8372 13050 8424
rect 18322 8372 18328 8424
rect 18380 8412 18386 8424
rect 18966 8421 18972 8424
rect 18693 8415 18751 8421
rect 18693 8412 18705 8415
rect 18380 8384 18705 8412
rect 18380 8372 18386 8384
rect 18693 8381 18705 8384
rect 18739 8381 18751 8415
rect 18960 8412 18972 8421
rect 18927 8384 18972 8412
rect 18693 8375 18751 8381
rect 18960 8375 18972 8384
rect 18966 8372 18972 8375
rect 19024 8372 19030 8424
rect 19242 8372 19248 8424
rect 19300 8412 19306 8424
rect 21545 8415 21603 8421
rect 21545 8412 21557 8415
rect 19300 8384 21557 8412
rect 19300 8372 19306 8384
rect 21545 8381 21557 8384
rect 21591 8412 21603 8415
rect 22189 8415 22247 8421
rect 22189 8412 22201 8415
rect 21591 8384 22201 8412
rect 21591 8381 21603 8384
rect 21545 8375 21603 8381
rect 22189 8381 22201 8384
rect 22235 8412 22247 8415
rect 23014 8412 23020 8424
rect 22235 8384 23020 8412
rect 22235 8381 22247 8384
rect 22189 8375 22247 8381
rect 23014 8372 23020 8384
rect 23072 8372 23078 8424
rect 23860 8412 23888 8508
rect 24670 8440 24676 8492
rect 24728 8480 24734 8492
rect 25240 8480 25268 8508
rect 24728 8452 25268 8480
rect 24728 8440 24734 8452
rect 25225 8415 25283 8421
rect 23860 8384 24256 8412
rect 11793 8347 11851 8353
rect 11793 8344 11805 8347
rect 10980 8316 11805 8344
rect 4479 8248 4660 8276
rect 7377 8279 7435 8285
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 7377 8245 7389 8279
rect 7423 8245 7435 8279
rect 7377 8239 7435 8245
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10413 8279 10471 8285
rect 10413 8276 10425 8279
rect 10192 8248 10425 8276
rect 10192 8236 10198 8248
rect 10413 8245 10425 8248
rect 10459 8245 10471 8279
rect 10413 8239 10471 8245
rect 10870 8236 10876 8288
rect 10928 8276 10934 8288
rect 10980 8276 11008 8316
rect 11793 8313 11805 8316
rect 11839 8344 11851 8347
rect 12161 8347 12219 8353
rect 12161 8344 12173 8347
rect 11839 8316 12173 8344
rect 11839 8313 11851 8316
rect 11793 8307 11851 8313
rect 12161 8313 12173 8316
rect 12207 8313 12219 8347
rect 12161 8307 12219 8313
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 12682 8347 12740 8353
rect 12682 8344 12694 8347
rect 12584 8316 12694 8344
rect 12584 8304 12590 8316
rect 12682 8313 12694 8316
rect 12728 8313 12740 8347
rect 12682 8307 12740 8313
rect 14182 8304 14188 8356
rect 14240 8344 14246 8356
rect 14737 8347 14795 8353
rect 14737 8344 14749 8347
rect 14240 8316 14749 8344
rect 14240 8304 14246 8316
rect 14737 8313 14749 8316
rect 14783 8313 14795 8347
rect 16022 8344 16028 8356
rect 15983 8316 16028 8344
rect 14737 8307 14795 8313
rect 16022 8304 16028 8316
rect 16080 8304 16086 8356
rect 16206 8344 16212 8356
rect 16167 8316 16212 8344
rect 16206 8304 16212 8316
rect 16264 8304 16270 8356
rect 16666 8304 16672 8356
rect 16724 8344 16730 8356
rect 20809 8347 20867 8353
rect 20809 8344 20821 8347
rect 16724 8316 20821 8344
rect 16724 8304 16730 8316
rect 20809 8313 20821 8316
rect 20855 8313 20867 8347
rect 20809 8307 20867 8313
rect 21821 8347 21879 8353
rect 21821 8313 21833 8347
rect 21867 8344 21879 8347
rect 22002 8344 22008 8356
rect 21867 8316 22008 8344
rect 21867 8313 21879 8316
rect 21821 8307 21879 8313
rect 22002 8304 22008 8316
rect 22060 8304 22066 8356
rect 23106 8344 23112 8356
rect 23067 8316 23112 8344
rect 23106 8304 23112 8316
rect 23164 8344 23170 8356
rect 24228 8353 24256 8384
rect 25225 8381 25237 8415
rect 25271 8412 25283 8415
rect 25884 8412 25912 8579
rect 25958 8576 25964 8588
rect 26016 8576 26022 8628
rect 26142 8616 26148 8628
rect 26103 8588 26148 8616
rect 26142 8576 26148 8588
rect 26200 8576 26206 8628
rect 25271 8384 25912 8412
rect 25271 8381 25283 8384
rect 25225 8375 25283 8381
rect 24029 8347 24087 8353
rect 24029 8344 24041 8347
rect 23164 8316 24041 8344
rect 23164 8304 23170 8316
rect 24029 8313 24041 8316
rect 24075 8313 24087 8347
rect 24029 8307 24087 8313
rect 24213 8347 24271 8353
rect 24213 8313 24225 8347
rect 24259 8313 24271 8347
rect 24213 8307 24271 8313
rect 24305 8347 24363 8353
rect 24305 8313 24317 8347
rect 24351 8344 24363 8347
rect 24394 8344 24400 8356
rect 24351 8316 24400 8344
rect 24351 8313 24363 8316
rect 24305 8307 24363 8313
rect 24394 8304 24400 8316
rect 24452 8304 24458 8356
rect 10928 8248 11008 8276
rect 11149 8279 11207 8285
rect 10928 8236 10934 8248
rect 11149 8245 11161 8279
rect 11195 8276 11207 8279
rect 13078 8276 13084 8288
rect 11195 8248 13084 8276
rect 11195 8245 11207 8248
rect 11149 8239 11207 8245
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 18322 8236 18328 8288
rect 18380 8276 18386 8288
rect 18509 8279 18567 8285
rect 18509 8276 18521 8279
rect 18380 8248 18521 8276
rect 18380 8236 18386 8248
rect 18509 8245 18521 8248
rect 18555 8245 18567 8279
rect 18509 8239 18567 8245
rect 21450 8236 21456 8288
rect 21508 8276 21514 8288
rect 21729 8279 21787 8285
rect 21729 8276 21741 8279
rect 21508 8248 21741 8276
rect 21508 8236 21514 8248
rect 21729 8245 21741 8248
rect 21775 8245 21787 8279
rect 21729 8239 21787 8245
rect 22278 8236 22284 8288
rect 22336 8276 22342 8288
rect 22554 8276 22560 8288
rect 22336 8248 22560 8276
rect 22336 8236 22342 8248
rect 22554 8236 22560 8248
rect 22612 8236 22618 8288
rect 22741 8279 22799 8285
rect 22741 8245 22753 8279
rect 22787 8276 22799 8279
rect 23382 8276 23388 8288
rect 22787 8248 23388 8276
rect 22787 8245 22799 8248
rect 22741 8239 22799 8245
rect 23382 8236 23388 8248
rect 23440 8236 23446 8288
rect 23934 8236 23940 8288
rect 23992 8276 23998 8288
rect 24118 8276 24124 8288
rect 23992 8248 24124 8276
rect 23992 8236 23998 8248
rect 24118 8236 24124 8248
rect 24176 8236 24182 8288
rect 25222 8236 25228 8288
rect 25280 8276 25286 8288
rect 25406 8276 25412 8288
rect 25280 8248 25412 8276
rect 25280 8236 25286 8248
rect 25406 8236 25412 8248
rect 25464 8236 25470 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 3050 8072 3056 8084
rect 1995 8044 3056 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 3050 8032 3056 8044
rect 3108 8072 3114 8084
rect 3418 8072 3424 8084
rect 3108 8044 3424 8072
rect 3108 8032 3114 8044
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 5074 8072 5080 8084
rect 5035 8044 5080 8072
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 9125 8075 9183 8081
rect 9125 8041 9137 8075
rect 9171 8072 9183 8075
rect 9214 8072 9220 8084
rect 9171 8044 9220 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 9214 8032 9220 8044
rect 9272 8072 9278 8084
rect 9398 8072 9404 8084
rect 9272 8044 9404 8072
rect 9272 8032 9278 8044
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10042 8072 10048 8084
rect 9916 8044 10048 8072
rect 9916 8032 9922 8044
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 12066 8072 12072 8084
rect 12027 8044 12072 8072
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12526 8072 12532 8084
rect 12487 8044 12532 8072
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 14458 8032 14464 8084
rect 14516 8072 14522 8084
rect 14826 8072 14832 8084
rect 14516 8044 14832 8072
rect 14516 8032 14522 8044
rect 14826 8032 14832 8044
rect 14884 8072 14890 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 15749 8075 15807 8081
rect 15749 8041 15761 8075
rect 15795 8072 15807 8075
rect 16298 8072 16304 8084
rect 15795 8044 16304 8072
rect 15795 8041 15807 8044
rect 15749 8035 15807 8041
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 18966 8072 18972 8084
rect 18927 8044 18972 8072
rect 18966 8032 18972 8044
rect 19024 8032 19030 8084
rect 19334 8072 19340 8084
rect 19295 8044 19340 8072
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19981 8075 20039 8081
rect 19981 8072 19993 8075
rect 19484 8044 19993 8072
rect 19484 8032 19490 8044
rect 19981 8041 19993 8044
rect 20027 8041 20039 8075
rect 19981 8035 20039 8041
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 20901 8075 20959 8081
rect 20901 8072 20913 8075
rect 20864 8044 20913 8072
rect 20864 8032 20870 8044
rect 20901 8041 20913 8044
rect 20947 8041 20959 8075
rect 20901 8035 20959 8041
rect 21266 8032 21272 8084
rect 21324 8072 21330 8084
rect 21729 8075 21787 8081
rect 21729 8072 21741 8075
rect 21324 8044 21741 8072
rect 21324 8032 21330 8044
rect 21729 8041 21741 8044
rect 21775 8041 21787 8075
rect 21729 8035 21787 8041
rect 21818 8032 21824 8084
rect 21876 8072 21882 8084
rect 24210 8072 24216 8084
rect 21876 8044 22508 8072
rect 21876 8032 21882 8044
rect 2958 8004 2964 8016
rect 2919 7976 2964 8004
rect 2958 7964 2964 7976
rect 3016 7964 3022 8016
rect 4430 7964 4436 8016
rect 4488 8004 4494 8016
rect 4617 8007 4675 8013
rect 4617 8004 4629 8007
rect 4488 7976 4629 8004
rect 4488 7964 4494 7976
rect 4617 7973 4629 7976
rect 4663 8004 4675 8007
rect 4890 8004 4896 8016
rect 4663 7976 4896 8004
rect 4663 7973 4675 7976
rect 4617 7967 4675 7973
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 7374 8013 7380 8016
rect 7368 8004 7380 8013
rect 7335 7976 7380 8004
rect 7368 7967 7380 7976
rect 7374 7964 7380 7967
rect 7432 7964 7438 8016
rect 10134 8013 10140 8016
rect 10128 8004 10140 8013
rect 10095 7976 10140 8004
rect 10128 7967 10140 7976
rect 10134 7964 10140 7967
rect 10192 7964 10198 8016
rect 12986 8004 12992 8016
rect 12636 7976 12992 8004
rect 2590 7896 2596 7948
rect 2648 7936 2654 7948
rect 2777 7939 2835 7945
rect 2777 7936 2789 7939
rect 2648 7908 2789 7936
rect 2648 7896 2654 7908
rect 2777 7905 2789 7908
rect 2823 7905 2835 7939
rect 5258 7936 5264 7948
rect 2777 7899 2835 7905
rect 4632 7908 5264 7936
rect 4632 7880 4660 7908
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7936 5871 7939
rect 6822 7936 6828 7948
rect 5859 7908 6828 7936
rect 5859 7905 5871 7908
rect 5813 7899 5871 7905
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 12636 7945 12664 7976
rect 12986 7964 12992 7976
rect 13044 7964 13050 8016
rect 16577 8007 16635 8013
rect 16577 7973 16589 8007
rect 16623 8004 16635 8007
rect 16942 8004 16948 8016
rect 16623 7976 16948 8004
rect 16623 7973 16635 7976
rect 16577 7967 16635 7973
rect 16942 7964 16948 7976
rect 17000 7964 17006 8016
rect 18417 8007 18475 8013
rect 18417 7973 18429 8007
rect 18463 8004 18475 8007
rect 18598 8004 18604 8016
rect 18463 7976 18604 8004
rect 18463 7973 18475 7976
rect 18417 7967 18475 7973
rect 18598 7964 18604 7976
rect 18656 7964 18662 8016
rect 21358 7964 21364 8016
rect 21416 8004 21422 8016
rect 22002 8004 22008 8016
rect 21416 7976 22008 8004
rect 21416 7964 21422 7976
rect 22002 7964 22008 7976
rect 22060 7964 22066 8016
rect 22186 8013 22192 8016
rect 22180 8004 22192 8013
rect 22147 7976 22192 8004
rect 22180 7967 22192 7976
rect 22186 7964 22192 7967
rect 22244 7964 22250 8016
rect 22480 8004 22508 8044
rect 23400 8044 24216 8072
rect 23400 8004 23428 8044
rect 24210 8032 24216 8044
rect 24268 8032 24274 8084
rect 24854 8032 24860 8084
rect 24912 8072 24918 8084
rect 24949 8075 25007 8081
rect 24949 8072 24961 8075
rect 24912 8044 24961 8072
rect 24912 8032 24918 8044
rect 24949 8041 24961 8044
rect 24995 8041 25007 8075
rect 24949 8035 25007 8041
rect 25682 8032 25688 8084
rect 25740 8072 25746 8084
rect 25777 8075 25835 8081
rect 25777 8072 25789 8075
rect 25740 8044 25789 8072
rect 25740 8032 25746 8044
rect 25777 8041 25789 8044
rect 25823 8041 25835 8075
rect 26234 8072 26240 8084
rect 26195 8044 26240 8072
rect 25777 8035 25835 8041
rect 26234 8032 26240 8044
rect 26292 8032 26298 8084
rect 22480 7976 23428 8004
rect 23750 7964 23756 8016
rect 23808 8004 23814 8016
rect 24302 8004 24308 8016
rect 23808 7976 24308 8004
rect 23808 7964 23814 7976
rect 24302 7964 24308 7976
rect 24360 7964 24366 8016
rect 25406 8004 25412 8016
rect 25367 7976 25412 8004
rect 25406 7964 25412 7976
rect 25464 7964 25470 8016
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7905 12679 7939
rect 12888 7939 12946 7945
rect 12888 7936 12900 7939
rect 12621 7899 12679 7905
rect 12728 7908 12900 7936
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 4614 7868 4620 7880
rect 4575 7840 4620 7868
rect 3053 7831 3111 7837
rect 2501 7803 2559 7809
rect 2501 7769 2513 7803
rect 2547 7800 2559 7803
rect 2774 7800 2780 7812
rect 2547 7772 2780 7800
rect 2547 7769 2559 7772
rect 2501 7763 2559 7769
rect 2774 7760 2780 7772
rect 2832 7760 2838 7812
rect 2317 7735 2375 7741
rect 2317 7701 2329 7735
rect 2363 7732 2375 7735
rect 2406 7732 2412 7744
rect 2363 7704 2412 7732
rect 2363 7701 2375 7704
rect 2317 7695 2375 7701
rect 2406 7692 2412 7704
rect 2464 7732 2470 7744
rect 3068 7732 3096 7831
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6638 7868 6644 7880
rect 6135 7840 6644 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 3970 7760 3976 7812
rect 4028 7800 4034 7812
rect 4157 7803 4215 7809
rect 4157 7800 4169 7803
rect 4028 7772 4169 7800
rect 4028 7760 4034 7772
rect 4157 7769 4169 7772
rect 4203 7769 4215 7803
rect 4157 7763 4215 7769
rect 3510 7732 3516 7744
rect 2464 7704 3096 7732
rect 3471 7704 3516 7732
rect 2464 7692 2470 7704
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 4338 7732 4344 7744
rect 3927 7704 4344 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 4338 7692 4344 7704
rect 4396 7732 4402 7744
rect 4724 7732 4752 7831
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 9858 7868 9864 7880
rect 9819 7840 9864 7868
rect 7101 7831 7159 7837
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 7116 7800 7144 7831
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 12728 7868 12756 7908
rect 12888 7905 12900 7908
rect 12934 7936 12946 7939
rect 13722 7936 13728 7948
rect 12934 7908 13728 7936
rect 12934 7905 12946 7908
rect 12888 7899 12946 7905
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 18509 7939 18567 7945
rect 18509 7936 18521 7939
rect 17920 7908 18521 7936
rect 17920 7896 17926 7908
rect 18509 7905 18521 7908
rect 18555 7905 18567 7939
rect 19426 7936 19432 7948
rect 19387 7908 19432 7936
rect 18509 7899 18567 7905
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 20717 7939 20775 7945
rect 20717 7905 20729 7939
rect 20763 7936 20775 7939
rect 21634 7936 21640 7948
rect 20763 7908 21640 7936
rect 20763 7905 20775 7908
rect 20717 7899 20775 7905
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 23566 7896 23572 7948
rect 23624 7936 23630 7948
rect 23845 7939 23903 7945
rect 23845 7936 23857 7939
rect 23624 7908 23857 7936
rect 23624 7896 23630 7908
rect 23845 7905 23857 7908
rect 23891 7936 23903 7939
rect 24394 7936 24400 7948
rect 23891 7908 24400 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24394 7896 24400 7908
rect 24452 7896 24458 7948
rect 12308 7840 12756 7868
rect 16577 7871 16635 7877
rect 12308 7828 12314 7840
rect 16577 7837 16589 7871
rect 16623 7837 16635 7871
rect 16577 7831 16635 7837
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7868 16727 7871
rect 17586 7868 17592 7880
rect 16715 7840 17592 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 11238 7800 11244 7812
rect 6420 7772 7144 7800
rect 11151 7772 11244 7800
rect 6420 7760 6426 7772
rect 11238 7760 11244 7772
rect 11296 7800 11302 7812
rect 12526 7800 12532 7812
rect 11296 7772 12532 7800
rect 11296 7760 11302 7772
rect 12526 7760 12532 7772
rect 12584 7760 12590 7812
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 14001 7803 14059 7809
rect 14001 7800 14013 7803
rect 13872 7772 14013 7800
rect 13872 7760 13878 7772
rect 14001 7769 14013 7772
rect 14047 7800 14059 7803
rect 14918 7800 14924 7812
rect 14047 7772 14924 7800
rect 14047 7769 14059 7772
rect 14001 7763 14059 7769
rect 14918 7760 14924 7772
rect 14976 7760 14982 7812
rect 16592 7800 16620 7831
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 18414 7868 18420 7880
rect 18375 7840 18420 7868
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 21818 7828 21824 7880
rect 21876 7868 21882 7880
rect 21913 7871 21971 7877
rect 21913 7868 21925 7871
rect 21876 7840 21925 7868
rect 21876 7828 21882 7840
rect 21913 7837 21925 7840
rect 21959 7837 21971 7871
rect 24854 7868 24860 7880
rect 24815 7840 24860 7868
rect 21913 7831 21971 7837
rect 24854 7828 24860 7840
rect 24912 7828 24918 7880
rect 25041 7871 25099 7877
rect 25041 7837 25053 7871
rect 25087 7837 25099 7871
rect 25041 7831 25099 7837
rect 16850 7800 16856 7812
rect 16592 7772 16856 7800
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 19613 7803 19671 7809
rect 19613 7769 19625 7803
rect 19659 7800 19671 7803
rect 21174 7800 21180 7812
rect 19659 7772 21180 7800
rect 19659 7769 19671 7772
rect 19613 7763 19671 7769
rect 21174 7760 21180 7772
rect 21232 7760 21238 7812
rect 23198 7800 23204 7812
rect 23124 7772 23204 7800
rect 4396 7704 4752 7732
rect 4396 7692 4402 7704
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 5629 7735 5687 7741
rect 5629 7732 5641 7735
rect 5592 7704 5641 7732
rect 5592 7692 5598 7704
rect 5629 7701 5641 7704
rect 5675 7732 5687 7735
rect 6454 7732 6460 7744
rect 5675 7704 6460 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 6914 7732 6920 7744
rect 6875 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8481 7735 8539 7741
rect 8481 7732 8493 7735
rect 8352 7704 8493 7732
rect 8352 7692 8358 7704
rect 8481 7701 8493 7704
rect 8527 7701 8539 7735
rect 8481 7695 8539 7701
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 8720 7704 9413 7732
rect 8720 7692 8726 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 11698 7732 11704 7744
rect 11204 7704 11704 7732
rect 11204 7692 11210 7704
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14148 7704 14657 7732
rect 14148 7692 14154 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 16114 7732 16120 7744
rect 16075 7704 16120 7732
rect 14645 7695 14703 7701
rect 16114 7692 16120 7704
rect 16172 7692 16178 7744
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 17037 7735 17095 7741
rect 17037 7732 17049 7735
rect 16632 7704 17049 7732
rect 16632 7692 16638 7704
rect 17037 7701 17049 7704
rect 17083 7701 17095 7735
rect 17402 7732 17408 7744
rect 17363 7704 17408 7732
rect 17037 7695 17095 7701
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 17957 7735 18015 7741
rect 17957 7701 17969 7735
rect 18003 7732 18015 7735
rect 18506 7732 18512 7744
rect 18003 7704 18512 7732
rect 18003 7701 18015 7704
rect 17957 7695 18015 7701
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 21450 7732 21456 7744
rect 21411 7704 21456 7732
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 21634 7692 21640 7744
rect 21692 7732 21698 7744
rect 23124 7732 23152 7772
rect 23198 7760 23204 7772
rect 23256 7800 23262 7812
rect 23256 7772 23520 7800
rect 23256 7760 23262 7772
rect 23290 7732 23296 7744
rect 21692 7704 23152 7732
rect 23251 7704 23296 7732
rect 21692 7692 21698 7704
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 23492 7732 23520 7772
rect 24118 7760 24124 7812
rect 24176 7800 24182 7812
rect 24489 7803 24547 7809
rect 24489 7800 24501 7803
rect 24176 7772 24501 7800
rect 24176 7760 24182 7772
rect 24489 7769 24501 7772
rect 24535 7769 24547 7803
rect 24489 7763 24547 7769
rect 24670 7732 24676 7744
rect 23492 7704 24676 7732
rect 24670 7692 24676 7704
rect 24728 7732 24734 7744
rect 25056 7732 25084 7831
rect 24728 7704 25084 7732
rect 24728 7692 24734 7704
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 2958 7528 2964 7540
rect 2271 7500 2964 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 4890 7528 4896 7540
rect 4851 7500 4896 7528
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 6362 7528 6368 7540
rect 6319 7500 6368 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 6362 7488 6368 7500
rect 6420 7528 6426 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6420 7500 6561 7528
rect 6420 7488 6426 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 4338 7352 4344 7404
rect 4396 7392 4402 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 4396 7364 5457 7392
rect 4396 7352 4402 7364
rect 5445 7361 5457 7364
rect 5491 7392 5503 7395
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5491 7364 5825 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 6564 7392 6592 7491
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 9401 7531 9459 7537
rect 9401 7528 9413 7531
rect 8536 7500 9413 7528
rect 8536 7488 8542 7500
rect 9401 7497 9413 7500
rect 9447 7497 9459 7531
rect 9401 7491 9459 7497
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10689 7531 10747 7537
rect 10689 7528 10701 7531
rect 10192 7500 10701 7528
rect 10192 7488 10198 7500
rect 10689 7497 10701 7500
rect 10735 7528 10747 7531
rect 10778 7528 10784 7540
rect 10735 7500 10784 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 11054 7528 11060 7540
rect 11015 7500 11060 7528
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 11606 7488 11612 7540
rect 11664 7528 11670 7540
rect 11882 7528 11888 7540
rect 11664 7500 11888 7528
rect 11664 7488 11670 7500
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12894 7488 12900 7540
rect 12952 7528 12958 7540
rect 13722 7528 13728 7540
rect 12952 7500 13728 7528
rect 12952 7488 12958 7500
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16393 7531 16451 7537
rect 16393 7528 16405 7531
rect 15988 7500 16405 7528
rect 15988 7488 15994 7500
rect 16393 7497 16405 7500
rect 16439 7497 16451 7531
rect 16942 7528 16948 7540
rect 16903 7500 16948 7528
rect 16393 7491 16451 7497
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 18230 7528 18236 7540
rect 18191 7500 18236 7528
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 18690 7528 18696 7540
rect 18651 7500 18696 7528
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 21082 7528 21088 7540
rect 21043 7500 21088 7528
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 21726 7528 21732 7540
rect 21687 7500 21732 7528
rect 21726 7488 21732 7500
rect 21784 7488 21790 7540
rect 22186 7488 22192 7540
rect 22244 7528 22250 7540
rect 22554 7528 22560 7540
rect 22244 7500 22560 7528
rect 22244 7488 22250 7500
rect 22554 7488 22560 7500
rect 22612 7488 22618 7540
rect 22738 7528 22744 7540
rect 22699 7500 22744 7528
rect 22738 7488 22744 7500
rect 22796 7528 22802 7540
rect 23474 7528 23480 7540
rect 22796 7500 23336 7528
rect 23435 7500 23480 7528
rect 22796 7488 22802 7500
rect 9858 7420 9864 7472
rect 9916 7460 9922 7472
rect 10321 7463 10379 7469
rect 10321 7460 10333 7463
rect 9916 7432 10333 7460
rect 9916 7420 9922 7432
rect 10321 7429 10333 7432
rect 10367 7460 10379 7463
rect 10870 7460 10876 7472
rect 10367 7432 10876 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 10870 7420 10876 7432
rect 10928 7420 10934 7472
rect 12986 7460 12992 7472
rect 12947 7432 12992 7460
rect 12986 7420 12992 7432
rect 13044 7420 13050 7472
rect 13538 7460 13544 7472
rect 13499 7432 13544 7460
rect 13538 7420 13544 7432
rect 13596 7420 13602 7472
rect 18322 7420 18328 7472
rect 18380 7460 18386 7472
rect 18969 7463 19027 7469
rect 18969 7460 18981 7463
rect 18380 7432 18981 7460
rect 18380 7420 18386 7432
rect 18969 7429 18981 7432
rect 19015 7460 19027 7463
rect 21100 7460 21128 7488
rect 22002 7460 22008 7472
rect 19015 7432 19196 7460
rect 21100 7432 22008 7460
rect 19015 7429 19027 7432
rect 18969 7423 19027 7429
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 6564 7364 6837 7392
rect 5813 7355 5871 7361
rect 6825 7361 6837 7364
rect 6871 7361 6883 7395
rect 9214 7392 9220 7404
rect 9127 7364 9220 7392
rect 6825 7355 6883 7361
rect 9214 7352 9220 7364
rect 9272 7392 9278 7404
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9272 7364 9965 7392
rect 9272 7352 9278 7364
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 13004 7392 13032 7420
rect 19168 7401 19196 7432
rect 22002 7420 22008 7432
rect 22060 7460 22066 7472
rect 23308 7460 23336 7500
rect 23474 7488 23480 7500
rect 23532 7528 23538 7540
rect 24670 7528 24676 7540
rect 23532 7500 24348 7528
rect 24631 7500 24676 7528
rect 23532 7488 23538 7500
rect 23382 7460 23388 7472
rect 22060 7432 22324 7460
rect 23308 7432 23388 7460
rect 22060 7420 22066 7432
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 12492 7364 12537 7392
rect 13004 7364 14841 7392
rect 12492 7352 12498 7364
rect 14829 7361 14841 7364
rect 14875 7392 14887 7395
rect 15013 7395 15071 7401
rect 15013 7392 15025 7395
rect 14875 7364 15025 7392
rect 14875 7361 14887 7364
rect 14829 7355 14887 7361
rect 15013 7361 15025 7364
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 19153 7395 19211 7401
rect 19153 7361 19165 7395
rect 19199 7361 19211 7395
rect 19153 7355 19211 7361
rect 20346 7352 20352 7404
rect 20404 7392 20410 7404
rect 22296 7401 22324 7432
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 23566 7420 23572 7472
rect 23624 7460 23630 7472
rect 23753 7463 23811 7469
rect 23753 7460 23765 7463
rect 23624 7432 23765 7460
rect 23624 7420 23630 7432
rect 23753 7429 23765 7432
rect 23799 7429 23811 7463
rect 23753 7423 23811 7429
rect 21453 7395 21511 7401
rect 21453 7392 21465 7395
rect 20404 7364 21465 7392
rect 20404 7352 20410 7364
rect 21453 7361 21465 7364
rect 21499 7392 21511 7395
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 21499 7364 22109 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 24210 7392 24216 7404
rect 24171 7364 24216 7392
rect 22281 7355 22339 7361
rect 24210 7352 24216 7364
rect 24268 7352 24274 7404
rect 24320 7401 24348 7500
rect 24670 7488 24676 7500
rect 24728 7488 24734 7540
rect 24946 7488 24952 7540
rect 25004 7528 25010 7540
rect 25041 7531 25099 7537
rect 25041 7528 25053 7531
rect 25004 7500 25053 7528
rect 25004 7488 25010 7500
rect 25041 7497 25053 7500
rect 25087 7497 25099 7531
rect 25041 7491 25099 7497
rect 25409 7531 25467 7537
rect 25409 7497 25421 7531
rect 25455 7528 25467 7531
rect 25774 7528 25780 7540
rect 25455 7500 25780 7528
rect 25455 7497 25467 7500
rect 25409 7491 25467 7497
rect 25774 7488 25780 7500
rect 25832 7488 25838 7540
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 26237 7395 26295 7401
rect 26237 7392 26249 7395
rect 24305 7355 24363 7361
rect 25148 7364 26249 7392
rect 1854 7324 1860 7336
rect 1767 7296 1860 7324
rect 1854 7284 1860 7296
rect 1912 7324 1918 7336
rect 2317 7327 2375 7333
rect 2317 7324 2329 7327
rect 1912 7296 2329 7324
rect 1912 7284 1918 7296
rect 2317 7293 2329 7296
rect 2363 7324 2375 7327
rect 2363 7296 2728 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 2700 7268 2728 7296
rect 3970 7284 3976 7336
rect 4028 7324 4034 7336
rect 4614 7324 4620 7336
rect 4028 7296 4620 7324
rect 4028 7284 4034 7296
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 5132 7296 5181 7324
rect 5132 7284 5138 7296
rect 5169 7293 5181 7296
rect 5215 7293 5227 7327
rect 5169 7287 5227 7293
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7092 7327 7150 7333
rect 7092 7324 7104 7327
rect 6972 7296 7104 7324
rect 6972 7284 6978 7296
rect 7092 7293 7104 7296
rect 7138 7324 7150 7327
rect 8202 7324 8208 7336
rect 7138 7296 8208 7324
rect 7138 7293 7150 7296
rect 7092 7287 7150 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 9677 7327 9735 7333
rect 9677 7293 9689 7327
rect 9723 7324 9735 7327
rect 9766 7324 9772 7336
rect 9723 7296 9772 7324
rect 9723 7293 9735 7296
rect 9677 7287 9735 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 11229 7327 11287 7333
rect 11229 7324 11241 7327
rect 10468 7296 11241 7324
rect 10468 7284 10474 7296
rect 1670 7216 1676 7268
rect 1728 7256 1734 7268
rect 2406 7256 2412 7268
rect 1728 7228 2412 7256
rect 1728 7216 1734 7228
rect 2406 7216 2412 7228
rect 2464 7256 2470 7268
rect 2562 7259 2620 7265
rect 2562 7256 2574 7259
rect 2464 7228 2574 7256
rect 2464 7216 2470 7228
rect 2562 7225 2574 7228
rect 2608 7225 2620 7259
rect 2562 7219 2620 7225
rect 2682 7216 2688 7268
rect 2740 7216 2746 7268
rect 4154 7216 4160 7268
rect 4212 7256 4218 7268
rect 5353 7259 5411 7265
rect 5353 7256 5365 7259
rect 4212 7228 5365 7256
rect 4212 7216 4218 7228
rect 5353 7225 5365 7228
rect 5399 7225 5411 7259
rect 5353 7219 5411 7225
rect 9861 7259 9919 7265
rect 9861 7225 9873 7259
rect 9907 7256 9919 7259
rect 10042 7256 10048 7268
rect 9907 7228 10048 7256
rect 9907 7225 9919 7228
rect 9861 7219 9919 7225
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 11164 7256 11192 7296
rect 11229 7293 11241 7296
rect 11275 7293 11287 7327
rect 11229 7287 11287 7293
rect 13998 7284 14004 7336
rect 14056 7324 14062 7336
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 14056 7296 14105 7324
rect 14056 7284 14062 7296
rect 14093 7293 14105 7296
rect 14139 7324 14151 7327
rect 14366 7324 14372 7336
rect 14139 7296 14372 7324
rect 14139 7293 14151 7296
rect 14093 7287 14151 7293
rect 14366 7284 14372 7296
rect 14424 7284 14430 7336
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7324 18107 7327
rect 18690 7324 18696 7336
rect 18095 7296 18696 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18690 7284 18696 7296
rect 18748 7284 18754 7336
rect 19242 7284 19248 7336
rect 19300 7324 19306 7336
rect 21818 7324 21824 7336
rect 19300 7296 21824 7324
rect 19300 7284 19306 7296
rect 21818 7284 21824 7296
rect 21876 7284 21882 7336
rect 23109 7327 23167 7333
rect 23109 7293 23121 7327
rect 23155 7324 23167 7327
rect 23155 7296 24164 7324
rect 23155 7293 23167 7296
rect 23109 7287 23167 7293
rect 24136 7268 24164 7296
rect 11885 7259 11943 7265
rect 11885 7256 11897 7259
rect 11164 7228 11897 7256
rect 11885 7225 11897 7228
rect 11931 7256 11943 7259
rect 12250 7256 12256 7268
rect 11931 7228 12256 7256
rect 11931 7225 11943 7228
rect 11885 7219 11943 7225
rect 12250 7216 12256 7228
rect 12308 7216 12314 7268
rect 13817 7259 13875 7265
rect 13817 7225 13829 7259
rect 13863 7256 13875 7259
rect 13863 7228 14596 7256
rect 13863 7225 13875 7228
rect 13817 7219 13875 7225
rect 3050 7148 3056 7200
rect 3108 7188 3114 7200
rect 3418 7188 3424 7200
rect 3108 7160 3424 7188
rect 3108 7148 3114 7160
rect 3418 7148 3424 7160
rect 3476 7188 3482 7200
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 3476 7160 3709 7188
rect 3476 7148 3482 7160
rect 3697 7157 3709 7160
rect 3743 7157 3755 7191
rect 3697 7151 3755 7157
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4430 7188 4436 7200
rect 4387 7160 4436 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 8205 7191 8263 7197
rect 8205 7188 8217 7191
rect 7432 7160 8217 7188
rect 7432 7148 7438 7160
rect 8205 7157 8217 7160
rect 8251 7157 8263 7191
rect 8205 7151 8263 7157
rect 8849 7191 8907 7197
rect 8849 7157 8861 7191
rect 8895 7188 8907 7191
rect 9674 7188 9680 7200
rect 8895 7160 9680 7188
rect 8895 7157 8907 7160
rect 8849 7151 8907 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 11425 7191 11483 7197
rect 11425 7157 11437 7191
rect 11471 7188 11483 7191
rect 11698 7188 11704 7200
rect 11471 7160 11704 7188
rect 11471 7157 11483 7160
rect 11425 7151 11483 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 13357 7191 13415 7197
rect 13357 7157 13369 7191
rect 13403 7188 13415 7191
rect 13538 7188 13544 7200
rect 13403 7160 13544 7188
rect 13403 7157 13415 7160
rect 13357 7151 13415 7157
rect 13538 7148 13544 7160
rect 13596 7188 13602 7200
rect 14568 7197 14596 7228
rect 15194 7216 15200 7268
rect 15252 7265 15258 7268
rect 15252 7259 15316 7265
rect 15252 7225 15270 7259
rect 15304 7225 15316 7259
rect 15252 7219 15316 7225
rect 15252 7216 15258 7219
rect 17770 7216 17776 7268
rect 17828 7256 17834 7268
rect 18322 7256 18328 7268
rect 17828 7228 18328 7256
rect 17828 7216 17834 7228
rect 18322 7216 18328 7228
rect 18380 7216 18386 7268
rect 19058 7216 19064 7268
rect 19116 7256 19122 7268
rect 19398 7259 19456 7265
rect 19398 7256 19410 7259
rect 19116 7228 19410 7256
rect 19116 7216 19122 7228
rect 19398 7225 19410 7228
rect 19444 7225 19456 7259
rect 22186 7256 22192 7268
rect 22099 7228 22192 7256
rect 19398 7219 19456 7225
rect 22186 7216 22192 7228
rect 22244 7256 22250 7268
rect 22244 7228 23428 7256
rect 22244 7216 22250 7228
rect 14001 7191 14059 7197
rect 14001 7188 14013 7191
rect 13596 7160 14013 7188
rect 13596 7148 13602 7160
rect 14001 7157 14013 7160
rect 14047 7157 14059 7191
rect 14001 7151 14059 7157
rect 14553 7191 14611 7197
rect 14553 7157 14565 7191
rect 14599 7188 14611 7191
rect 15102 7188 15108 7200
rect 14599 7160 15108 7188
rect 14599 7157 14611 7160
rect 14553 7151 14611 7157
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 16666 7188 16672 7200
rect 15436 7160 16672 7188
rect 15436 7148 15442 7160
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 17405 7191 17463 7197
rect 17405 7157 17417 7191
rect 17451 7188 17463 7191
rect 17586 7188 17592 7200
rect 17451 7160 17592 7188
rect 17451 7157 17463 7160
rect 17405 7151 17463 7157
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 17862 7188 17868 7200
rect 17823 7160 17868 7188
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 20533 7191 20591 7197
rect 20533 7188 20545 7191
rect 20312 7160 20545 7188
rect 20312 7148 20318 7160
rect 20533 7157 20545 7160
rect 20579 7157 20591 7191
rect 23400 7188 23428 7228
rect 24118 7216 24124 7268
rect 24176 7256 24182 7268
rect 24213 7259 24271 7265
rect 24213 7256 24225 7259
rect 24176 7228 24225 7256
rect 24176 7216 24182 7228
rect 24213 7225 24225 7228
rect 24259 7225 24271 7259
rect 25148 7256 25176 7364
rect 26237 7361 26249 7364
rect 26283 7361 26295 7395
rect 26237 7355 26295 7361
rect 25225 7327 25283 7333
rect 25225 7293 25237 7327
rect 25271 7324 25283 7327
rect 25271 7296 25544 7324
rect 25271 7293 25283 7296
rect 25225 7287 25283 7293
rect 24213 7219 24271 7225
rect 24596 7228 25176 7256
rect 24596 7188 24624 7228
rect 25516 7200 25544 7296
rect 23400 7160 24624 7188
rect 20533 7151 20591 7157
rect 25498 7148 25504 7200
rect 25556 7188 25562 7200
rect 25777 7191 25835 7197
rect 25777 7188 25789 7191
rect 25556 7160 25789 7188
rect 25556 7148 25562 7160
rect 25777 7157 25789 7160
rect 25823 7157 25835 7191
rect 25777 7151 25835 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 3786 6944 3792 6996
rect 3844 6984 3850 6996
rect 3844 6956 6960 6984
rect 3844 6944 3850 6956
rect 2961 6919 3019 6925
rect 2961 6885 2973 6919
rect 3007 6885 3019 6919
rect 4890 6916 4896 6928
rect 2961 6879 3019 6885
rect 4080 6888 4896 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 1443 6820 2329 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2317 6817 2329 6820
rect 2363 6848 2375 6851
rect 2590 6848 2596 6860
rect 2363 6820 2596 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 2590 6808 2596 6820
rect 2648 6808 2654 6860
rect 2976 6848 3004 6879
rect 4080 6848 4108 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 5261 6919 5319 6925
rect 5261 6885 5273 6919
rect 5307 6885 5319 6919
rect 5261 6879 5319 6885
rect 6825 6919 6883 6925
rect 6825 6885 6837 6919
rect 6871 6885 6883 6919
rect 6932 6916 6960 6956
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 7653 6987 7711 6993
rect 7653 6984 7665 6987
rect 7432 6956 7665 6984
rect 7432 6944 7438 6956
rect 7653 6953 7665 6956
rect 7699 6953 7711 6987
rect 7653 6947 7711 6953
rect 8389 6987 8447 6993
rect 8389 6953 8401 6987
rect 8435 6984 8447 6987
rect 8570 6984 8576 6996
rect 8435 6956 8576 6984
rect 8435 6953 8447 6956
rect 8389 6947 8447 6953
rect 8570 6944 8576 6956
rect 8628 6944 8634 6996
rect 9692 6956 11376 6984
rect 9692 6916 9720 6956
rect 6932 6888 9720 6916
rect 10229 6919 10287 6925
rect 6825 6879 6883 6885
rect 10229 6885 10241 6919
rect 10275 6885 10287 6919
rect 11238 6916 11244 6928
rect 10229 6879 10287 6885
rect 11164 6888 11244 6916
rect 2976 6820 4108 6848
rect 5276 6848 5304 6879
rect 5442 6848 5448 6860
rect 5276 6820 5448 6848
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 6362 6808 6368 6860
rect 6420 6848 6426 6860
rect 6840 6848 6868 6879
rect 6420 6820 6868 6848
rect 7377 6851 7435 6857
rect 6420 6808 6426 6820
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7466 6848 7472 6860
rect 7423 6820 7472 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8260 6820 8524 6848
rect 8260 6808 8266 6820
rect 8496 6792 8524 6820
rect 10042 6808 10048 6860
rect 10100 6848 10106 6860
rect 10244 6848 10272 6879
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 10100 6820 11069 6848
rect 10100 6808 10106 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 2866 6780 2872 6792
rect 2827 6752 2872 6780
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 3050 6780 3056 6792
rect 3011 6752 3056 6780
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 5258 6780 5264 6792
rect 5219 6752 5264 6780
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5534 6780 5540 6792
rect 5399 6752 5540 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 6454 6780 6460 6792
rect 5859 6752 6460 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6749 6791 6783
rect 6733 6743 6791 6749
rect 2130 6672 2136 6724
rect 2188 6712 2194 6724
rect 2498 6712 2504 6724
rect 2188 6684 2504 6712
rect 2188 6672 2194 6684
rect 2498 6672 2504 6684
rect 2556 6672 2562 6724
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 1857 6647 1915 6653
rect 1857 6644 1869 6647
rect 1728 6616 1869 6644
rect 1728 6604 1734 6616
rect 1857 6613 1869 6616
rect 1903 6613 1915 6647
rect 1857 6607 1915 6613
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 2648 6616 3433 6644
rect 2648 6604 2654 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 3881 6647 3939 6653
rect 3881 6613 3893 6647
rect 3927 6644 3939 6647
rect 4062 6644 4068 6656
rect 3927 6616 4068 6644
rect 3927 6613 3939 6616
rect 3881 6607 3939 6613
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 4338 6644 4344 6656
rect 4299 6616 4344 6644
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 4798 6644 4804 6656
rect 4759 6616 4804 6644
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 5276 6644 5304 6740
rect 6181 6715 6239 6721
rect 6181 6681 6193 6715
rect 6227 6712 6239 6715
rect 6638 6712 6644 6724
rect 6227 6684 6644 6712
rect 6227 6681 6239 6684
rect 6181 6675 6239 6681
rect 6638 6672 6644 6684
rect 6696 6672 6702 6724
rect 6748 6712 6776 6743
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 6917 6783 6975 6789
rect 6917 6780 6929 6783
rect 6880 6752 6929 6780
rect 6880 6740 6886 6752
rect 6917 6749 6929 6752
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6749 8355 6783
rect 8478 6780 8484 6792
rect 8439 6752 8484 6780
rect 8297 6743 8355 6749
rect 7006 6712 7012 6724
rect 6748 6684 7012 6712
rect 7006 6672 7012 6684
rect 7064 6712 7070 6724
rect 7374 6712 7380 6724
rect 7064 6684 7380 6712
rect 7064 6672 7070 6684
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 7558 6672 7564 6724
rect 7616 6712 7622 6724
rect 7929 6715 7987 6721
rect 7929 6712 7941 6715
rect 7616 6684 7941 6712
rect 7616 6672 7622 6684
rect 7929 6681 7941 6684
rect 7975 6681 7987 6715
rect 7929 6675 7987 6681
rect 8202 6672 8208 6724
rect 8260 6712 8266 6724
rect 8312 6712 8340 6743
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 9490 6740 9496 6792
rect 9548 6740 9554 6792
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9732 6752 10149 6780
rect 9732 6740 9738 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6780 10379 6783
rect 10870 6780 10876 6792
rect 10367 6752 10876 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 10870 6740 10876 6752
rect 10928 6780 10934 6792
rect 11164 6780 11192 6888
rect 11238 6876 11244 6888
rect 11296 6876 11302 6928
rect 11348 6848 11376 6956
rect 13538 6944 13544 6996
rect 13596 6984 13602 6996
rect 13596 6956 14320 6984
rect 13596 6944 13602 6956
rect 12986 6916 12992 6928
rect 12544 6888 12992 6916
rect 12544 6857 12572 6888
rect 12986 6876 12992 6888
rect 13044 6876 13050 6928
rect 13814 6916 13820 6928
rect 13740 6888 13820 6916
rect 12802 6857 12808 6860
rect 11425 6851 11483 6857
rect 11425 6848 11437 6851
rect 11348 6820 11437 6848
rect 10928 6752 11192 6780
rect 10928 6740 10934 6752
rect 11238 6740 11244 6792
rect 11296 6780 11302 6792
rect 11348 6780 11376 6820
rect 11425 6817 11437 6820
rect 11471 6817 11483 6851
rect 11425 6811 11483 6817
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6817 12587 6851
rect 12796 6848 12808 6857
rect 12715 6820 12808 6848
rect 12529 6811 12587 6817
rect 12796 6811 12808 6820
rect 12860 6848 12866 6860
rect 13740 6848 13768 6888
rect 13814 6876 13820 6888
rect 13872 6876 13878 6928
rect 14292 6916 14320 6956
rect 14366 6944 14372 6996
rect 14424 6984 14430 6996
rect 14461 6987 14519 6993
rect 14461 6984 14473 6987
rect 14424 6956 14473 6984
rect 14424 6944 14430 6956
rect 14461 6953 14473 6956
rect 14507 6953 14519 6987
rect 14461 6947 14519 6953
rect 15105 6987 15163 6993
rect 15105 6953 15117 6987
rect 15151 6984 15163 6987
rect 15194 6984 15200 6996
rect 15151 6956 15200 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 15194 6944 15200 6956
rect 15252 6944 15258 6996
rect 21634 6984 21640 6996
rect 15755 6956 21640 6984
rect 14918 6916 14924 6928
rect 14292 6888 14924 6916
rect 14918 6876 14924 6888
rect 14976 6876 14982 6928
rect 15755 6916 15783 6956
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 22373 6987 22431 6993
rect 22373 6953 22385 6987
rect 22419 6984 22431 6987
rect 22554 6984 22560 6996
rect 22419 6956 22560 6984
rect 22419 6953 22431 6956
rect 22373 6947 22431 6953
rect 22554 6944 22560 6956
rect 22612 6944 22618 6996
rect 22848 6956 23152 6984
rect 15120 6888 15783 6916
rect 15933 6919 15991 6925
rect 15120 6848 15148 6888
rect 15933 6885 15945 6919
rect 15979 6885 15991 6919
rect 15933 6879 15991 6885
rect 12860 6820 13768 6848
rect 15028 6820 15148 6848
rect 12802 6808 12808 6811
rect 12860 6808 12866 6820
rect 11296 6752 11376 6780
rect 11296 6740 11302 6752
rect 9508 6712 9536 6740
rect 14090 6712 14096 6724
rect 8260 6684 9536 6712
rect 13464 6684 14096 6712
rect 8260 6672 8266 6684
rect 6365 6647 6423 6653
rect 6365 6644 6377 6647
rect 5276 6616 6377 6644
rect 6365 6613 6377 6616
rect 6411 6613 6423 6647
rect 8938 6644 8944 6656
rect 8899 6616 8944 6644
rect 6365 6607 6423 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9490 6644 9496 6656
rect 9451 6616 9496 6644
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9766 6644 9772 6656
rect 9727 6616 9772 6644
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 10686 6644 10692 6656
rect 10647 6616 10692 6644
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 11606 6644 11612 6656
rect 11567 6616 11612 6644
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 12069 6647 12127 6653
rect 12069 6613 12081 6647
rect 12115 6644 12127 6647
rect 12342 6644 12348 6656
rect 12115 6616 12348 6644
rect 12115 6613 12127 6616
rect 12069 6607 12127 6613
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 13464 6644 13492 6684
rect 14090 6672 14096 6684
rect 14148 6672 14154 6724
rect 14274 6672 14280 6724
rect 14332 6712 14338 6724
rect 14734 6712 14740 6724
rect 14332 6684 14740 6712
rect 14332 6672 14338 6684
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 12492 6616 13492 6644
rect 12492 6604 12498 6616
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 13909 6647 13967 6653
rect 13909 6644 13921 6647
rect 13872 6616 13921 6644
rect 13872 6604 13878 6616
rect 13909 6613 13921 6616
rect 13955 6644 13967 6647
rect 15028 6644 15056 6820
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 15749 6851 15807 6857
rect 15749 6848 15761 6851
rect 15436 6820 15761 6848
rect 15436 6808 15442 6820
rect 15749 6817 15761 6820
rect 15795 6817 15807 6851
rect 15749 6811 15807 6817
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 15948 6848 15976 6879
rect 16206 6876 16212 6928
rect 16264 6916 16270 6928
rect 16393 6919 16451 6925
rect 16393 6916 16405 6919
rect 16264 6888 16405 6916
rect 16264 6876 16270 6888
rect 16393 6885 16405 6888
rect 16439 6916 16451 6919
rect 16850 6916 16856 6928
rect 16439 6888 16856 6916
rect 16439 6885 16451 6888
rect 16393 6879 16451 6885
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 17144 6888 17724 6916
rect 16945 6851 17003 6857
rect 15896 6820 16160 6848
rect 15896 6808 15902 6820
rect 15194 6740 15200 6792
rect 15252 6780 15258 6792
rect 15856 6780 15884 6808
rect 16022 6780 16028 6792
rect 15252 6752 15884 6780
rect 15983 6752 16028 6780
rect 15252 6740 15258 6752
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16132 6780 16160 6820
rect 16945 6817 16957 6851
rect 16991 6848 17003 6851
rect 17144 6848 17172 6888
rect 16991 6820 17172 6848
rect 17212 6851 17270 6857
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17212 6817 17224 6851
rect 17258 6848 17270 6851
rect 17586 6848 17592 6860
rect 17258 6820 17592 6848
rect 17258 6817 17270 6820
rect 17212 6811 17270 6817
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 17696 6848 17724 6888
rect 19794 6876 19800 6928
rect 19852 6916 19858 6928
rect 20346 6916 20352 6928
rect 19852 6888 20352 6916
rect 19852 6876 19858 6888
rect 20346 6876 20352 6888
rect 20404 6876 20410 6928
rect 21453 6919 21511 6925
rect 21453 6916 21465 6919
rect 20456 6888 21465 6916
rect 20456 6860 20484 6888
rect 21453 6885 21465 6888
rect 21499 6885 21511 6919
rect 21453 6879 21511 6885
rect 22002 6876 22008 6928
rect 22060 6916 22066 6928
rect 22646 6916 22652 6928
rect 22060 6888 22652 6916
rect 22060 6876 22066 6888
rect 22646 6876 22652 6888
rect 22704 6916 22710 6928
rect 22848 6916 22876 6956
rect 23014 6916 23020 6928
rect 22704 6888 22876 6916
rect 22975 6888 23020 6916
rect 22704 6876 22710 6888
rect 23014 6876 23020 6888
rect 23072 6876 23078 6928
rect 23124 6925 23152 6956
rect 23109 6919 23167 6925
rect 23109 6885 23121 6919
rect 23155 6916 23167 6919
rect 24578 6916 24584 6928
rect 23155 6888 23612 6916
rect 24491 6888 24584 6916
rect 23155 6885 23167 6888
rect 23109 6879 23167 6885
rect 17770 6848 17776 6860
rect 17696 6820 17776 6848
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 19058 6808 19064 6860
rect 19116 6848 19122 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 19116 6820 19257 6848
rect 19116 6808 19122 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 19518 6808 19524 6860
rect 19576 6848 19582 6860
rect 19705 6851 19763 6857
rect 19705 6848 19717 6851
rect 19576 6820 19717 6848
rect 19576 6808 19582 6820
rect 19705 6817 19717 6820
rect 19751 6848 19763 6851
rect 20438 6848 20444 6860
rect 19751 6820 20444 6848
rect 19751 6817 19763 6820
rect 19705 6811 19763 6817
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 20806 6808 20812 6860
rect 20864 6848 20870 6860
rect 21726 6848 21732 6860
rect 20864 6820 21732 6848
rect 20864 6808 20870 6820
rect 21726 6808 21732 6820
rect 21784 6848 21790 6860
rect 21913 6851 21971 6857
rect 21913 6848 21925 6851
rect 21784 6820 21925 6848
rect 21784 6808 21790 6820
rect 21913 6817 21925 6820
rect 21959 6817 21971 6851
rect 23474 6848 23480 6860
rect 23435 6820 23480 6848
rect 21913 6811 21971 6817
rect 16482 6780 16488 6792
rect 16132 6752 16488 6780
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 19426 6740 19432 6792
rect 19484 6780 19490 6792
rect 19613 6783 19671 6789
rect 19613 6780 19625 6783
rect 19484 6752 19625 6780
rect 19484 6740 19490 6752
rect 19613 6749 19625 6752
rect 19659 6780 19671 6783
rect 20530 6780 20536 6792
rect 19659 6752 20536 6780
rect 19659 6749 19671 6752
rect 19613 6743 19671 6749
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 20622 6740 20628 6792
rect 20680 6780 20686 6792
rect 21450 6780 21456 6792
rect 20680 6752 21456 6780
rect 20680 6740 20686 6752
rect 21450 6740 21456 6752
rect 21508 6740 21514 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6749 21603 6783
rect 21928 6780 21956 6811
rect 23474 6808 23480 6820
rect 23532 6808 23538 6860
rect 23584 6848 23612 6888
rect 24578 6876 24584 6888
rect 24636 6916 24642 6928
rect 25682 6916 25688 6928
rect 24636 6888 25688 6916
rect 24636 6876 24642 6888
rect 25682 6876 25688 6888
rect 25740 6876 25746 6928
rect 23845 6851 23903 6857
rect 23845 6848 23857 6851
rect 23584 6820 23857 6848
rect 23845 6817 23857 6820
rect 23891 6848 23903 6851
rect 24210 6848 24216 6860
rect 23891 6820 24216 6848
rect 23891 6817 23903 6820
rect 23845 6811 23903 6817
rect 24210 6808 24216 6820
rect 24268 6848 24274 6860
rect 24673 6851 24731 6857
rect 24673 6848 24685 6851
rect 24268 6820 24685 6848
rect 24268 6808 24274 6820
rect 24673 6817 24685 6820
rect 24719 6817 24731 6851
rect 25406 6848 25412 6860
rect 25367 6820 25412 6848
rect 24673 6811 24731 6817
rect 25406 6808 25412 6820
rect 25464 6808 25470 6860
rect 26237 6851 26295 6857
rect 26237 6817 26249 6851
rect 26283 6848 26295 6851
rect 26418 6848 26424 6860
rect 26283 6820 26424 6848
rect 26283 6817 26295 6820
rect 26237 6811 26295 6817
rect 26418 6808 26424 6820
rect 26476 6808 26482 6860
rect 23017 6783 23075 6789
rect 21928 6752 22692 6780
rect 21545 6743 21603 6749
rect 19889 6715 19947 6721
rect 19889 6681 19901 6715
rect 19935 6712 19947 6715
rect 20346 6712 20352 6724
rect 19935 6684 20352 6712
rect 19935 6681 19947 6684
rect 19889 6675 19947 6681
rect 20346 6672 20352 6684
rect 20404 6672 20410 6724
rect 20990 6712 20996 6724
rect 20951 6684 20996 6712
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 15470 6644 15476 6656
rect 13955 6616 15056 6644
rect 15431 6616 15476 6644
rect 13955 6613 13967 6616
rect 13909 6607 13967 6613
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 16942 6644 16948 6656
rect 16899 6616 16948 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 18325 6647 18383 6653
rect 18325 6644 18337 6647
rect 17920 6616 18337 6644
rect 17920 6604 17926 6616
rect 18325 6613 18337 6616
rect 18371 6644 18383 6647
rect 18690 6644 18696 6656
rect 18371 6616 18696 6644
rect 18371 6613 18383 6616
rect 18325 6607 18383 6613
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 20254 6644 20260 6656
rect 20215 6616 20260 6644
rect 20254 6604 20260 6616
rect 20312 6644 20318 6656
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 20312 6616 20637 6644
rect 20312 6604 20318 6616
rect 20625 6613 20637 6616
rect 20671 6644 20683 6647
rect 21560 6644 21588 6743
rect 21910 6672 21916 6724
rect 21968 6712 21974 6724
rect 22557 6715 22615 6721
rect 22557 6712 22569 6715
rect 21968 6684 22569 6712
rect 21968 6672 21974 6684
rect 22557 6681 22569 6684
rect 22603 6681 22615 6715
rect 22557 6675 22615 6681
rect 21818 6644 21824 6656
rect 20671 6616 21824 6644
rect 20671 6613 20683 6616
rect 20625 6607 20683 6613
rect 21818 6604 21824 6616
rect 21876 6604 21882 6656
rect 22664 6644 22692 6752
rect 23017 6749 23029 6783
rect 23063 6780 23075 6783
rect 23198 6780 23204 6792
rect 23063 6752 23204 6780
rect 23063 6749 23075 6752
rect 23017 6743 23075 6749
rect 23198 6740 23204 6752
rect 23256 6740 23262 6792
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 25038 6780 25044 6792
rect 24627 6752 25044 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 24026 6672 24032 6724
rect 24084 6712 24090 6724
rect 24121 6715 24179 6721
rect 24121 6712 24133 6715
rect 24084 6684 24133 6712
rect 24084 6672 24090 6684
rect 24121 6681 24133 6684
rect 24167 6681 24179 6715
rect 24121 6675 24179 6681
rect 24596 6644 24624 6743
rect 25038 6740 25044 6752
rect 25096 6740 25102 6792
rect 25774 6780 25780 6792
rect 25735 6752 25780 6780
rect 25774 6740 25780 6752
rect 25832 6740 25838 6792
rect 22664 6616 24624 6644
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25041 6647 25099 6653
rect 25041 6644 25053 6647
rect 24912 6616 25053 6644
rect 24912 6604 24918 6616
rect 25041 6613 25053 6616
rect 25087 6613 25099 6647
rect 25041 6607 25099 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 5442 6440 5448 6452
rect 4479 6412 5448 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 5442 6400 5448 6412
rect 5500 6440 5506 6452
rect 6086 6440 6092 6452
rect 5500 6412 6092 6440
rect 5500 6400 5506 6412
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6914 6440 6920 6452
rect 6875 6412 6920 6440
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 7926 6440 7932 6452
rect 7887 6412 7932 6440
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8573 6443 8631 6449
rect 8573 6440 8585 6443
rect 8168 6412 8585 6440
rect 8168 6400 8174 6412
rect 8573 6409 8585 6412
rect 8619 6409 8631 6443
rect 8573 6403 8631 6409
rect 4982 6372 4988 6384
rect 4908 6344 4988 6372
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6304 1823 6307
rect 1854 6304 1860 6316
rect 1811 6276 1860 6304
rect 1811 6273 1823 6276
rect 1765 6267 1823 6273
rect 1854 6264 1860 6276
rect 1912 6264 1918 6316
rect 4908 6313 4936 6344
rect 4982 6332 4988 6344
rect 5040 6332 5046 6384
rect 5997 6375 6055 6381
rect 5997 6341 6009 6375
rect 6043 6372 6055 6375
rect 7006 6372 7012 6384
rect 6043 6344 7012 6372
rect 6043 6341 6055 6344
rect 5997 6335 6055 6341
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6304 7435 6307
rect 7466 6304 7472 6316
rect 7423 6276 7472 6304
rect 7423 6273 7435 6276
rect 7377 6267 7435 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 8588 6304 8616 6403
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 9456 6412 10149 6440
rect 9456 6400 9462 6412
rect 10137 6409 10149 6412
rect 10183 6409 10195 6443
rect 10137 6403 10195 6409
rect 10781 6443 10839 6449
rect 10781 6409 10793 6443
rect 10827 6440 10839 6443
rect 10870 6440 10876 6452
rect 10827 6412 10876 6440
rect 10827 6409 10839 6412
rect 10781 6403 10839 6409
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11296 6412 11805 6440
rect 11296 6400 11302 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12802 6440 12808 6452
rect 12299 6412 12808 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 12986 6440 12992 6452
rect 12947 6412 12992 6440
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 14366 6400 14372 6452
rect 14424 6400 14430 6452
rect 14734 6400 14740 6452
rect 14792 6440 14798 6452
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 14792 6412 14841 6440
rect 14792 6400 14798 6412
rect 14829 6409 14841 6412
rect 14875 6440 14887 6443
rect 15746 6440 15752 6452
rect 14875 6412 15752 6440
rect 14875 6409 14887 6412
rect 14829 6403 14887 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 15838 6400 15844 6452
rect 15896 6440 15902 6452
rect 15896 6412 15941 6440
rect 15896 6400 15902 6412
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 18506 6440 18512 6452
rect 17000 6412 18512 6440
rect 17000 6400 17006 6412
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 19518 6440 19524 6452
rect 19479 6412 19524 6440
rect 19518 6400 19524 6412
rect 19576 6400 19582 6452
rect 20438 6400 20444 6452
rect 20496 6440 20502 6452
rect 20901 6443 20959 6449
rect 20901 6440 20913 6443
rect 20496 6412 20913 6440
rect 20496 6400 20502 6412
rect 20901 6409 20913 6412
rect 20947 6440 20959 6443
rect 21082 6440 21088 6452
rect 20947 6412 21088 6440
rect 20947 6409 20959 6412
rect 20901 6403 20959 6409
rect 21082 6400 21088 6412
rect 21140 6400 21146 6452
rect 22554 6400 22560 6452
rect 22612 6440 22618 6452
rect 25406 6440 25412 6452
rect 22612 6412 25412 6440
rect 22612 6400 22618 6412
rect 25406 6400 25412 6412
rect 25464 6400 25470 6452
rect 14384 6372 14412 6400
rect 16209 6375 16267 6381
rect 16209 6372 16221 6375
rect 14384 6344 16221 6372
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 8588 6276 8769 6304
rect 8757 6273 8769 6276
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 2124 6239 2182 6245
rect 2124 6205 2136 6239
rect 2170 6236 2182 6239
rect 2498 6236 2504 6248
rect 2170 6208 2504 6236
rect 2170 6205 2182 6208
rect 2124 6199 2182 6205
rect 2498 6196 2504 6208
rect 2556 6236 2562 6248
rect 3050 6236 3056 6248
rect 2556 6208 3056 6236
rect 2556 6196 2562 6208
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3418 6236 3424 6248
rect 3292 6208 3424 6236
rect 3292 6196 3298 6208
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4614 6236 4620 6248
rect 4295 6208 4620 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4614 6196 4620 6208
rect 4672 6236 4678 6248
rect 4985 6239 5043 6245
rect 4985 6236 4997 6239
rect 4672 6208 4997 6236
rect 4672 6196 4678 6208
rect 4985 6205 4997 6208
rect 5031 6205 5043 6239
rect 8772 6236 8800 6267
rect 10594 6264 10600 6316
rect 10652 6304 10658 6316
rect 10870 6304 10876 6316
rect 10652 6276 10876 6304
rect 10652 6264 10658 6276
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 11054 6264 11060 6316
rect 11112 6304 11118 6316
rect 11149 6307 11207 6313
rect 11149 6304 11161 6307
rect 11112 6276 11161 6304
rect 11112 6264 11118 6276
rect 11149 6273 11161 6276
rect 11195 6304 11207 6307
rect 12250 6304 12256 6316
rect 11195 6276 12256 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11256 6245 11284 6276
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 11241 6239 11299 6245
rect 8772 6208 9168 6236
rect 4985 6199 5043 6205
rect 4893 6171 4951 6177
rect 4893 6137 4905 6171
rect 4939 6168 4951 6171
rect 5166 6168 5172 6180
rect 4939 6140 5172 6168
rect 4939 6137 4951 6140
rect 4893 6131 4951 6137
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 6822 6128 6828 6180
rect 6880 6168 6886 6180
rect 7466 6168 7472 6180
rect 6880 6140 7472 6168
rect 6880 6128 6886 6140
rect 7466 6128 7472 6140
rect 7524 6128 7530 6180
rect 9002 6171 9060 6177
rect 9002 6168 9014 6171
rect 8312 6140 9014 6168
rect 8312 6112 8340 6140
rect 9002 6137 9014 6140
rect 9048 6137 9060 6171
rect 9140 6168 9168 6208
rect 11241 6205 11253 6239
rect 11287 6236 11299 6239
rect 13449 6239 13507 6245
rect 11287 6208 11321 6236
rect 11287 6205 11299 6208
rect 11241 6199 11299 6205
rect 13449 6205 13461 6239
rect 13495 6205 13507 6239
rect 13449 6199 13507 6205
rect 12986 6168 12992 6180
rect 9140 6140 12992 6168
rect 9002 6131 9060 6137
rect 12986 6128 12992 6140
rect 13044 6168 13050 6180
rect 13265 6171 13323 6177
rect 13265 6168 13277 6171
rect 13044 6140 13277 6168
rect 13044 6128 13050 6140
rect 13265 6137 13277 6140
rect 13311 6168 13323 6171
rect 13464 6168 13492 6199
rect 13538 6168 13544 6180
rect 13311 6140 13544 6168
rect 13311 6137 13323 6140
rect 13265 6131 13323 6137
rect 13538 6128 13544 6140
rect 13596 6128 13602 6180
rect 13716 6171 13774 6177
rect 13716 6137 13728 6171
rect 13762 6168 13774 6171
rect 13814 6168 13820 6180
rect 13762 6140 13820 6168
rect 13762 6137 13774 6140
rect 13716 6131 13774 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 15948 6168 15976 6344
rect 16209 6341 16221 6344
rect 16255 6341 16267 6375
rect 16209 6335 16267 6341
rect 16485 6375 16543 6381
rect 16485 6341 16497 6375
rect 16531 6372 16543 6375
rect 17034 6372 17040 6384
rect 16531 6344 17040 6372
rect 16531 6341 16543 6344
rect 16485 6335 16543 6341
rect 17034 6332 17040 6344
rect 17092 6332 17098 6384
rect 18138 6372 18144 6384
rect 18099 6344 18144 6372
rect 18138 6332 18144 6344
rect 18196 6332 18202 6384
rect 19702 6372 19708 6384
rect 18616 6344 19708 6372
rect 16850 6304 16856 6316
rect 16811 6276 16856 6304
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 18616 6313 18644 6344
rect 19702 6332 19708 6344
rect 19760 6332 19766 6384
rect 21266 6372 21272 6384
rect 21227 6344 21272 6372
rect 21266 6332 21272 6344
rect 21324 6332 21330 6384
rect 22002 6332 22008 6384
rect 22060 6372 22066 6384
rect 23382 6372 23388 6384
rect 22060 6344 23388 6372
rect 22060 6332 22066 6344
rect 23382 6332 23388 6344
rect 23440 6372 23446 6384
rect 23845 6375 23903 6381
rect 23845 6372 23857 6375
rect 23440 6344 23857 6372
rect 23440 6332 23446 6344
rect 23845 6341 23857 6344
rect 23891 6341 23903 6375
rect 23845 6335 23903 6341
rect 18601 6307 18659 6313
rect 18601 6273 18613 6307
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 18690 6264 18696 6316
rect 18748 6304 18754 6316
rect 19153 6307 19211 6313
rect 19153 6304 19165 6307
rect 18748 6276 19165 6304
rect 18748 6264 18754 6276
rect 19153 6273 19165 6276
rect 19199 6304 19211 6307
rect 20257 6307 20315 6313
rect 20257 6304 20269 6307
rect 19199 6276 20269 6304
rect 19199 6273 19211 6276
rect 19153 6267 19211 6273
rect 20257 6273 20269 6276
rect 20303 6273 20315 6307
rect 20257 6267 20315 6273
rect 16022 6196 16028 6248
rect 16080 6236 16086 6248
rect 17037 6239 17095 6245
rect 17037 6236 17049 6239
rect 16080 6208 17049 6236
rect 16080 6196 16086 6208
rect 17037 6205 17049 6208
rect 17083 6236 17095 6239
rect 17586 6236 17592 6248
rect 17083 6208 17592 6236
rect 17083 6205 17095 6208
rect 17037 6199 17095 6205
rect 17586 6196 17592 6208
rect 17644 6236 17650 6248
rect 17773 6239 17831 6245
rect 17773 6236 17785 6239
rect 17644 6208 17785 6236
rect 17644 6196 17650 6208
rect 17773 6205 17785 6208
rect 17819 6205 17831 6239
rect 19978 6236 19984 6248
rect 19939 6208 19984 6236
rect 17773 6199 17831 6205
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 21284 6236 21312 6332
rect 21818 6304 21824 6316
rect 21779 6276 21824 6304
rect 21818 6264 21824 6276
rect 21876 6264 21882 6316
rect 23860 6304 23888 6335
rect 24029 6307 24087 6313
rect 24029 6304 24041 6307
rect 23860 6276 24041 6304
rect 24029 6273 24041 6276
rect 24075 6273 24087 6307
rect 25958 6304 25964 6316
rect 25919 6276 25964 6304
rect 24029 6267 24087 6273
rect 25958 6264 25964 6276
rect 26016 6264 26022 6316
rect 20180 6208 21312 6236
rect 21545 6239 21603 6245
rect 16945 6171 17003 6177
rect 16945 6168 16957 6171
rect 15948 6140 16957 6168
rect 16945 6137 16957 6140
rect 16991 6137 17003 6171
rect 18690 6168 18696 6180
rect 18651 6140 18696 6168
rect 16945 6131 17003 6137
rect 18690 6128 18696 6140
rect 18748 6128 18754 6180
rect 20180 6177 20208 6208
rect 21545 6205 21557 6239
rect 21591 6236 21603 6239
rect 22094 6236 22100 6248
rect 21591 6208 22100 6236
rect 21591 6205 21603 6208
rect 21545 6199 21603 6205
rect 20165 6171 20223 6177
rect 20165 6137 20177 6171
rect 20211 6137 20223 6171
rect 20165 6131 20223 6137
rect 20806 6128 20812 6180
rect 20864 6168 20870 6180
rect 21560 6168 21588 6199
rect 22094 6196 22100 6208
rect 22152 6236 22158 6248
rect 26602 6236 26608 6248
rect 22152 6208 26608 6236
rect 22152 6196 22158 6208
rect 26602 6196 26608 6208
rect 26660 6196 26666 6248
rect 21726 6168 21732 6180
rect 20864 6140 21588 6168
rect 21687 6140 21732 6168
rect 20864 6128 20870 6140
rect 21726 6128 21732 6140
rect 21784 6128 21790 6180
rect 22557 6171 22615 6177
rect 22557 6137 22569 6171
rect 22603 6168 22615 6171
rect 23014 6168 23020 6180
rect 22603 6140 23020 6168
rect 22603 6137 22615 6140
rect 22557 6131 22615 6137
rect 23014 6128 23020 6140
rect 23072 6128 23078 6180
rect 24210 6128 24216 6180
rect 24268 6177 24274 6180
rect 24268 6171 24332 6177
rect 24268 6137 24286 6171
rect 24320 6137 24332 6171
rect 24268 6131 24332 6137
rect 24268 6128 24274 6131
rect 24486 6128 24492 6180
rect 24544 6168 24550 6180
rect 25866 6168 25872 6180
rect 24544 6140 25872 6168
rect 24544 6128 24550 6140
rect 25866 6128 25872 6140
rect 25924 6128 25930 6180
rect 3234 6100 3240 6112
rect 3195 6072 3240 6100
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 3881 6103 3939 6109
rect 3881 6069 3893 6103
rect 3927 6100 3939 6103
rect 5074 6100 5080 6112
rect 3927 6072 5080 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5445 6103 5503 6109
rect 5445 6069 5457 6103
rect 5491 6100 5503 6103
rect 5534 6100 5540 6112
rect 5491 6072 5540 6100
rect 5491 6069 5503 6072
rect 5445 6063 5503 6069
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 5902 6060 5908 6112
rect 5960 6100 5966 6112
rect 6273 6103 6331 6109
rect 6273 6100 6285 6103
rect 5960 6072 6285 6100
rect 5960 6060 5966 6072
rect 6273 6069 6285 6072
rect 6319 6100 6331 6103
rect 6362 6100 6368 6112
rect 6319 6072 6368 6100
rect 6319 6069 6331 6072
rect 6273 6063 6331 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 7377 6103 7435 6109
rect 7377 6069 7389 6103
rect 7423 6100 7435 6103
rect 7926 6100 7932 6112
rect 7423 6072 7932 6100
rect 7423 6069 7435 6072
rect 7377 6063 7435 6069
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8294 6100 8300 6112
rect 8255 6072 8300 6100
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 11425 6103 11483 6109
rect 11425 6069 11437 6103
rect 11471 6100 11483 6103
rect 11514 6100 11520 6112
rect 11471 6072 11520 6100
rect 11471 6069 11483 6072
rect 11425 6063 11483 6069
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12492 6072 12537 6100
rect 12492 6060 12498 6072
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 15378 6100 15384 6112
rect 12860 6072 15384 6100
rect 12860 6060 12866 6072
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 17497 6103 17555 6109
rect 17497 6069 17509 6103
rect 17543 6100 17555 6103
rect 17770 6100 17776 6112
rect 17543 6072 17776 6100
rect 17543 6069 17555 6072
rect 17497 6063 17555 6069
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 18598 6100 18604 6112
rect 18559 6072 18604 6100
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 22925 6103 22983 6109
rect 22925 6069 22937 6103
rect 22971 6100 22983 6103
rect 23198 6100 23204 6112
rect 22971 6072 23204 6100
rect 22971 6069 22983 6072
rect 22925 6063 22983 6069
rect 23198 6060 23204 6072
rect 23256 6060 23262 6112
rect 23477 6103 23535 6109
rect 23477 6069 23489 6103
rect 23523 6100 23535 6103
rect 25682 6100 25688 6112
rect 23523 6072 25688 6100
rect 23523 6069 23535 6072
rect 23477 6063 23535 6069
rect 25682 6060 25688 6072
rect 25740 6060 25746 6112
rect 26326 6100 26332 6112
rect 26287 6072 26332 6100
rect 26326 6060 26332 6072
rect 26384 6060 26390 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2498 5896 2504 5908
rect 2056 5868 2504 5896
rect 1762 5828 1768 5840
rect 1723 5800 1768 5828
rect 1762 5788 1768 5800
rect 1820 5788 1826 5840
rect 2056 5837 2084 5868
rect 2498 5856 2504 5868
rect 2556 5896 2562 5908
rect 2777 5899 2835 5905
rect 2777 5896 2789 5899
rect 2556 5868 2789 5896
rect 2556 5856 2562 5868
rect 2777 5865 2789 5868
rect 2823 5865 2835 5899
rect 2777 5859 2835 5865
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 7098 5896 7104 5908
rect 3384 5868 7104 5896
rect 3384 5856 3390 5868
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8536 5868 8861 5896
rect 8536 5856 8542 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 10229 5899 10287 5905
rect 10229 5896 10241 5899
rect 9548 5868 10241 5896
rect 9548 5856 9554 5868
rect 10229 5865 10241 5868
rect 10275 5896 10287 5899
rect 11315 5899 11373 5905
rect 11315 5896 11327 5899
rect 10275 5868 11327 5896
rect 10275 5865 10287 5868
rect 10229 5859 10287 5865
rect 11315 5865 11327 5868
rect 11361 5865 11373 5899
rect 11315 5859 11373 5865
rect 12529 5899 12587 5905
rect 12529 5865 12541 5899
rect 12575 5896 12587 5899
rect 12618 5896 12624 5908
rect 12575 5868 12624 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 13814 5896 13820 5908
rect 13587 5868 13820 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 14734 5896 14740 5908
rect 13924 5868 14320 5896
rect 14695 5868 14740 5896
rect 2041 5831 2099 5837
rect 2041 5797 2053 5831
rect 2087 5797 2099 5831
rect 2041 5791 2099 5797
rect 4614 5788 4620 5840
rect 4672 5837 4678 5840
rect 4672 5831 4736 5837
rect 4672 5797 4690 5831
rect 4724 5797 4736 5831
rect 6914 5828 6920 5840
rect 4672 5791 4736 5797
rect 6012 5800 6920 5828
rect 4672 5788 4678 5791
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 6012 5760 6040 5800
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 8110 5828 8116 5840
rect 7024 5800 8116 5828
rect 6822 5760 6828 5772
rect 2832 5732 6040 5760
rect 6748 5732 6828 5760
rect 2832 5720 2838 5732
rect 2958 5692 2964 5704
rect 2919 5664 2964 5692
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5661 4491 5695
rect 4433 5655 4491 5661
rect 1489 5627 1547 5633
rect 1489 5593 1501 5627
rect 1535 5624 1547 5627
rect 1946 5624 1952 5636
rect 1535 5596 1952 5624
rect 1535 5593 1547 5596
rect 1489 5587 1547 5593
rect 1946 5584 1952 5596
rect 2004 5624 2010 5636
rect 2590 5624 2596 5636
rect 2004 5596 2596 5624
rect 2004 5584 2010 5596
rect 2590 5584 2596 5596
rect 2648 5584 2654 5636
rect 3234 5516 3240 5568
rect 3292 5556 3298 5568
rect 3513 5559 3571 5565
rect 3513 5556 3525 5559
rect 3292 5528 3525 5556
rect 3292 5516 3298 5528
rect 3513 5525 3525 5528
rect 3559 5556 3571 5559
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 3559 5528 3893 5556
rect 3559 5525 3571 5528
rect 3513 5519 3571 5525
rect 3881 5525 3893 5528
rect 3927 5556 3939 5559
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 3927 5528 4261 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 4249 5525 4261 5528
rect 4295 5525 4307 5559
rect 4448 5556 4476 5655
rect 4798 5556 4804 5568
rect 4448 5528 4804 5556
rect 4249 5519 4307 5525
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 6270 5556 6276 5568
rect 5859 5528 6276 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 6270 5516 6276 5528
rect 6328 5556 6334 5568
rect 6748 5565 6776 5732
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 6914 5692 6920 5704
rect 6827 5664 6920 5692
rect 6914 5652 6920 5664
rect 6972 5692 6978 5704
rect 7024 5692 7052 5800
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 10045 5831 10103 5837
rect 10045 5828 10057 5831
rect 9824 5800 10057 5828
rect 9824 5788 9830 5800
rect 10045 5797 10057 5800
rect 10091 5828 10103 5831
rect 10686 5828 10692 5840
rect 10091 5800 10692 5828
rect 10091 5797 10103 5800
rect 10045 5791 10103 5797
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 10778 5788 10784 5840
rect 10836 5828 10842 5840
rect 10836 5800 10881 5828
rect 10836 5788 10842 5800
rect 11422 5788 11428 5840
rect 11480 5828 11486 5840
rect 11609 5831 11667 5837
rect 11609 5828 11621 5831
rect 11480 5800 11621 5828
rect 11480 5788 11486 5800
rect 11609 5797 11621 5800
rect 11655 5797 11667 5831
rect 11790 5828 11796 5840
rect 11751 5800 11796 5828
rect 11609 5791 11667 5797
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 7184 5763 7242 5769
rect 7184 5729 7196 5763
rect 7230 5760 7242 5763
rect 7466 5760 7472 5772
rect 7230 5732 7472 5760
rect 7230 5729 7242 5732
rect 7184 5723 7242 5729
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10796 5760 10824 5788
rect 10367 5732 10824 5760
rect 11164 5732 13768 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 6972 5664 7052 5692
rect 6972 5652 6978 5664
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 11164 5692 11192 5732
rect 9364 5664 11192 5692
rect 9364 5652 9370 5664
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 11885 5695 11943 5701
rect 11885 5692 11897 5695
rect 11296 5664 11897 5692
rect 11296 5652 11302 5664
rect 11885 5661 11897 5664
rect 11931 5661 11943 5695
rect 13740 5692 13768 5732
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 13924 5760 13952 5868
rect 14292 5837 14320 5868
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 16022 5896 16028 5908
rect 15151 5868 16028 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 16022 5856 16028 5868
rect 16080 5856 16086 5908
rect 16298 5896 16304 5908
rect 16259 5868 16304 5896
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 17586 5896 17592 5908
rect 17547 5868 17592 5896
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 17957 5899 18015 5905
rect 17957 5865 17969 5899
rect 18003 5896 18015 5899
rect 18690 5896 18696 5908
rect 18003 5868 18696 5896
rect 18003 5865 18015 5868
rect 17957 5859 18015 5865
rect 18690 5856 18696 5868
rect 18748 5896 18754 5908
rect 19061 5899 19119 5905
rect 19061 5896 19073 5899
rect 18748 5868 19073 5896
rect 18748 5856 18754 5868
rect 19061 5865 19073 5868
rect 19107 5865 19119 5899
rect 19061 5859 19119 5865
rect 19889 5899 19947 5905
rect 19889 5865 19901 5899
rect 19935 5896 19947 5899
rect 20438 5896 20444 5908
rect 19935 5868 20444 5896
rect 19935 5865 19947 5868
rect 19889 5859 19947 5865
rect 20438 5856 20444 5868
rect 20496 5856 20502 5908
rect 20717 5899 20775 5905
rect 20717 5865 20729 5899
rect 20763 5896 20775 5899
rect 20806 5896 20812 5908
rect 20763 5868 20812 5896
rect 20763 5865 20775 5868
rect 20717 5859 20775 5865
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 21177 5899 21235 5905
rect 21177 5865 21189 5899
rect 21223 5896 21235 5899
rect 21634 5896 21640 5908
rect 21223 5868 21640 5896
rect 21223 5865 21235 5868
rect 21177 5859 21235 5865
rect 21634 5856 21640 5868
rect 21692 5856 21698 5908
rect 22646 5896 22652 5908
rect 22607 5868 22652 5896
rect 22646 5856 22652 5868
rect 22704 5896 22710 5908
rect 23201 5899 23259 5905
rect 23201 5896 23213 5899
rect 22704 5868 23213 5896
rect 22704 5856 22710 5868
rect 23201 5865 23213 5868
rect 23247 5896 23259 5899
rect 23569 5899 23627 5905
rect 23569 5896 23581 5899
rect 23247 5868 23581 5896
rect 23247 5865 23259 5868
rect 23201 5859 23259 5865
rect 23569 5865 23581 5868
rect 23615 5865 23627 5899
rect 23569 5859 23627 5865
rect 24305 5899 24363 5905
rect 24305 5865 24317 5899
rect 24351 5896 24363 5899
rect 25130 5896 25136 5908
rect 24351 5868 25136 5896
rect 24351 5865 24363 5868
rect 24305 5859 24363 5865
rect 14185 5831 14243 5837
rect 14185 5797 14197 5831
rect 14231 5797 14243 5831
rect 14185 5791 14243 5797
rect 14277 5831 14335 5837
rect 14277 5797 14289 5831
rect 14323 5828 14335 5831
rect 14550 5828 14556 5840
rect 14323 5800 14556 5828
rect 14323 5797 14335 5800
rect 14277 5791 14335 5797
rect 13872 5732 13952 5760
rect 14200 5760 14228 5791
rect 14550 5788 14556 5800
rect 14608 5788 14614 5840
rect 17034 5828 17040 5840
rect 16995 5800 17040 5828
rect 17034 5788 17040 5800
rect 17092 5788 17098 5840
rect 17129 5831 17187 5837
rect 17129 5797 17141 5831
rect 17175 5828 17187 5831
rect 17402 5828 17408 5840
rect 17175 5800 17408 5828
rect 17175 5797 17187 5800
rect 17129 5791 17187 5797
rect 17402 5788 17408 5800
rect 17460 5828 17466 5840
rect 17862 5828 17868 5840
rect 17460 5800 17868 5828
rect 17460 5788 17466 5800
rect 17862 5788 17868 5800
rect 17920 5788 17926 5840
rect 18138 5788 18144 5840
rect 18196 5828 18202 5840
rect 18601 5831 18659 5837
rect 18601 5828 18613 5831
rect 18196 5800 18613 5828
rect 18196 5788 18202 5800
rect 18601 5797 18613 5800
rect 18647 5828 18659 5831
rect 18966 5828 18972 5840
rect 18647 5800 18972 5828
rect 18647 5797 18659 5800
rect 18601 5791 18659 5797
rect 18966 5788 18972 5800
rect 19024 5788 19030 5840
rect 22738 5788 22744 5840
rect 22796 5828 22802 5840
rect 23382 5828 23388 5840
rect 22796 5800 23388 5828
rect 22796 5788 22802 5800
rect 23382 5788 23388 5800
rect 23440 5828 23446 5840
rect 24320 5828 24348 5859
rect 25130 5856 25136 5868
rect 25188 5856 25194 5908
rect 25866 5896 25872 5908
rect 25827 5868 25872 5896
rect 25866 5856 25872 5868
rect 25924 5856 25930 5908
rect 23440 5800 24348 5828
rect 23440 5788 23446 5800
rect 14366 5760 14372 5772
rect 14200 5732 14372 5760
rect 13872 5720 13878 5732
rect 14366 5720 14372 5732
rect 14424 5760 14430 5772
rect 15381 5763 15439 5769
rect 15381 5760 15393 5763
rect 14424 5732 15393 5760
rect 14424 5720 14430 5732
rect 15381 5729 15393 5732
rect 15427 5760 15439 5763
rect 15654 5760 15660 5772
rect 15427 5732 15660 5760
rect 15427 5729 15439 5732
rect 15381 5723 15439 5729
rect 15654 5720 15660 5732
rect 15712 5760 15718 5772
rect 15933 5763 15991 5769
rect 15933 5760 15945 5763
rect 15712 5732 15945 5760
rect 15712 5720 15718 5732
rect 15933 5729 15945 5732
rect 15979 5729 15991 5763
rect 15933 5723 15991 5729
rect 16758 5720 16764 5772
rect 16816 5760 16822 5772
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 16816 5732 16865 5760
rect 16816 5720 16822 5732
rect 16853 5729 16865 5732
rect 16899 5729 16911 5763
rect 16853 5723 16911 5729
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18012 5732 18736 5760
rect 18012 5720 18018 5732
rect 13740 5664 13860 5692
rect 11885 5655 11943 5661
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 9769 5627 9827 5633
rect 9769 5624 9781 5627
rect 9732 5596 9781 5624
rect 9732 5584 9738 5596
rect 9769 5593 9781 5596
rect 9815 5593 9827 5627
rect 9769 5587 9827 5593
rect 13170 5584 13176 5636
rect 13228 5624 13234 5636
rect 13725 5627 13783 5633
rect 13725 5624 13737 5627
rect 13228 5596 13737 5624
rect 13228 5584 13234 5596
rect 13725 5593 13737 5596
rect 13771 5593 13783 5627
rect 13725 5587 13783 5593
rect 6365 5559 6423 5565
rect 6365 5556 6377 5559
rect 6328 5528 6377 5556
rect 6328 5516 6334 5528
rect 6365 5525 6377 5528
rect 6411 5556 6423 5559
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6411 5528 6745 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 8110 5516 8116 5568
rect 8168 5556 8174 5568
rect 8297 5559 8355 5565
rect 8297 5556 8309 5559
rect 8168 5528 8309 5556
rect 8168 5516 8174 5528
rect 8297 5525 8309 5528
rect 8343 5525 8355 5559
rect 9306 5556 9312 5568
rect 9267 5528 9312 5556
rect 8297 5519 8355 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 11054 5556 11060 5568
rect 11015 5528 11060 5556
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 12897 5559 12955 5565
rect 12897 5525 12909 5559
rect 12943 5556 12955 5559
rect 13078 5556 13084 5568
rect 12943 5528 13084 5556
rect 12943 5525 12955 5528
rect 12897 5519 12955 5525
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 13832 5556 13860 5664
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14185 5695 14243 5701
rect 14185 5692 14197 5695
rect 13964 5664 14197 5692
rect 13964 5652 13970 5664
rect 14185 5661 14197 5664
rect 14231 5692 14243 5695
rect 18598 5692 18604 5704
rect 14231 5664 17448 5692
rect 18559 5664 18604 5692
rect 14231 5661 14243 5664
rect 14185 5655 14243 5661
rect 15565 5627 15623 5633
rect 15565 5593 15577 5627
rect 15611 5624 15623 5627
rect 16482 5624 16488 5636
rect 15611 5596 16488 5624
rect 15611 5593 15623 5596
rect 15565 5587 15623 5593
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 16022 5556 16028 5568
rect 13832 5528 16028 5556
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 16577 5559 16635 5565
rect 16577 5525 16589 5559
rect 16623 5556 16635 5559
rect 17310 5556 17316 5568
rect 16623 5528 17316 5556
rect 16623 5525 16635 5528
rect 16577 5519 16635 5525
rect 17310 5516 17316 5528
rect 17368 5516 17374 5568
rect 17420 5556 17448 5664
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 18708 5701 18736 5732
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 19702 5760 19708 5772
rect 19392 5732 19708 5760
rect 19392 5720 19398 5732
rect 19702 5720 19708 5732
rect 19760 5720 19766 5772
rect 20070 5720 20076 5772
rect 20128 5760 20134 5772
rect 21358 5760 21364 5772
rect 20128 5732 21364 5760
rect 20128 5720 20134 5732
rect 21358 5720 21364 5732
rect 21416 5760 21422 5772
rect 21525 5763 21583 5769
rect 21525 5760 21537 5763
rect 21416 5732 21537 5760
rect 21416 5720 21422 5732
rect 21525 5729 21537 5732
rect 21571 5729 21583 5763
rect 21525 5723 21583 5729
rect 24121 5763 24179 5769
rect 24121 5729 24133 5763
rect 24167 5760 24179 5763
rect 24210 5760 24216 5772
rect 24167 5732 24216 5760
rect 24167 5729 24179 5732
rect 24121 5723 24179 5729
rect 24210 5720 24216 5732
rect 24268 5760 24274 5772
rect 24486 5760 24492 5772
rect 24268 5732 24492 5760
rect 24268 5720 24274 5732
rect 24486 5720 24492 5732
rect 24544 5720 24550 5772
rect 25222 5720 25228 5772
rect 25280 5760 25286 5772
rect 25317 5763 25375 5769
rect 25317 5760 25329 5763
rect 25280 5732 25329 5760
rect 25280 5720 25286 5732
rect 25317 5729 25329 5732
rect 25363 5760 25375 5763
rect 25866 5760 25872 5772
rect 25363 5732 25872 5760
rect 25363 5729 25375 5732
rect 25317 5723 25375 5729
rect 25866 5720 25872 5732
rect 25924 5720 25930 5772
rect 18693 5695 18751 5701
rect 18693 5661 18705 5695
rect 18739 5692 18751 5695
rect 21269 5695 21327 5701
rect 18739 5664 20300 5692
rect 18739 5661 18751 5664
rect 18693 5655 18751 5661
rect 18141 5627 18199 5633
rect 18141 5593 18153 5627
rect 18187 5624 18199 5627
rect 19242 5624 19248 5636
rect 18187 5596 19248 5624
rect 18187 5593 18199 5596
rect 18141 5587 18199 5593
rect 19242 5584 19248 5596
rect 19300 5584 19306 5636
rect 19613 5627 19671 5633
rect 19613 5593 19625 5627
rect 19659 5624 19671 5627
rect 20070 5624 20076 5636
rect 19659 5596 20076 5624
rect 19659 5593 19671 5596
rect 19613 5587 19671 5593
rect 20070 5584 20076 5596
rect 20128 5584 20134 5636
rect 20272 5568 20300 5664
rect 21269 5661 21281 5695
rect 21315 5661 21327 5695
rect 21269 5655 21327 5661
rect 24397 5695 24455 5701
rect 24397 5661 24409 5695
rect 24443 5692 24455 5695
rect 24670 5692 24676 5704
rect 24443 5664 24676 5692
rect 24443 5661 24455 5664
rect 24397 5655 24455 5661
rect 19518 5556 19524 5568
rect 17420 5528 19524 5556
rect 19518 5516 19524 5528
rect 19576 5516 19582 5568
rect 20254 5556 20260 5568
rect 20215 5528 20260 5556
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20622 5516 20628 5568
rect 20680 5556 20686 5568
rect 21284 5556 21312 5655
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 25130 5692 25136 5704
rect 25091 5664 25136 5692
rect 25130 5652 25136 5664
rect 25188 5652 25194 5704
rect 24857 5627 24915 5633
rect 24857 5593 24869 5627
rect 24903 5624 24915 5627
rect 25038 5624 25044 5636
rect 24903 5596 25044 5624
rect 24903 5593 24915 5596
rect 24857 5587 24915 5593
rect 25038 5584 25044 5596
rect 25096 5624 25102 5636
rect 25958 5624 25964 5636
rect 25096 5596 25964 5624
rect 25096 5584 25102 5596
rect 25958 5584 25964 5596
rect 26016 5584 26022 5636
rect 22002 5556 22008 5568
rect 20680 5528 22008 5556
rect 20680 5516 20686 5528
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 23845 5559 23903 5565
rect 23845 5525 23857 5559
rect 23891 5556 23903 5559
rect 23934 5556 23940 5568
rect 23891 5528 23940 5556
rect 23891 5525 23903 5528
rect 23845 5519 23903 5525
rect 23934 5516 23940 5528
rect 23992 5516 23998 5568
rect 25314 5516 25320 5568
rect 25372 5556 25378 5568
rect 25501 5559 25559 5565
rect 25501 5556 25513 5559
rect 25372 5528 25513 5556
rect 25372 5516 25378 5528
rect 25501 5525 25513 5528
rect 25547 5525 25559 5559
rect 26234 5556 26240 5568
rect 26195 5528 26240 5556
rect 25501 5519 25559 5525
rect 26234 5516 26240 5528
rect 26292 5516 26298 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1486 5352 1492 5364
rect 1447 5324 1492 5352
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 2498 5352 2504 5364
rect 2459 5324 2504 5352
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 4614 5352 4620 5364
rect 4387 5324 4620 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 4614 5312 4620 5324
rect 4672 5352 4678 5364
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 4672 5324 5273 5352
rect 4672 5312 4678 5324
rect 5261 5321 5273 5324
rect 5307 5321 5319 5355
rect 5261 5315 5319 5321
rect 6917 5355 6975 5361
rect 6917 5321 6929 5355
rect 6963 5352 6975 5355
rect 8202 5352 8208 5364
rect 6963 5324 8208 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 10042 5352 10048 5364
rect 10003 5324 10048 5352
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11422 5352 11428 5364
rect 11379 5324 11428 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 11606 5352 11612 5364
rect 11567 5324 11612 5352
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 13725 5355 13783 5361
rect 13725 5321 13737 5355
rect 13771 5352 13783 5355
rect 13906 5352 13912 5364
rect 13771 5324 13912 5352
rect 13771 5321 13783 5324
rect 13725 5315 13783 5321
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 14093 5355 14151 5361
rect 14093 5321 14105 5355
rect 14139 5352 14151 5355
rect 14366 5352 14372 5364
rect 14139 5324 14372 5352
rect 14139 5321 14151 5324
rect 14093 5315 14151 5321
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 17678 5352 17684 5364
rect 17543 5324 17684 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 7282 5284 7288 5296
rect 5684 5256 7288 5284
rect 5684 5244 5690 5256
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 8481 5287 8539 5293
rect 8481 5253 8493 5287
rect 8527 5284 8539 5287
rect 12526 5284 12532 5296
rect 8527 5256 10456 5284
rect 12487 5256 12532 5284
rect 8527 5253 8539 5256
rect 8481 5247 8539 5253
rect 1946 5216 1952 5228
rect 1907 5188 1952 5216
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2958 5216 2964 5228
rect 2919 5188 2964 5216
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5216 5779 5219
rect 6730 5216 6736 5228
rect 5767 5188 6736 5216
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5216 7987 5219
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 7975 5188 9045 5216
rect 7975 5185 7987 5188
rect 7929 5179 7987 5185
rect 9033 5185 9045 5188
rect 9079 5216 9091 5219
rect 9398 5216 9404 5228
rect 9079 5188 9404 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 10428 5225 10456 5256
rect 12526 5244 12532 5256
rect 12584 5244 12590 5296
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5216 10471 5219
rect 11606 5216 11612 5228
rect 10459 5188 11612 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13044 5188 13089 5216
rect 13044 5176 13050 5188
rect 13538 5176 13544 5228
rect 13596 5216 13602 5228
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 13596 5188 14381 5216
rect 13596 5176 13602 5188
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 3234 5157 3240 5160
rect 3228 5148 3240 5157
rect 3160 5120 3240 5148
rect 2041 5083 2099 5089
rect 2041 5049 2053 5083
rect 2087 5080 2099 5083
rect 2682 5080 2688 5092
rect 2087 5052 2688 5080
rect 2087 5049 2099 5052
rect 2041 5043 2099 5049
rect 2682 5040 2688 5052
rect 2740 5080 2746 5092
rect 3160 5080 3188 5120
rect 3228 5111 3240 5120
rect 3234 5108 3240 5111
rect 3292 5108 3298 5160
rect 5442 5148 5448 5160
rect 5403 5120 5448 5148
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 5810 5148 5816 5160
rect 5592 5120 5816 5148
rect 5592 5108 5598 5120
rect 5810 5108 5816 5120
rect 5868 5148 5874 5160
rect 7469 5151 7527 5157
rect 7469 5148 7481 5151
rect 5868 5120 7481 5148
rect 5868 5108 5874 5120
rect 7469 5117 7481 5120
rect 7515 5148 7527 5151
rect 8110 5148 8116 5160
rect 7515 5120 8116 5148
rect 7515 5117 7527 5120
rect 7469 5111 7527 5117
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 9769 5151 9827 5157
rect 9769 5117 9781 5151
rect 9815 5148 9827 5151
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 9815 5120 10609 5148
rect 9815 5117 9827 5120
rect 9769 5111 9827 5117
rect 10597 5117 10609 5120
rect 10643 5148 10655 5151
rect 10778 5148 10784 5160
rect 10643 5120 10784 5148
rect 10643 5117 10655 5120
rect 10597 5111 10655 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 13004 5148 13032 5176
rect 12299 5120 13032 5148
rect 14384 5148 14412 5179
rect 14458 5148 14464 5160
rect 14384 5120 14464 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5148 16911 5151
rect 17512 5148 17540 5315
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 17862 5352 17868 5364
rect 17823 5324 17868 5352
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 18141 5355 18199 5361
rect 18141 5321 18153 5355
rect 18187 5352 18199 5355
rect 18598 5352 18604 5364
rect 18187 5324 18604 5352
rect 18187 5321 18199 5324
rect 18141 5315 18199 5321
rect 18598 5312 18604 5324
rect 18656 5312 18662 5364
rect 19702 5352 19708 5364
rect 19663 5324 19708 5352
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 20622 5352 20628 5364
rect 19996 5324 20628 5352
rect 18322 5244 18328 5296
rect 18380 5284 18386 5296
rect 19429 5287 19487 5293
rect 19429 5284 19441 5287
rect 18380 5256 19441 5284
rect 18380 5244 18386 5256
rect 19429 5253 19441 5256
rect 19475 5284 19487 5287
rect 19996 5284 20024 5324
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 21358 5352 21364 5364
rect 21319 5324 21364 5352
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 22002 5352 22008 5364
rect 21963 5324 22008 5352
rect 22002 5312 22008 5324
rect 22060 5312 22066 5364
rect 23109 5355 23167 5361
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23382 5352 23388 5364
rect 23155 5324 23388 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23382 5312 23388 5324
rect 23440 5312 23446 5364
rect 23753 5355 23811 5361
rect 23753 5321 23765 5355
rect 23799 5352 23811 5355
rect 24854 5352 24860 5364
rect 23799 5324 24860 5352
rect 23799 5321 23811 5324
rect 23753 5315 23811 5321
rect 24854 5312 24860 5324
rect 24912 5312 24918 5364
rect 25866 5312 25872 5364
rect 25924 5352 25930 5364
rect 25961 5355 26019 5361
rect 25961 5352 25973 5355
rect 25924 5324 25973 5352
rect 25924 5312 25930 5324
rect 25961 5321 25973 5324
rect 26007 5321 26019 5355
rect 25961 5315 26019 5321
rect 19475 5256 20024 5284
rect 19475 5253 19487 5256
rect 19429 5247 19487 5253
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 18506 5216 18512 5228
rect 17828 5188 18512 5216
rect 17828 5176 17834 5188
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 18690 5216 18696 5228
rect 18651 5188 18696 5216
rect 18690 5176 18696 5188
rect 18748 5176 18754 5228
rect 19996 5225 20024 5256
rect 23014 5244 23020 5296
rect 23072 5284 23078 5296
rect 26694 5284 26700 5296
rect 23072 5256 26700 5284
rect 23072 5244 23078 5256
rect 26694 5244 26700 5256
rect 26752 5244 26758 5296
rect 19981 5219 20039 5225
rect 19981 5185 19993 5219
rect 20027 5185 20039 5219
rect 19981 5179 20039 5185
rect 22278 5176 22284 5228
rect 22336 5216 22342 5228
rect 24305 5219 24363 5225
rect 24305 5216 24317 5219
rect 22336 5188 24317 5216
rect 22336 5176 22342 5188
rect 24305 5185 24317 5188
rect 24351 5216 24363 5219
rect 24765 5219 24823 5225
rect 24765 5216 24777 5219
rect 24351 5188 24777 5216
rect 24351 5185 24363 5188
rect 24305 5179 24363 5185
rect 24765 5185 24777 5188
rect 24811 5185 24823 5219
rect 25498 5216 25504 5228
rect 25459 5188 25504 5216
rect 24765 5179 24823 5185
rect 25498 5176 25504 5188
rect 25556 5176 25562 5228
rect 20254 5157 20260 5160
rect 20248 5148 20260 5157
rect 16899 5120 17540 5148
rect 20215 5120 20260 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 20248 5111 20260 5120
rect 20254 5108 20260 5111
rect 20312 5108 20318 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22296 5120 22477 5148
rect 22296 5092 22324 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 23474 5108 23480 5160
rect 23532 5148 23538 5160
rect 23532 5120 24164 5148
rect 23532 5108 23538 5120
rect 2740 5052 3188 5080
rect 4985 5083 5043 5089
rect 2740 5040 2746 5052
rect 4985 5049 4997 5083
rect 5031 5080 5043 5083
rect 6914 5080 6920 5092
rect 5031 5052 6920 5080
rect 5031 5049 5043 5052
rect 4985 5043 5043 5049
rect 1949 5015 2007 5021
rect 1949 4981 1961 5015
rect 1995 5012 2007 5015
rect 2130 5012 2136 5024
rect 1995 4984 2136 5012
rect 1995 4981 2007 4984
rect 1949 4975 2007 4981
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2869 5015 2927 5021
rect 2869 4981 2881 5015
rect 2915 5012 2927 5015
rect 2958 5012 2964 5024
rect 2915 4984 2964 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 2958 4972 2964 4984
rect 3016 5012 3022 5024
rect 3234 5012 3240 5024
rect 3016 4984 3240 5012
rect 3016 4972 3022 4984
rect 3234 4972 3240 4984
rect 3292 5012 3298 5024
rect 4798 5012 4804 5024
rect 3292 4984 4804 5012
rect 3292 4972 3298 4984
rect 4798 4972 4804 4984
rect 4856 5012 4862 5024
rect 5000 5012 5028 5043
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 7193 5083 7251 5089
rect 7193 5049 7205 5083
rect 7239 5049 7251 5083
rect 7193 5043 7251 5049
rect 8297 5083 8355 5089
rect 8297 5049 8309 5083
rect 8343 5080 8355 5083
rect 8754 5080 8760 5092
rect 8343 5052 8760 5080
rect 8343 5049 8355 5052
rect 8297 5043 8355 5049
rect 6270 5012 6276 5024
rect 4856 4984 5028 5012
rect 6231 4984 6276 5012
rect 4856 4972 4862 4984
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 6546 4972 6552 4984
rect 6604 5012 6610 5024
rect 7208 5012 7236 5043
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 8938 5080 8944 5092
rect 8899 5052 8944 5080
rect 8938 5040 8944 5052
rect 8996 5040 9002 5092
rect 13078 5080 13084 5092
rect 13039 5052 13084 5080
rect 13078 5040 13084 5052
rect 13136 5040 13142 5092
rect 14636 5083 14694 5089
rect 14636 5049 14648 5083
rect 14682 5080 14694 5083
rect 14734 5080 14740 5092
rect 14682 5052 14740 5080
rect 14682 5049 14694 5052
rect 14636 5043 14694 5049
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 16485 5083 16543 5089
rect 16485 5080 16497 5083
rect 15304 5052 16497 5080
rect 6604 4984 7236 5012
rect 7377 5015 7435 5021
rect 6604 4972 6610 4984
rect 7377 4981 7389 5015
rect 7423 5012 7435 5015
rect 7650 5012 7656 5024
rect 7423 4984 7656 5012
rect 7423 4981 7435 4984
rect 7377 4975 7435 4981
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 10192 4984 10517 5012
rect 10192 4972 10198 4984
rect 10505 4981 10517 4984
rect 10551 5012 10563 5015
rect 11054 5012 11060 5024
rect 10551 4984 11060 5012
rect 10551 4981 10563 4984
rect 10505 4975 10563 4981
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 12989 5015 13047 5021
rect 12989 5012 13001 5015
rect 12676 4984 13001 5012
rect 12676 4972 12682 4984
rect 12989 4981 13001 4984
rect 13035 4981 13047 5015
rect 12989 4975 13047 4981
rect 13906 4972 13912 5024
rect 13964 5012 13970 5024
rect 15304 5012 15332 5052
rect 16485 5049 16497 5052
rect 16531 5080 16543 5083
rect 16758 5080 16764 5092
rect 16531 5052 16764 5080
rect 16531 5049 16543 5052
rect 16485 5043 16543 5049
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 18598 5080 18604 5092
rect 18559 5052 18604 5080
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 22278 5080 22284 5092
rect 22239 5052 22284 5080
rect 22278 5040 22284 5052
rect 22336 5040 22342 5092
rect 24029 5083 24087 5089
rect 24029 5049 24041 5083
rect 24075 5049 24087 5083
rect 24136 5080 24164 5120
rect 24670 5108 24676 5160
rect 24728 5148 24734 5160
rect 25041 5151 25099 5157
rect 25041 5148 25053 5151
rect 24728 5120 25053 5148
rect 24728 5108 24734 5120
rect 25041 5117 25053 5120
rect 25087 5117 25099 5151
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 25041 5111 25099 5117
rect 25222 5108 25228 5120
rect 25280 5108 25286 5160
rect 25498 5080 25504 5092
rect 24136 5052 25504 5080
rect 24029 5043 24087 5049
rect 13964 4984 15332 5012
rect 13964 4972 13970 4984
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15749 5015 15807 5021
rect 15749 5012 15761 5015
rect 15436 4984 15761 5012
rect 15436 4972 15442 4984
rect 15749 4981 15761 4984
rect 15795 4981 15807 5015
rect 15749 4975 15807 4981
rect 17037 5015 17095 5021
rect 17037 4981 17049 5015
rect 17083 5012 17095 5015
rect 17310 5012 17316 5024
rect 17083 4984 17316 5012
rect 17083 4981 17095 4984
rect 17037 4975 17095 4981
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 19978 4972 19984 5024
rect 20036 5012 20042 5024
rect 22370 5012 22376 5024
rect 20036 4984 22376 5012
rect 20036 4972 20042 4984
rect 22370 4972 22376 4984
rect 22428 4972 22434 5024
rect 22646 5012 22652 5024
rect 22607 4984 22652 5012
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 23474 5012 23480 5024
rect 23435 4984 23480 5012
rect 23474 4972 23480 4984
rect 23532 5012 23538 5024
rect 24044 5012 24072 5043
rect 25498 5040 25504 5052
rect 25556 5040 25562 5092
rect 24210 5012 24216 5024
rect 23532 4984 24072 5012
rect 24171 4984 24216 5012
rect 23532 4972 23538 4984
rect 24210 4972 24216 4984
rect 24268 4972 24274 5024
rect 26326 5012 26332 5024
rect 26287 4984 26332 5012
rect 26326 4972 26332 4984
rect 26384 4972 26390 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 2133 4811 2191 4817
rect 2133 4777 2145 4811
rect 2179 4808 2191 4811
rect 2498 4808 2504 4820
rect 2179 4780 2504 4808
rect 2179 4777 2191 4780
rect 2133 4771 2191 4777
rect 2498 4768 2504 4780
rect 2556 4808 2562 4820
rect 5074 4808 5080 4820
rect 2556 4780 2912 4808
rect 5035 4780 5080 4808
rect 2556 4768 2562 4780
rect 2884 4749 2912 4780
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 5721 4811 5779 4817
rect 5721 4777 5733 4811
rect 5767 4808 5779 4811
rect 5810 4808 5816 4820
rect 5767 4780 5816 4808
rect 5767 4777 5779 4780
rect 5721 4771 5779 4777
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 5994 4768 6000 4820
rect 6052 4808 6058 4820
rect 6362 4808 6368 4820
rect 6052 4780 6368 4808
rect 6052 4768 6058 4780
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 6914 4808 6920 4820
rect 6875 4780 6920 4808
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 8294 4768 8300 4820
rect 8352 4768 8358 4820
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 8846 4808 8852 4820
rect 8619 4780 8852 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 9125 4811 9183 4817
rect 9125 4777 9137 4811
rect 9171 4808 9183 4811
rect 9398 4808 9404 4820
rect 9171 4780 9404 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 9398 4768 9404 4780
rect 9456 4808 9462 4820
rect 11238 4808 11244 4820
rect 9456 4780 11244 4808
rect 9456 4768 9462 4780
rect 2777 4743 2835 4749
rect 2777 4709 2789 4743
rect 2823 4709 2835 4743
rect 2777 4703 2835 4709
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4709 2927 4743
rect 2869 4703 2927 4709
rect 2792 4672 2820 4703
rect 3510 4700 3516 4752
rect 3568 4740 3574 4752
rect 4617 4743 4675 4749
rect 4617 4740 4629 4743
rect 3568 4712 4629 4740
rect 3568 4700 3574 4712
rect 4617 4709 4629 4712
rect 4663 4740 4675 4743
rect 6546 4740 6552 4752
rect 4663 4712 6552 4740
rect 4663 4709 4675 4712
rect 4617 4703 4675 4709
rect 6546 4700 6552 4712
rect 6604 4700 6610 4752
rect 7929 4743 7987 4749
rect 7929 4709 7941 4743
rect 7975 4740 7987 4743
rect 8312 4740 8340 4768
rect 10042 4740 10048 4752
rect 7975 4712 8708 4740
rect 10003 4712 10048 4740
rect 7975 4709 7987 4712
rect 7929 4703 7987 4709
rect 4154 4672 4160 4684
rect 2792 4644 4160 4672
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 5994 4632 6000 4684
rect 6052 4672 6058 4684
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 6052 4644 6193 4672
rect 6052 4632 6058 4644
rect 6181 4641 6193 4644
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 8680 4681 8708 4712
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 10226 4740 10232 4752
rect 10187 4712 10232 4740
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 10336 4749 10364 4780
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11606 4808 11612 4820
rect 11567 4780 11612 4808
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 12621 4811 12679 4817
rect 12621 4777 12633 4811
rect 12667 4808 12679 4811
rect 12802 4808 12808 4820
rect 12667 4780 12808 4808
rect 12667 4777 12679 4780
rect 12621 4771 12679 4777
rect 12802 4768 12808 4780
rect 12860 4808 12866 4820
rect 13630 4808 13636 4820
rect 12860 4780 13636 4808
rect 12860 4768 12866 4780
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14458 4768 14464 4820
rect 14516 4808 14522 4820
rect 14645 4811 14703 4817
rect 14645 4808 14657 4811
rect 14516 4780 14657 4808
rect 14516 4768 14522 4780
rect 14645 4777 14657 4780
rect 14691 4808 14703 4811
rect 14734 4808 14740 4820
rect 14691 4780 14740 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 15252 4780 15853 4808
rect 15252 4768 15258 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 15841 4771 15899 4777
rect 16577 4811 16635 4817
rect 16577 4777 16589 4811
rect 16623 4808 16635 4811
rect 17402 4808 17408 4820
rect 16623 4780 17408 4808
rect 16623 4777 16635 4780
rect 16577 4771 16635 4777
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 19705 4811 19763 4817
rect 19705 4777 19717 4811
rect 19751 4808 19763 4811
rect 20254 4808 20260 4820
rect 19751 4780 20260 4808
rect 19751 4777 19763 4780
rect 19705 4771 19763 4777
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 21358 4768 21364 4820
rect 21416 4808 21422 4820
rect 22281 4811 22339 4817
rect 22281 4808 22293 4811
rect 21416 4780 22293 4808
rect 21416 4768 21422 4780
rect 22281 4777 22293 4780
rect 22327 4777 22339 4811
rect 22281 4771 22339 4777
rect 23845 4811 23903 4817
rect 23845 4777 23857 4811
rect 23891 4808 23903 4811
rect 24118 4808 24124 4820
rect 23891 4780 24124 4808
rect 23891 4777 23903 4780
rect 23845 4771 23903 4777
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 24581 4811 24639 4817
rect 24581 4777 24593 4811
rect 24627 4808 24639 4811
rect 25130 4808 25136 4820
rect 24627 4780 25136 4808
rect 24627 4777 24639 4780
rect 24581 4771 24639 4777
rect 25130 4768 25136 4780
rect 25188 4768 25194 4820
rect 25222 4768 25228 4820
rect 25280 4808 25286 4820
rect 25777 4811 25835 4817
rect 25777 4808 25789 4811
rect 25280 4780 25789 4808
rect 25280 4768 25286 4780
rect 25777 4777 25789 4780
rect 25823 4777 25835 4811
rect 26234 4808 26240 4820
rect 26195 4780 26240 4808
rect 25777 4771 25835 4777
rect 26234 4768 26240 4780
rect 26292 4768 26298 4820
rect 10321 4743 10379 4749
rect 10321 4709 10333 4743
rect 10367 4709 10379 4743
rect 10778 4740 10784 4752
rect 10739 4712 10784 4740
rect 10321 4703 10379 4709
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 13541 4743 13599 4749
rect 13541 4709 13553 4743
rect 13587 4740 13599 4743
rect 13814 4740 13820 4752
rect 13587 4712 13820 4740
rect 13587 4709 13599 4712
rect 13541 4703 13599 4709
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 14185 4743 14243 4749
rect 14185 4709 14197 4743
rect 14231 4709 14243 4743
rect 14185 4703 14243 4709
rect 14277 4743 14335 4749
rect 14277 4709 14289 4743
rect 14323 4740 14335 4743
rect 15378 4740 15384 4752
rect 14323 4712 15384 4740
rect 14323 4709 14335 4712
rect 14277 4703 14335 4709
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 8352 4644 8401 4672
rect 8352 4632 8358 4644
rect 8389 4641 8401 4644
rect 8435 4641 8447 4675
rect 8389 4635 8447 4641
rect 8665 4675 8723 4681
rect 8665 4641 8677 4675
rect 8711 4672 8723 4675
rect 10796 4672 10824 4700
rect 8711 4644 10824 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 10870 4632 10876 4684
rect 10928 4672 10934 4684
rect 11238 4672 11244 4684
rect 10928 4644 11244 4672
rect 10928 4632 10934 4644
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 14200 4672 14228 4703
rect 15378 4700 15384 4712
rect 15436 4700 15442 4752
rect 15654 4740 15660 4752
rect 15615 4712 15660 4740
rect 15654 4700 15660 4712
rect 15712 4700 15718 4752
rect 16666 4740 16672 4752
rect 15755 4712 16672 4740
rect 14550 4672 14556 4684
rect 12308 4644 12756 4672
rect 14200 4644 14556 4672
rect 12308 4632 12314 4644
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 2777 4607 2835 4613
rect 2777 4604 2789 4607
rect 2556 4576 2789 4604
rect 2556 4564 2562 4576
rect 2777 4573 2789 4576
rect 2823 4604 2835 4607
rect 3326 4604 3332 4616
rect 2823 4576 3332 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4614 4604 4620 4616
rect 4028 4576 4620 4604
rect 4028 4564 4034 4576
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 2314 4536 2320 4548
rect 2275 4508 2320 4536
rect 2314 4496 2320 4508
rect 2372 4496 2378 4548
rect 4338 4536 4344 4548
rect 3436 4508 4344 4536
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4468 1734 4480
rect 3436 4477 3464 4508
rect 4338 4496 4344 4508
rect 4396 4536 4402 4548
rect 4724 4536 4752 4567
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6328 4576 6469 4604
rect 6328 4564 6334 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 10226 4604 10232 4616
rect 9732 4576 10232 4604
rect 9732 4564 9738 4576
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 12618 4604 12624 4616
rect 12579 4576 12624 4604
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 12728 4613 12756 4644
rect 14550 4632 14556 4644
rect 14608 4672 14614 4684
rect 15755 4672 15783 4712
rect 16666 4700 16672 4712
rect 16724 4700 16730 4752
rect 18592 4743 18650 4749
rect 18592 4709 18604 4743
rect 18638 4740 18650 4743
rect 18690 4740 18696 4752
rect 18638 4712 18696 4740
rect 18638 4709 18650 4712
rect 18592 4703 18650 4709
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 21174 4700 21180 4752
rect 21232 4740 21238 4752
rect 21453 4743 21511 4749
rect 21453 4740 21465 4743
rect 21232 4712 21465 4740
rect 21232 4700 21238 4712
rect 21453 4709 21465 4712
rect 21499 4709 21511 4743
rect 22830 4740 22836 4752
rect 22791 4712 22836 4740
rect 21453 4703 21511 4709
rect 22830 4700 22836 4712
rect 22888 4700 22894 4752
rect 23014 4740 23020 4752
rect 22975 4712 23020 4740
rect 23014 4700 23020 4712
rect 23072 4700 23078 4752
rect 23109 4743 23167 4749
rect 23109 4709 23121 4743
rect 23155 4740 23167 4743
rect 24486 4740 24492 4752
rect 23155 4712 24492 4740
rect 23155 4709 23167 4712
rect 23109 4703 23167 4709
rect 14608 4644 15783 4672
rect 14608 4632 14614 4644
rect 16298 4632 16304 4684
rect 16356 4672 16362 4684
rect 16945 4675 17003 4681
rect 16945 4672 16957 4675
rect 16356 4644 16957 4672
rect 16356 4632 16362 4644
rect 16945 4641 16957 4644
rect 16991 4641 17003 4675
rect 18138 4672 18144 4684
rect 18051 4644 18144 4672
rect 16945 4635 17003 4641
rect 18138 4632 18144 4644
rect 18196 4672 18202 4684
rect 18322 4672 18328 4684
rect 18196 4644 18328 4672
rect 18196 4632 18202 4644
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 20898 4632 20904 4684
rect 20956 4672 20962 4684
rect 21358 4672 21364 4684
rect 20956 4644 21364 4672
rect 20956 4632 20962 4644
rect 21358 4632 21364 4644
rect 21416 4632 21422 4684
rect 22002 4672 22008 4684
rect 21468 4644 22008 4672
rect 12713 4607 12771 4613
rect 12713 4573 12725 4607
rect 12759 4604 12771 4607
rect 12986 4604 12992 4616
rect 12759 4576 12992 4604
rect 12759 4573 12771 4576
rect 12713 4567 12771 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 14185 4607 14243 4613
rect 14185 4573 14197 4607
rect 14231 4573 14243 4607
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 14185 4567 14243 4573
rect 15028 4576 15945 4604
rect 5442 4536 5448 4548
rect 4396 4508 5448 4536
rect 4396 4496 4402 4508
rect 5442 4496 5448 4508
rect 5500 4496 5506 4548
rect 5905 4539 5963 4545
rect 5905 4505 5917 4539
rect 5951 4536 5963 4539
rect 7650 4536 7656 4548
rect 5951 4508 7656 4536
rect 5951 4505 5963 4508
rect 5905 4499 5963 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 8113 4539 8171 4545
rect 8113 4505 8125 4539
rect 8159 4536 8171 4539
rect 8938 4536 8944 4548
rect 8159 4508 8944 4536
rect 8159 4505 8171 4508
rect 8113 4499 8171 4505
rect 8938 4496 8944 4508
rect 8996 4496 9002 4548
rect 9766 4536 9772 4548
rect 9727 4508 9772 4536
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 12158 4536 12164 4548
rect 12119 4508 12164 4536
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 12434 4496 12440 4548
rect 12492 4536 12498 4548
rect 13725 4539 13783 4545
rect 13725 4536 13737 4539
rect 12492 4508 13737 4536
rect 12492 4496 12498 4508
rect 13725 4505 13737 4508
rect 13771 4536 13783 4539
rect 13814 4536 13820 4548
rect 13771 4508 13820 4536
rect 13771 4505 13783 4508
rect 13725 4499 13783 4505
rect 13814 4496 13820 4508
rect 13872 4496 13878 4548
rect 14200 4536 14228 4567
rect 14458 4536 14464 4548
rect 14200 4508 14464 4536
rect 14458 4496 14464 4508
rect 14516 4496 14522 4548
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 1728 4440 3433 4468
rect 1728 4428 1734 4440
rect 3421 4437 3433 4440
rect 3467 4437 3479 4471
rect 3421 4431 3479 4437
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4062 4468 4068 4480
rect 3927 4440 4068 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 7282 4468 7288 4480
rect 4212 4440 4257 4468
rect 7243 4440 7288 4468
rect 4212 4428 4218 4440
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 13173 4471 13231 4477
rect 13173 4437 13185 4471
rect 13219 4468 13231 4471
rect 13998 4468 14004 4480
rect 13219 4440 14004 4468
rect 13219 4437 13231 4440
rect 13173 4431 13231 4437
rect 13998 4428 14004 4440
rect 14056 4468 14062 4480
rect 15028 4477 15056 4576
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 16482 4564 16488 4616
rect 16540 4564 16546 4616
rect 17126 4604 17132 4616
rect 17087 4576 17132 4604
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 21468 4613 21496 4644
rect 22002 4632 22008 4644
rect 22060 4632 22066 4684
rect 22186 4632 22192 4684
rect 22244 4672 22250 4684
rect 23124 4672 23152 4703
rect 24486 4700 24492 4712
rect 24544 4700 24550 4752
rect 22244 4644 23152 4672
rect 22244 4632 22250 4644
rect 24118 4632 24124 4684
rect 24176 4672 24182 4684
rect 24673 4675 24731 4681
rect 24673 4672 24685 4675
rect 24176 4644 24685 4672
rect 24176 4632 24182 4644
rect 24673 4641 24685 4644
rect 24719 4641 24731 4675
rect 24673 4635 24731 4641
rect 21453 4607 21511 4613
rect 19484 4576 21128 4604
rect 19484 4564 19490 4576
rect 15381 4539 15439 4545
rect 15381 4505 15393 4539
rect 15427 4536 15439 4539
rect 15838 4536 15844 4548
rect 15427 4508 15844 4536
rect 15427 4505 15439 4508
rect 15381 4499 15439 4505
rect 15838 4496 15844 4508
rect 15896 4536 15902 4548
rect 16500 4536 16528 4564
rect 20990 4536 20996 4548
rect 15896 4508 16528 4536
rect 20951 4508 20996 4536
rect 15896 4496 15902 4508
rect 20990 4496 20996 4508
rect 21048 4496 21054 4548
rect 21100 4536 21128 4576
rect 21453 4573 21465 4607
rect 21499 4573 21511 4607
rect 21453 4567 21511 4573
rect 21542 4564 21548 4616
rect 21600 4604 21606 4616
rect 21913 4607 21971 4613
rect 21913 4604 21925 4607
rect 21600 4576 21925 4604
rect 21600 4564 21606 4576
rect 21913 4573 21925 4576
rect 21959 4573 21971 4607
rect 24578 4604 24584 4616
rect 24539 4576 24584 4604
rect 21913 4567 21971 4573
rect 24578 4564 24584 4576
rect 24636 4564 24642 4616
rect 22462 4536 22468 4548
rect 21100 4508 22468 4536
rect 22462 4496 22468 4508
rect 22520 4496 22526 4548
rect 24121 4539 24179 4545
rect 24121 4505 24133 4539
rect 24167 4536 24179 4539
rect 24210 4536 24216 4548
rect 24167 4508 24216 4536
rect 24167 4505 24179 4508
rect 24121 4499 24179 4505
rect 24210 4496 24216 4508
rect 24268 4536 24274 4548
rect 25041 4539 25099 4545
rect 25041 4536 25053 4539
rect 24268 4508 25053 4536
rect 24268 4496 24274 4508
rect 25041 4505 25053 4508
rect 25087 4505 25099 4539
rect 25041 4499 25099 4505
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14056 4440 15025 4468
rect 14056 4428 14062 4440
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15013 4431 15071 4437
rect 17773 4471 17831 4477
rect 17773 4437 17785 4471
rect 17819 4468 17831 4471
rect 17862 4468 17868 4480
rect 17819 4440 17868 4468
rect 17819 4437 17831 4440
rect 17773 4431 17831 4437
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 20622 4468 20628 4480
rect 20583 4440 20628 4468
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 22554 4428 22560 4480
rect 22612 4468 22618 4480
rect 25406 4468 25412 4480
rect 22612 4440 22657 4468
rect 25367 4440 25412 4468
rect 22612 4428 22618 4440
rect 25406 4428 25412 4440
rect 25464 4428 25470 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2130 4264 2136 4276
rect 2091 4236 2136 4264
rect 2130 4224 2136 4236
rect 2188 4224 2194 4276
rect 3234 4264 3240 4276
rect 3195 4236 3240 4264
rect 3234 4224 3240 4236
rect 3292 4224 3298 4276
rect 5442 4264 5448 4276
rect 5403 4236 5448 4264
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 6362 4264 6368 4276
rect 6323 4236 6368 4264
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 7101 4267 7159 4273
rect 7101 4264 7113 4267
rect 7064 4236 7113 4264
rect 7064 4224 7070 4236
rect 7101 4233 7113 4236
rect 7147 4233 7159 4267
rect 7101 4227 7159 4233
rect 8481 4267 8539 4273
rect 8481 4233 8493 4267
rect 8527 4264 8539 4267
rect 8846 4264 8852 4276
rect 8527 4236 8852 4264
rect 8527 4233 8539 4236
rect 8481 4227 8539 4233
rect 8846 4224 8852 4236
rect 8904 4224 8910 4276
rect 9033 4267 9091 4273
rect 9033 4233 9045 4267
rect 9079 4264 9091 4267
rect 10134 4264 10140 4276
rect 9079 4236 10140 4264
rect 9079 4233 9091 4236
rect 9033 4227 9091 4233
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 12158 4264 12164 4276
rect 12071 4236 12164 4264
rect 12158 4224 12164 4236
rect 12216 4264 12222 4276
rect 12618 4264 12624 4276
rect 12216 4236 12624 4264
rect 12216 4224 12222 4236
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 12713 4267 12771 4273
rect 12713 4233 12725 4267
rect 12759 4264 12771 4267
rect 12802 4264 12808 4276
rect 12759 4236 12808 4264
rect 12759 4233 12771 4236
rect 12713 4227 12771 4233
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 13449 4267 13507 4273
rect 13449 4233 13461 4267
rect 13495 4264 13507 4267
rect 14182 4264 14188 4276
rect 13495 4236 14188 4264
rect 13495 4233 13507 4236
rect 13449 4227 13507 4233
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 14369 4267 14427 4273
rect 14369 4233 14381 4267
rect 14415 4264 14427 4267
rect 14550 4264 14556 4276
rect 14415 4236 14556 4264
rect 14415 4233 14427 4236
rect 14369 4227 14427 4233
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 14734 4264 14740 4276
rect 14695 4236 14740 4264
rect 14734 4224 14740 4236
rect 14792 4224 14798 4276
rect 17402 4264 17408 4276
rect 17363 4236 17408 4264
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 21634 4264 21640 4276
rect 21547 4236 21640 4264
rect 21634 4224 21640 4236
rect 21692 4264 21698 4276
rect 22005 4267 22063 4273
rect 22005 4264 22017 4267
rect 21692 4236 22017 4264
rect 21692 4224 21698 4236
rect 22005 4233 22017 4236
rect 22051 4264 22063 4267
rect 22186 4264 22192 4276
rect 22051 4236 22192 4264
rect 22051 4233 22063 4236
rect 22005 4227 22063 4233
rect 22186 4224 22192 4236
rect 22244 4224 22250 4276
rect 22925 4267 22983 4273
rect 22925 4233 22937 4267
rect 22971 4264 22983 4267
rect 23014 4264 23020 4276
rect 22971 4236 23020 4264
rect 22971 4233 22983 4236
rect 22925 4227 22983 4233
rect 23014 4224 23020 4236
rect 23072 4224 23078 4276
rect 23750 4264 23756 4276
rect 23711 4236 23756 4264
rect 23750 4224 23756 4236
rect 23808 4224 23814 4276
rect 3510 4196 3516 4208
rect 2240 4168 3516 4196
rect 2240 4072 2268 4168
rect 3510 4156 3516 4168
rect 3568 4196 3574 4208
rect 3973 4199 4031 4205
rect 3973 4196 3985 4199
rect 3568 4168 3985 4196
rect 3568 4156 3574 4168
rect 3973 4165 3985 4168
rect 4019 4165 4031 4199
rect 8754 4196 8760 4208
rect 8715 4168 8760 4196
rect 3973 4159 4031 4165
rect 8754 4156 8760 4168
rect 8812 4156 8818 4208
rect 10045 4199 10103 4205
rect 10045 4165 10057 4199
rect 10091 4196 10103 4199
rect 10226 4196 10232 4208
rect 10091 4168 10232 4196
rect 10091 4165 10103 4168
rect 10045 4159 10103 4165
rect 10226 4156 10232 4168
rect 10284 4156 10290 4208
rect 10778 4156 10784 4208
rect 10836 4196 10842 4208
rect 14458 4196 14464 4208
rect 10836 4168 11100 4196
rect 10836 4156 10842 4168
rect 2682 4128 2688 4140
rect 2643 4100 2688 4128
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 3602 4088 3608 4140
rect 3660 4128 3666 4140
rect 3878 4128 3884 4140
rect 3660 4100 3884 4128
rect 3660 4088 3666 4100
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 8021 4131 8079 4137
rect 8021 4128 8033 4131
rect 7432 4100 8033 4128
rect 7432 4088 7438 4100
rect 8021 4097 8033 4100
rect 8067 4128 8079 4131
rect 8294 4128 8300 4140
rect 8067 4100 8300 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9585 4131 9643 4137
rect 9585 4128 9597 4131
rect 9456 4100 9597 4128
rect 9456 4088 9462 4100
rect 9585 4097 9597 4100
rect 9631 4097 9643 4131
rect 9585 4091 9643 4097
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 10962 4128 10968 4140
rect 9916 4100 10732 4128
rect 10923 4100 10968 4128
rect 9916 4088 9922 4100
rect 2222 4020 2228 4072
rect 2280 4020 2286 4072
rect 2406 4060 2412 4072
rect 2367 4032 2412 4060
rect 2406 4020 2412 4032
rect 2464 4020 2470 4072
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4029 4123 4063
rect 4065 4023 4123 4029
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 2593 3995 2651 4001
rect 2593 3992 2605 3995
rect 2372 3964 2605 3992
rect 2372 3952 2378 3964
rect 2593 3961 2605 3964
rect 2639 3961 2651 3995
rect 3605 3995 3663 4001
rect 3605 3992 3617 3995
rect 2593 3955 2651 3961
rect 2884 3964 3617 3992
rect 1670 3924 1676 3936
rect 1583 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3924 1734 3936
rect 2038 3924 2044 3936
rect 1728 3896 2044 3924
rect 1728 3884 1734 3896
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2884 3924 2912 3964
rect 3605 3961 3617 3964
rect 3651 3992 3663 3995
rect 3970 3992 3976 4004
rect 3651 3964 3976 3992
rect 3651 3961 3663 3964
rect 3605 3955 3663 3961
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 4080 3936 4108 4023
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4321 4063 4379 4069
rect 4321 4060 4333 4063
rect 4212 4032 4333 4060
rect 4212 4020 4218 4032
rect 4321 4029 4333 4032
rect 4367 4029 4379 4063
rect 5994 4060 6000 4072
rect 5955 4032 6000 4060
rect 4321 4023 4379 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 7282 4060 7288 4072
rect 6972 4032 7288 4060
rect 6972 4020 6978 4032
rect 7282 4020 7288 4032
rect 7340 4060 7346 4072
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 7340 4032 7665 4060
rect 7340 4020 7346 4032
rect 7653 4029 7665 4032
rect 7699 4029 7711 4063
rect 9306 4060 9312 4072
rect 9267 4032 9312 4060
rect 7653 4023 7711 4029
rect 9306 4020 9312 4032
rect 9364 4060 9370 4072
rect 10579 4063 10637 4069
rect 10579 4060 10591 4063
rect 9364 4032 10591 4060
rect 9364 4020 9370 4032
rect 10579 4029 10591 4032
rect 10625 4029 10637 4063
rect 10704 4060 10732 4100
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11072 4128 11100 4168
rect 13648 4168 14464 4196
rect 11149 4131 11207 4137
rect 11149 4128 11161 4131
rect 11072 4100 11161 4128
rect 11149 4097 11161 4100
rect 11195 4097 11207 4131
rect 11149 4091 11207 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4128 11851 4131
rect 12250 4128 12256 4140
rect 11839 4100 12256 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 12250 4088 12256 4100
rect 12308 4088 12314 4140
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13648 4128 13676 4168
rect 14458 4156 14464 4168
rect 14516 4156 14522 4208
rect 13814 4128 13820 4140
rect 13311 4100 13676 4128
rect 13775 4100 13820 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 13998 4128 14004 4140
rect 13959 4100 14004 4128
rect 13998 4088 14004 4100
rect 14056 4128 14062 4140
rect 17420 4128 17448 4224
rect 22830 4156 22836 4208
rect 22888 4196 22894 4208
rect 23201 4199 23259 4205
rect 23201 4196 23213 4199
rect 22888 4168 23213 4196
rect 22888 4156 22894 4168
rect 23201 4165 23213 4168
rect 23247 4165 23259 4199
rect 23201 4159 23259 4165
rect 24118 4156 24124 4208
rect 24176 4196 24182 4208
rect 24176 4168 24808 4196
rect 24176 4156 24182 4168
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 14056 4100 15056 4128
rect 17420 4100 18184 4128
rect 14056 4088 14062 4100
rect 10704 4032 14228 4060
rect 10579 4023 10637 4029
rect 7377 3995 7435 4001
rect 7377 3961 7389 3995
rect 7423 3992 7435 3995
rect 7742 3992 7748 4004
rect 7423 3964 7748 3992
rect 7423 3961 7435 3964
rect 7377 3955 7435 3961
rect 7742 3952 7748 3964
rect 7800 3952 7806 4004
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 9490 3992 9496 4004
rect 8536 3964 9496 3992
rect 8536 3952 8542 3964
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 11882 3992 11888 4004
rect 10100 3964 11888 3992
rect 10100 3952 10106 3964
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 13909 3995 13967 4001
rect 13909 3961 13921 3995
rect 13955 3992 13967 3995
rect 14090 3992 14096 4004
rect 13955 3964 14096 3992
rect 13955 3961 13967 3964
rect 13909 3955 13967 3961
rect 14090 3952 14096 3964
rect 14148 3952 14154 4004
rect 14200 3992 14228 4032
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 14921 4063 14979 4069
rect 14921 4060 14933 4063
rect 14792 4032 14933 4060
rect 14792 4020 14798 4032
rect 14921 4029 14933 4032
rect 14967 4029 14979 4063
rect 15028 4060 15056 4100
rect 15177 4063 15235 4069
rect 15177 4060 15189 4063
rect 15028 4032 15189 4060
rect 14921 4023 14979 4029
rect 15177 4029 15189 4032
rect 15223 4060 15235 4063
rect 16298 4060 16304 4072
rect 15223 4032 16304 4060
rect 15223 4029 15235 4032
rect 15177 4023 15235 4029
rect 16298 4020 16304 4032
rect 16356 4060 16362 4072
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 16356 4032 16865 4060
rect 16356 4020 16362 4032
rect 16853 4029 16865 4032
rect 16899 4029 16911 4063
rect 16853 4023 16911 4029
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4060 17923 4063
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17911 4032 18061 4060
rect 17911 4029 17923 4032
rect 17865 4023 17923 4029
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18156 4060 18184 4100
rect 19904 4100 20269 4128
rect 18305 4063 18363 4069
rect 18305 4060 18317 4063
rect 18156 4032 18317 4060
rect 18049 4023 18107 4029
rect 18305 4029 18317 4032
rect 18351 4029 18363 4063
rect 18305 4023 18363 4029
rect 18064 3992 18092 4023
rect 18138 3992 18144 4004
rect 14200 3964 17908 3992
rect 18064 3964 18144 3992
rect 17880 3936 17908 3964
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 19904 3992 19932 4100
rect 20257 4097 20269 4100
rect 20303 4128 20315 4131
rect 20349 4131 20407 4137
rect 20349 4128 20361 4131
rect 20303 4100 20361 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 20349 4097 20361 4100
rect 20395 4097 20407 4131
rect 22278 4128 22284 4140
rect 22239 4100 22284 4128
rect 20349 4091 20407 4097
rect 22278 4088 22284 4100
rect 22336 4088 22342 4140
rect 24780 4128 24808 4168
rect 25777 4131 25835 4137
rect 25777 4128 25789 4131
rect 24780 4100 25789 4128
rect 25777 4097 25789 4100
rect 25823 4097 25835 4131
rect 25777 4091 25835 4097
rect 21177 4063 21235 4069
rect 21177 4060 21189 4063
rect 18248 3964 19932 3992
rect 19996 4032 21189 4060
rect 18248 3936 18276 3964
rect 19996 3936 20024 4032
rect 21177 4029 21189 4032
rect 21223 4060 21235 4063
rect 21542 4060 21548 4072
rect 21223 4032 21548 4060
rect 21223 4029 21235 4032
rect 21177 4023 21235 4029
rect 21542 4020 21548 4032
rect 21600 4020 21606 4072
rect 22097 4063 22155 4069
rect 22097 4029 22109 4063
rect 22143 4060 22155 4063
rect 22370 4060 22376 4072
rect 22143 4032 22376 4060
rect 22143 4029 22155 4032
rect 22097 4023 22155 4029
rect 22370 4020 22376 4032
rect 22428 4060 22434 4072
rect 23382 4060 23388 4072
rect 22428 4032 23388 4060
rect 22428 4020 22434 4032
rect 23382 4020 23388 4032
rect 23440 4020 23446 4072
rect 23750 4020 23756 4072
rect 23808 4060 23814 4072
rect 24029 4063 24087 4069
rect 24029 4060 24041 4063
rect 23808 4032 24041 4060
rect 23808 4020 23814 4032
rect 24029 4029 24041 4032
rect 24075 4060 24087 4063
rect 24578 4060 24584 4072
rect 24075 4032 24584 4060
rect 24075 4029 24087 4032
rect 24029 4023 24087 4029
rect 24578 4020 24584 4032
rect 24636 4020 24642 4072
rect 25130 4060 25136 4072
rect 25091 4032 25136 4060
rect 25130 4020 25136 4032
rect 25188 4020 25194 4072
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 25406 4060 25412 4072
rect 25271 4032 25412 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25406 4020 25412 4032
rect 25464 4020 25470 4072
rect 20162 3952 20168 4004
rect 20220 3992 20226 4004
rect 20607 3995 20665 4001
rect 20607 3992 20619 3995
rect 20220 3964 20619 3992
rect 20220 3952 20226 3964
rect 20607 3961 20619 3964
rect 20653 3961 20665 3995
rect 20898 3992 20904 4004
rect 20859 3964 20904 3992
rect 20607 3955 20665 3961
rect 20898 3952 20904 3964
rect 20956 3952 20962 4004
rect 22738 3952 22744 4004
rect 22796 3992 22802 4004
rect 24210 3992 24216 4004
rect 22796 3964 24216 3992
rect 22796 3952 22802 3964
rect 24210 3952 24216 3964
rect 24268 3952 24274 4004
rect 24302 3952 24308 4004
rect 24360 3992 24366 4004
rect 25498 3992 25504 4004
rect 24360 3964 25504 3992
rect 24360 3952 24366 3964
rect 25498 3952 25504 3964
rect 25556 3952 25562 4004
rect 2832 3896 2912 3924
rect 2832 3884 2838 3896
rect 3234 3884 3240 3936
rect 3292 3924 3298 3936
rect 4062 3924 4068 3936
rect 3292 3896 4068 3924
rect 3292 3884 3298 3896
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 7561 3927 7619 3933
rect 7561 3924 7573 3927
rect 6696 3896 7573 3924
rect 6696 3884 6702 3896
rect 7561 3893 7573 3896
rect 7607 3924 7619 3927
rect 7926 3924 7932 3936
rect 7607 3896 7932 3924
rect 7607 3893 7619 3896
rect 7561 3887 7619 3893
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 10413 3927 10471 3933
rect 10413 3893 10425 3927
rect 10459 3924 10471 3927
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10459 3896 11069 3924
rect 10459 3893 10471 3896
rect 10413 3887 10471 3893
rect 11057 3893 11069 3896
rect 11103 3924 11115 3927
rect 11330 3924 11336 3936
rect 11103 3896 11336 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 15286 3884 15292 3936
rect 15344 3924 15350 3936
rect 15930 3924 15936 3936
rect 15344 3896 15936 3924
rect 15344 3884 15350 3896
rect 15930 3884 15936 3896
rect 15988 3924 15994 3936
rect 16301 3927 16359 3933
rect 16301 3924 16313 3927
rect 15988 3896 16313 3924
rect 15988 3884 15994 3896
rect 16301 3893 16313 3896
rect 16347 3893 16359 3927
rect 16301 3887 16359 3893
rect 17862 3884 17868 3936
rect 17920 3884 17926 3936
rect 18230 3884 18236 3936
rect 18288 3884 18294 3936
rect 18690 3884 18696 3936
rect 18748 3924 18754 3936
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 18748 3896 19441 3924
rect 18748 3884 18754 3896
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 19978 3924 19984 3936
rect 19939 3896 19984 3924
rect 19429 3887 19487 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20257 3927 20315 3933
rect 20257 3893 20269 3927
rect 20303 3924 20315 3927
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20303 3896 21097 3924
rect 20303 3893 20315 3896
rect 20257 3887 20315 3893
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 22002 3884 22008 3936
rect 22060 3924 22066 3936
rect 22554 3924 22560 3936
rect 22060 3896 22560 3924
rect 22060 3884 22066 3896
rect 22554 3884 22560 3896
rect 22612 3924 22618 3936
rect 23382 3924 23388 3936
rect 22612 3896 23388 3924
rect 22612 3884 22618 3896
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 24670 3924 24676 3936
rect 24631 3896 24676 3924
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 25130 3884 25136 3936
rect 25188 3924 25194 3936
rect 25409 3927 25467 3933
rect 25409 3924 25421 3927
rect 25188 3896 25421 3924
rect 25188 3884 25194 3896
rect 25409 3893 25421 3896
rect 25455 3893 25467 3927
rect 25409 3887 25467 3893
rect 26237 3927 26295 3933
rect 26237 3893 26249 3927
rect 26283 3924 26295 3927
rect 26418 3924 26424 3936
rect 26283 3896 26424 3924
rect 26283 3893 26295 3896
rect 26237 3887 26295 3893
rect 26418 3884 26424 3896
rect 26476 3884 26482 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 5442 3720 5448 3732
rect 4212 3692 5448 3720
rect 4212 3680 4218 3692
rect 5442 3680 5448 3692
rect 5500 3720 5506 3732
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 5500 3692 5641 3720
rect 5500 3680 5506 3692
rect 5629 3689 5641 3692
rect 5675 3689 5687 3723
rect 6270 3720 6276 3732
rect 6231 3692 6276 3720
rect 5629 3683 5687 3689
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 10597 3723 10655 3729
rect 10597 3689 10609 3723
rect 10643 3720 10655 3723
rect 10962 3720 10968 3732
rect 10643 3692 10968 3720
rect 10643 3689 10655 3692
rect 10597 3683 10655 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 13449 3723 13507 3729
rect 13449 3720 13461 3723
rect 13044 3692 13461 3720
rect 13044 3680 13050 3692
rect 13449 3689 13461 3692
rect 13495 3720 13507 3723
rect 14921 3723 14979 3729
rect 14921 3720 14933 3723
rect 13495 3692 14933 3720
rect 13495 3689 13507 3692
rect 13449 3683 13507 3689
rect 14921 3689 14933 3692
rect 14967 3720 14979 3723
rect 15378 3720 15384 3732
rect 14967 3692 15384 3720
rect 14967 3689 14979 3692
rect 14921 3683 14979 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15838 3720 15844 3732
rect 15799 3692 15844 3720
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 17126 3720 17132 3732
rect 17087 3692 17132 3720
rect 17126 3680 17132 3692
rect 17184 3680 17190 3732
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 17497 3723 17555 3729
rect 17497 3720 17509 3723
rect 17460 3692 17509 3720
rect 17460 3680 17466 3692
rect 17497 3689 17509 3692
rect 17543 3720 17555 3723
rect 18690 3720 18696 3732
rect 17543 3692 18368 3720
rect 18651 3692 18696 3720
rect 17543 3689 17555 3692
rect 17497 3683 17555 3689
rect 1670 3652 1676 3664
rect 1583 3624 1676 3652
rect 1670 3612 1676 3624
rect 1728 3652 1734 3664
rect 2866 3652 2872 3664
rect 1728 3624 2872 3652
rect 1728 3612 1734 3624
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 4522 3661 4528 3664
rect 2961 3655 3019 3661
rect 2961 3621 2973 3655
rect 3007 3652 3019 3655
rect 3237 3655 3295 3661
rect 3237 3652 3249 3655
rect 3007 3624 3249 3652
rect 3007 3621 3019 3624
rect 2961 3615 3019 3621
rect 3237 3621 3249 3624
rect 3283 3621 3295 3655
rect 3237 3615 3295 3621
rect 3789 3655 3847 3661
rect 3789 3621 3801 3655
rect 3835 3652 3847 3655
rect 4516 3652 4528 3661
rect 3835 3624 4528 3652
rect 3835 3621 3847 3624
rect 3789 3615 3847 3621
rect 4516 3615 4528 3624
rect 4522 3612 4528 3615
rect 4580 3612 4586 3664
rect 14093 3655 14151 3661
rect 14093 3621 14105 3655
rect 14139 3621 14151 3655
rect 15654 3652 15660 3664
rect 15615 3624 15660 3652
rect 14093 3615 14151 3621
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3584 2835 3587
rect 3878 3584 3884 3596
rect 2823 3556 3884 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 3878 3544 3884 3556
rect 3936 3544 3942 3596
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 4120 3556 4261 3584
rect 4120 3544 4126 3556
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4890 3584 4896 3596
rect 4249 3547 4307 3553
rect 4336 3556 4896 3584
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3326 3516 3332 3528
rect 3283 3488 3332 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 2498 3448 2504 3460
rect 2459 3420 2504 3448
rect 2498 3408 2504 3420
rect 2556 3408 2562 3460
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2096 3352 2237 3380
rect 2096 3340 2102 3352
rect 2225 3349 2237 3352
rect 2271 3380 2283 3383
rect 3068 3380 3096 3479
rect 3326 3476 3332 3488
rect 3384 3516 3390 3528
rect 4336 3516 4364 3556
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 7009 3587 7067 3593
rect 7009 3553 7021 3587
rect 7055 3584 7067 3587
rect 7098 3584 7104 3596
rect 7055 3556 7104 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 7282 3593 7288 3596
rect 7276 3584 7288 3593
rect 7243 3556 7288 3584
rect 7276 3547 7288 3556
rect 7282 3544 7288 3547
rect 7340 3544 7346 3596
rect 9766 3584 9772 3596
rect 9727 3556 9772 3584
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3584 10839 3587
rect 11313 3587 11371 3593
rect 11313 3584 11325 3587
rect 10827 3556 11325 3584
rect 10827 3553 10839 3556
rect 10781 3547 10839 3553
rect 11313 3553 11325 3556
rect 11359 3584 11371 3587
rect 11606 3584 11612 3596
rect 11359 3556 11612 3584
rect 11359 3553 11371 3556
rect 11313 3547 11371 3553
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 14108 3584 14136 3615
rect 15654 3612 15660 3624
rect 15712 3612 15718 3664
rect 15930 3652 15936 3664
rect 15891 3624 15936 3652
rect 15930 3612 15936 3624
rect 15988 3612 15994 3664
rect 17218 3612 17224 3664
rect 17276 3652 17282 3664
rect 18049 3655 18107 3661
rect 18049 3652 18061 3655
rect 17276 3624 18061 3652
rect 17276 3612 17282 3624
rect 18049 3621 18061 3624
rect 18095 3621 18107 3655
rect 18230 3652 18236 3664
rect 18191 3624 18236 3652
rect 18049 3615 18107 3621
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 18340 3661 18368 3692
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19484 3692 19809 3720
rect 19484 3680 19490 3692
rect 19797 3689 19809 3692
rect 19843 3689 19855 3723
rect 19797 3683 19855 3689
rect 20717 3723 20775 3729
rect 20717 3689 20729 3723
rect 20763 3720 20775 3723
rect 20806 3720 20812 3732
rect 20763 3692 20812 3720
rect 20763 3689 20775 3692
rect 20717 3683 20775 3689
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 21082 3680 21088 3732
rect 21140 3720 21146 3732
rect 21634 3720 21640 3732
rect 21140 3692 21640 3720
rect 21140 3680 21146 3692
rect 21634 3680 21640 3692
rect 21692 3720 21698 3732
rect 21913 3723 21971 3729
rect 21913 3720 21925 3723
rect 21692 3692 21925 3720
rect 21692 3680 21698 3692
rect 21913 3689 21925 3692
rect 21959 3689 21971 3723
rect 22370 3720 22376 3732
rect 22331 3692 22376 3720
rect 21913 3683 21971 3689
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 22646 3680 22652 3732
rect 22704 3720 22710 3732
rect 23017 3723 23075 3729
rect 23017 3720 23029 3723
rect 22704 3692 23029 3720
rect 22704 3680 22710 3692
rect 23017 3689 23029 3692
rect 23063 3689 23075 3723
rect 23017 3683 23075 3689
rect 23753 3723 23811 3729
rect 23753 3689 23765 3723
rect 23799 3720 23811 3723
rect 24302 3720 24308 3732
rect 23799 3692 24308 3720
rect 23799 3689 23811 3692
rect 23753 3683 23811 3689
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 25409 3723 25467 3729
rect 25409 3720 25421 3723
rect 24412 3692 25421 3720
rect 18325 3655 18383 3661
rect 18325 3621 18337 3655
rect 18371 3621 18383 3655
rect 20824 3652 20852 3680
rect 21453 3655 21511 3661
rect 21453 3652 21465 3655
rect 20824 3624 21465 3652
rect 18325 3615 18383 3621
rect 21453 3621 21465 3624
rect 21499 3621 21511 3655
rect 21453 3615 21511 3621
rect 21542 3612 21548 3664
rect 21600 3652 21606 3664
rect 21600 3624 21645 3652
rect 21600 3612 21606 3624
rect 23382 3612 23388 3664
rect 23440 3652 23446 3664
rect 24412 3652 24440 3692
rect 25409 3689 25421 3692
rect 25455 3689 25467 3723
rect 26234 3720 26240 3732
rect 26195 3692 26240 3720
rect 25409 3683 25467 3689
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 23440 3624 24440 3652
rect 24581 3655 24639 3661
rect 23440 3612 23446 3624
rect 24581 3621 24593 3655
rect 24627 3652 24639 3655
rect 26326 3652 26332 3664
rect 24627 3624 26332 3652
rect 24627 3621 24639 3624
rect 24581 3615 24639 3621
rect 26326 3612 26332 3624
rect 26384 3612 26390 3664
rect 14642 3584 14648 3596
rect 14108 3556 14648 3584
rect 14642 3544 14648 3556
rect 14700 3544 14706 3596
rect 16850 3584 16856 3596
rect 16763 3556 16856 3584
rect 16850 3544 16856 3556
rect 16908 3584 16914 3596
rect 19613 3587 19671 3593
rect 19613 3584 19625 3587
rect 16908 3556 19625 3584
rect 16908 3544 16914 3556
rect 19613 3553 19625 3556
rect 19659 3553 19671 3587
rect 19613 3547 19671 3553
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 21269 3587 21327 3593
rect 21269 3584 21281 3587
rect 20680 3556 21281 3584
rect 20680 3544 20686 3556
rect 21269 3553 21281 3556
rect 21315 3553 21327 3587
rect 21269 3547 21327 3553
rect 22462 3544 22468 3596
rect 22520 3584 22526 3596
rect 23109 3587 23167 3593
rect 23109 3584 23121 3587
rect 22520 3556 23121 3584
rect 22520 3544 22526 3556
rect 23109 3553 23121 3556
rect 23155 3553 23167 3587
rect 23109 3547 23167 3553
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 25777 3587 25835 3593
rect 25777 3584 25789 3587
rect 24268 3556 25789 3584
rect 24268 3544 24274 3556
rect 25777 3553 25789 3556
rect 25823 3553 25835 3587
rect 25777 3547 25835 3553
rect 3384 3488 4364 3516
rect 10045 3519 10103 3525
rect 3384 3476 3390 3488
rect 10045 3485 10057 3519
rect 10091 3516 10103 3519
rect 10962 3516 10968 3528
rect 10091 3488 10968 3516
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 13081 3519 13139 3525
rect 11112 3488 11157 3516
rect 11112 3476 11118 3488
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 14090 3516 14096 3528
rect 13127 3488 14096 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 14185 3519 14243 3525
rect 14185 3485 14197 3519
rect 14231 3516 14243 3519
rect 14366 3516 14372 3528
rect 14231 3488 14372 3516
rect 14231 3485 14243 3488
rect 14185 3479 14243 3485
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 19886 3516 19892 3528
rect 19847 3488 19892 3516
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 20349 3519 20407 3525
rect 20349 3485 20361 3519
rect 20395 3516 20407 3519
rect 21542 3516 21548 3528
rect 20395 3488 21548 3516
rect 20395 3485 20407 3488
rect 20349 3479 20407 3485
rect 21542 3476 21548 3488
rect 21600 3476 21606 3528
rect 23014 3516 23020 3528
rect 22975 3488 23020 3516
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3485 24731 3519
rect 25038 3516 25044 3528
rect 24999 3488 25044 3516
rect 24673 3479 24731 3485
rect 9490 3408 9496 3460
rect 9548 3448 9554 3460
rect 10781 3451 10839 3457
rect 10781 3448 10793 3451
rect 9548 3420 10793 3448
rect 9548 3408 9554 3420
rect 10781 3417 10793 3420
rect 10827 3448 10839 3451
rect 10873 3451 10931 3457
rect 10873 3448 10885 3451
rect 10827 3420 10885 3448
rect 10827 3417 10839 3420
rect 10781 3411 10839 3417
rect 10873 3417 10885 3420
rect 10919 3417 10931 3451
rect 13630 3448 13636 3460
rect 13591 3420 13636 3448
rect 10873 3411 10931 3417
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 15381 3451 15439 3457
rect 15381 3417 15393 3451
rect 15427 3448 15439 3451
rect 16574 3448 16580 3460
rect 15427 3420 16580 3448
rect 15427 3417 15439 3420
rect 15381 3411 15439 3417
rect 16574 3408 16580 3420
rect 16632 3408 16638 3460
rect 17770 3448 17776 3460
rect 17731 3420 17776 3448
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 19334 3448 19340 3460
rect 19295 3420 19340 3448
rect 19334 3408 19340 3420
rect 19392 3408 19398 3460
rect 20993 3451 21051 3457
rect 20993 3417 21005 3451
rect 21039 3448 21051 3451
rect 21174 3448 21180 3460
rect 21039 3420 21180 3448
rect 21039 3417 21051 3420
rect 20993 3411 21051 3417
rect 21174 3408 21180 3420
rect 21232 3408 21238 3460
rect 22370 3408 22376 3460
rect 22428 3448 22434 3460
rect 22922 3448 22928 3460
rect 22428 3420 22928 3448
rect 22428 3408 22434 3420
rect 22922 3408 22928 3420
rect 22980 3408 22986 3460
rect 24026 3408 24032 3460
rect 24084 3448 24090 3460
rect 24121 3451 24179 3457
rect 24121 3448 24133 3451
rect 24084 3420 24133 3448
rect 24084 3408 24090 3420
rect 24121 3417 24133 3420
rect 24167 3417 24179 3451
rect 24121 3411 24179 3417
rect 24302 3408 24308 3460
rect 24360 3448 24366 3460
rect 24688 3448 24716 3479
rect 25038 3476 25044 3488
rect 25096 3476 25102 3528
rect 24360 3420 24716 3448
rect 24360 3408 24366 3420
rect 3510 3380 3516 3392
rect 2271 3352 3096 3380
rect 3471 3352 3516 3380
rect 2271 3349 2283 3352
rect 2225 3343 2283 3349
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 6914 3380 6920 3392
rect 6875 3352 6920 3380
rect 6914 3340 6920 3352
rect 6972 3380 6978 3392
rect 8389 3383 8447 3389
rect 8389 3380 8401 3383
rect 6972 3352 8401 3380
rect 6972 3340 6978 3352
rect 8389 3349 8401 3352
rect 8435 3349 8447 3383
rect 9306 3380 9312 3392
rect 9267 3352 9312 3380
rect 8389 3343 8447 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 12492 3352 12537 3380
rect 12492 3340 12498 3352
rect 15286 3340 15292 3392
rect 15344 3380 15350 3392
rect 16482 3380 16488 3392
rect 15344 3352 16488 3380
rect 15344 3340 15350 3352
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 19058 3380 19064 3392
rect 19019 3352 19064 3380
rect 19058 3340 19064 3352
rect 19116 3340 19122 3392
rect 22554 3380 22560 3392
rect 22515 3352 22560 3380
rect 22554 3340 22560 3352
rect 22612 3340 22618 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1489 3179 1547 3185
rect 1489 3145 1501 3179
rect 1535 3176 1547 3179
rect 1762 3176 1768 3188
rect 1535 3148 1768 3176
rect 1535 3145 1547 3148
rect 1489 3139 1547 3145
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 3326 3176 3332 3188
rect 2915 3148 3332 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 3878 3176 3884 3188
rect 3835 3148 3884 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4062 3176 4068 3188
rect 4023 3148 4068 3176
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 4580 3148 5641 3176
rect 4580 3136 4586 3148
rect 5629 3145 5641 3148
rect 5675 3145 5687 3179
rect 5629 3139 5687 3145
rect 6273 3179 6331 3185
rect 6273 3145 6285 3179
rect 6319 3176 6331 3179
rect 6362 3176 6368 3188
rect 6319 3148 6368 3176
rect 6319 3145 6331 3148
rect 6273 3139 6331 3145
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 6917 3179 6975 3185
rect 6917 3145 6929 3179
rect 6963 3176 6975 3179
rect 7006 3176 7012 3188
rect 6963 3148 7012 3176
rect 6963 3145 6975 3148
rect 6917 3139 6975 3145
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7156 3148 7849 3176
rect 7156 3136 7162 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 7837 3139 7895 3145
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 8478 3176 8484 3188
rect 8435 3148 8484 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 3050 3068 3056 3120
rect 3108 3108 3114 3120
rect 3418 3108 3424 3120
rect 3108 3080 3424 3108
rect 3108 3068 3114 3080
rect 3418 3068 3424 3080
rect 3476 3068 3482 3120
rect 1762 3000 1768 3052
rect 1820 3040 1826 3052
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1820 3012 1961 3040
rect 1820 3000 1826 3012
rect 1949 3009 1961 3012
rect 1995 3040 2007 3043
rect 2498 3040 2504 3052
rect 1995 3012 2504 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 3234 3040 3240 3052
rect 3195 3012 3240 3040
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 4080 3040 4108 3136
rect 7852 3108 7880 3139
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 9582 3176 9588 3188
rect 8803 3148 9588 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 14366 3176 14372 3188
rect 11480 3148 14372 3176
rect 11480 3136 11486 3148
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 14734 3176 14740 3188
rect 14695 3148 14740 3176
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 15930 3136 15936 3188
rect 15988 3176 15994 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 15988 3148 16865 3176
rect 15988 3136 15994 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 17276 3148 17325 3176
rect 17276 3136 17282 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 17678 3176 17684 3188
rect 17639 3148 17684 3176
rect 17313 3139 17371 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 18138 3176 18144 3188
rect 18099 3148 18144 3176
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 22557 3179 22615 3185
rect 22557 3145 22569 3179
rect 22603 3176 22615 3179
rect 22646 3176 22652 3188
rect 22603 3148 22652 3176
rect 22603 3145 22615 3148
rect 22557 3139 22615 3145
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 23014 3136 23020 3188
rect 23072 3176 23078 3188
rect 23198 3176 23204 3188
rect 23072 3148 23204 3176
rect 23072 3136 23078 3148
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 24210 3136 24216 3188
rect 24268 3176 24274 3188
rect 24673 3179 24731 3185
rect 24673 3176 24685 3179
rect 24268 3148 24685 3176
rect 24268 3136 24274 3148
rect 24673 3145 24685 3148
rect 24719 3145 24731 3179
rect 26326 3176 26332 3188
rect 26287 3148 26332 3176
rect 24673 3139 24731 3145
rect 26326 3136 26332 3148
rect 26384 3136 26390 3188
rect 9033 3111 9091 3117
rect 9033 3108 9045 3111
rect 7852 3080 9045 3108
rect 9033 3077 9045 3080
rect 9079 3108 9091 3111
rect 9079 3080 9260 3108
rect 9079 3077 9091 3080
rect 9033 3071 9091 3077
rect 9232 3052 9260 3080
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 4080 3012 4261 3040
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 2958 2972 2964 2984
rect 2919 2944 2964 2972
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 4264 2972 4292 3003
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 7064 3012 7481 3040
rect 7064 3000 7070 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 9214 3040 9220 3052
rect 9127 3012 9220 3040
rect 7469 3003 7527 3009
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 14550 3040 14556 3052
rect 14424 3012 14556 3040
rect 14424 3000 14430 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14752 3040 14780 3136
rect 16298 3108 16304 3120
rect 16259 3080 16304 3108
rect 16298 3068 16304 3080
rect 16356 3068 16362 3120
rect 19334 3068 19340 3120
rect 19392 3108 19398 3120
rect 19705 3111 19763 3117
rect 19705 3108 19717 3111
rect 19392 3080 19717 3108
rect 19392 3068 19398 3080
rect 19705 3077 19717 3080
rect 19751 3077 19763 3111
rect 19705 3071 19763 3077
rect 20070 3068 20076 3120
rect 20128 3108 20134 3120
rect 21269 3111 21327 3117
rect 21269 3108 21281 3111
rect 20128 3080 21281 3108
rect 20128 3068 20134 3080
rect 21269 3077 21281 3080
rect 21315 3077 21327 3111
rect 21269 3071 21327 3077
rect 21542 3068 21548 3120
rect 21600 3108 21606 3120
rect 23750 3108 23756 3120
rect 21600 3080 21864 3108
rect 23711 3080 23756 3108
rect 21600 3068 21606 3080
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14752 3012 14933 3040
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 18012 3012 18613 3040
rect 18012 3000 18018 3012
rect 18601 3009 18613 3012
rect 18647 3040 18659 3043
rect 18690 3040 18696 3052
rect 18647 3012 18696 3040
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 18690 3000 18696 3012
rect 18748 3000 18754 3052
rect 20162 3040 20168 3052
rect 20123 3012 20168 3040
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 21634 3040 21640 3052
rect 21595 3012 21640 3040
rect 21634 3000 21640 3012
rect 21692 3000 21698 3052
rect 21836 3049 21864 3080
rect 23750 3068 23756 3080
rect 23808 3068 23814 3120
rect 24854 3108 24860 3120
rect 24228 3080 24860 3108
rect 24228 3049 24256 3080
rect 24854 3068 24860 3080
rect 24912 3068 24918 3120
rect 21821 3043 21879 3049
rect 21821 3009 21833 3043
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 24213 3043 24271 3049
rect 24213 3009 24225 3043
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 24305 3043 24363 3049
rect 24305 3009 24317 3043
rect 24351 3040 24363 3043
rect 24946 3040 24952 3052
rect 24351 3012 24952 3040
rect 24351 3009 24363 3012
rect 24305 3003 24363 3009
rect 24946 3000 24952 3012
rect 25004 3040 25010 3052
rect 25041 3043 25099 3049
rect 25041 3040 25053 3043
rect 25004 3012 25053 3040
rect 25004 3000 25010 3012
rect 25041 3009 25053 3012
rect 25087 3009 25099 3043
rect 25406 3040 25412 3052
rect 25367 3012 25412 3040
rect 25041 3003 25099 3009
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 5074 2972 5080 2984
rect 4264 2944 5080 2972
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 7282 2972 7288 2984
rect 6687 2944 7288 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 7282 2932 7288 2944
rect 7340 2972 7346 2984
rect 8202 2972 8208 2984
rect 7340 2944 8208 2972
rect 7340 2932 7346 2944
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9490 2981 9496 2984
rect 9473 2975 9496 2981
rect 9473 2972 9485 2975
rect 9364 2944 9485 2972
rect 9364 2932 9370 2944
rect 9473 2941 9485 2944
rect 9548 2972 9554 2984
rect 12069 2975 12127 2981
rect 9548 2944 9621 2972
rect 9473 2935 9496 2941
rect 9490 2932 9496 2935
rect 9548 2932 9554 2944
rect 12069 2941 12081 2975
rect 12115 2972 12127 2975
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12115 2944 12449 2972
rect 12115 2941 12127 2944
rect 12069 2935 12127 2941
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12704 2975 12762 2981
rect 12704 2972 12716 2975
rect 12437 2935 12495 2941
rect 12636 2944 12716 2972
rect 2038 2904 2044 2916
rect 1999 2876 2044 2904
rect 2038 2864 2044 2876
rect 2096 2864 2102 2916
rect 3510 2864 3516 2916
rect 3568 2904 3574 2916
rect 4494 2907 4552 2913
rect 4494 2904 4506 2907
rect 3568 2876 4506 2904
rect 3568 2864 3574 2876
rect 4494 2873 4506 2876
rect 4540 2904 4552 2907
rect 5350 2904 5356 2916
rect 4540 2876 5356 2904
rect 4540 2873 4552 2876
rect 4494 2867 4552 2873
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 7193 2907 7251 2913
rect 7193 2873 7205 2907
rect 7239 2904 7251 2907
rect 7742 2904 7748 2916
rect 7239 2876 7748 2904
rect 7239 2873 7251 2876
rect 7193 2867 7251 2873
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 11422 2904 11428 2916
rect 9732 2876 11428 2904
rect 9732 2864 9738 2876
rect 11422 2864 11428 2876
rect 11480 2864 11486 2916
rect 11885 2907 11943 2913
rect 11885 2873 11897 2907
rect 11931 2904 11943 2907
rect 12636 2904 12664 2944
rect 12704 2941 12716 2944
rect 12750 2972 12762 2975
rect 13446 2972 13452 2984
rect 12750 2944 13452 2972
rect 12750 2941 12762 2944
rect 12704 2935 12762 2941
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 19058 2932 19064 2984
rect 19116 2972 19122 2984
rect 19978 2972 19984 2984
rect 19116 2944 19984 2972
rect 19116 2932 19122 2944
rect 19978 2932 19984 2944
rect 20036 2972 20042 2984
rect 20257 2975 20315 2981
rect 20257 2972 20269 2975
rect 20036 2944 20269 2972
rect 20036 2932 20042 2944
rect 20257 2941 20269 2944
rect 20303 2941 20315 2975
rect 22833 2975 22891 2981
rect 22833 2972 22845 2975
rect 20257 2935 20315 2941
rect 21744 2944 22845 2972
rect 21744 2916 21772 2944
rect 22833 2941 22845 2944
rect 22879 2941 22891 2975
rect 25222 2972 25228 2984
rect 25135 2944 25228 2972
rect 22833 2935 22891 2941
rect 25222 2932 25228 2944
rect 25280 2972 25286 2984
rect 25961 2975 26019 2981
rect 25961 2972 25973 2975
rect 25280 2944 25973 2972
rect 25280 2932 25286 2944
rect 25961 2941 25973 2944
rect 26007 2941 26019 2975
rect 25961 2935 26019 2941
rect 11931 2876 12664 2904
rect 15188 2907 15246 2913
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 15188 2873 15200 2907
rect 15234 2904 15246 2907
rect 15378 2904 15384 2916
rect 15234 2876 15384 2904
rect 15234 2873 15246 2876
rect 15188 2867 15246 2873
rect 15378 2864 15384 2876
rect 15436 2864 15442 2916
rect 18598 2904 18604 2916
rect 18559 2876 18604 2904
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 18690 2864 18696 2916
rect 18748 2904 18754 2916
rect 19153 2907 19211 2913
rect 19153 2904 19165 2907
rect 18748 2876 19165 2904
rect 18748 2864 18754 2876
rect 19153 2873 19165 2876
rect 19199 2904 19211 2907
rect 19429 2907 19487 2913
rect 19429 2904 19441 2907
rect 19199 2876 19441 2904
rect 19199 2873 19211 2876
rect 19153 2867 19211 2873
rect 19429 2873 19441 2876
rect 19475 2904 19487 2907
rect 19886 2904 19892 2916
rect 19475 2876 19892 2904
rect 19475 2873 19487 2876
rect 19429 2867 19487 2873
rect 19886 2864 19892 2876
rect 19944 2864 19950 2916
rect 20070 2864 20076 2916
rect 20128 2904 20134 2916
rect 20165 2907 20223 2913
rect 20165 2904 20177 2907
rect 20128 2876 20177 2904
rect 20128 2864 20134 2876
rect 20165 2873 20177 2876
rect 20211 2873 20223 2907
rect 20165 2867 20223 2873
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 20901 2907 20959 2913
rect 20901 2904 20913 2907
rect 20680 2876 20913 2904
rect 20680 2864 20686 2876
rect 20901 2873 20913 2876
rect 20947 2873 20959 2907
rect 21726 2904 21732 2916
rect 21687 2876 21732 2904
rect 20901 2867 20959 2873
rect 21726 2864 21732 2876
rect 21784 2864 21790 2916
rect 24213 2907 24271 2913
rect 24213 2873 24225 2907
rect 24259 2904 24271 2907
rect 26142 2904 26148 2916
rect 24259 2876 26148 2904
rect 24259 2873 24271 2876
rect 24213 2867 24271 2873
rect 26142 2864 26148 2876
rect 26200 2864 26206 2916
rect 1210 2796 1216 2848
rect 1268 2836 1274 2848
rect 1670 2836 1676 2848
rect 1268 2808 1676 2836
rect 1268 2796 1274 2808
rect 1670 2796 1676 2808
rect 1728 2836 1734 2848
rect 1949 2839 2007 2845
rect 1949 2836 1961 2839
rect 1728 2808 1961 2836
rect 1728 2796 1734 2808
rect 1949 2805 1961 2808
rect 1995 2805 2007 2839
rect 2498 2836 2504 2848
rect 2459 2808 2504 2836
rect 1949 2799 2007 2805
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 7377 2839 7435 2845
rect 7377 2836 7389 2839
rect 5224 2808 7389 2836
rect 5224 2796 5230 2808
rect 7377 2805 7389 2808
rect 7423 2836 7435 2839
rect 7558 2836 7564 2848
rect 7423 2808 7564 2836
rect 7423 2805 7435 2808
rect 7377 2799 7435 2805
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 10597 2839 10655 2845
rect 10597 2805 10609 2839
rect 10643 2836 10655 2839
rect 10686 2836 10692 2848
rect 10643 2808 10692 2836
rect 10643 2805 10655 2808
rect 10597 2799 10655 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 10870 2796 10876 2848
rect 10928 2836 10934 2848
rect 11054 2836 11060 2848
rect 10928 2808 11060 2836
rect 10928 2796 10934 2808
rect 11054 2796 11060 2808
rect 11112 2836 11118 2848
rect 11149 2839 11207 2845
rect 11149 2836 11161 2839
rect 11112 2808 11161 2836
rect 11112 2796 11118 2808
rect 11149 2805 11161 2808
rect 11195 2836 11207 2839
rect 12069 2839 12127 2845
rect 12069 2836 12081 2839
rect 11195 2808 12081 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 12069 2805 12081 2808
rect 12115 2836 12127 2839
rect 12161 2839 12219 2845
rect 12161 2836 12173 2839
rect 12115 2808 12173 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 12161 2805 12173 2808
rect 12207 2805 12219 2839
rect 13814 2836 13820 2848
rect 13727 2808 13820 2836
rect 12161 2799 12219 2805
rect 13814 2796 13820 2808
rect 13872 2836 13878 2848
rect 14550 2836 14556 2848
rect 13872 2808 14556 2836
rect 13872 2796 13878 2808
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 25590 2836 25596 2848
rect 20036 2808 25596 2836
rect 20036 2796 20042 2808
rect 25590 2796 25596 2808
rect 25648 2796 25654 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 198 2592 204 2644
rect 256 2632 262 2644
rect 1578 2632 1584 2644
rect 256 2604 1584 2632
rect 256 2592 262 2604
rect 1578 2592 1584 2604
rect 1636 2632 1642 2644
rect 1949 2635 2007 2641
rect 1949 2632 1961 2635
rect 1636 2604 1961 2632
rect 1636 2592 1642 2604
rect 1949 2601 1961 2604
rect 1995 2632 2007 2635
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 1995 2604 2421 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2409 2595 2467 2601
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3476 2604 3801 2632
rect 3476 2592 3482 2604
rect 3789 2601 3801 2604
rect 3835 2632 3847 2635
rect 5442 2632 5448 2644
rect 3835 2604 4476 2632
rect 3835 2601 3847 2604
rect 3789 2595 3847 2601
rect 2038 2564 2044 2576
rect 1999 2536 2044 2564
rect 2038 2524 2044 2536
rect 2096 2524 2102 2576
rect 4448 2573 4476 2604
rect 4724 2604 5448 2632
rect 4724 2573 4752 2604
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 9214 2592 9220 2644
rect 9272 2632 9278 2644
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 9272 2604 9597 2632
rect 9272 2592 9278 2604
rect 9585 2601 9597 2604
rect 9631 2632 9643 2635
rect 10870 2632 10876 2644
rect 9631 2604 10876 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 4433 2567 4491 2573
rect 4433 2533 4445 2567
rect 4479 2533 4491 2567
rect 4433 2527 4491 2533
rect 4617 2567 4675 2573
rect 4617 2533 4629 2567
rect 4663 2533 4675 2567
rect 4617 2527 4675 2533
rect 4709 2567 4767 2573
rect 4709 2533 4721 2567
rect 4755 2533 4767 2567
rect 5074 2564 5080 2576
rect 5035 2536 5080 2564
rect 4709 2527 4767 2533
rect 658 2456 664 2508
rect 716 2496 722 2508
rect 1765 2499 1823 2505
rect 1765 2496 1777 2499
rect 716 2468 1777 2496
rect 716 2456 722 2468
rect 1765 2465 1777 2468
rect 1811 2496 1823 2499
rect 2869 2499 2927 2505
rect 2869 2496 2881 2499
rect 1811 2468 2881 2496
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 2869 2465 2881 2468
rect 2915 2496 2927 2499
rect 3418 2496 3424 2508
rect 2915 2468 3424 2496
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 3513 2499 3571 2505
rect 3513 2465 3525 2499
rect 3559 2496 3571 2499
rect 3786 2496 3792 2508
rect 3559 2468 3792 2496
rect 3559 2465 3571 2468
rect 3513 2459 3571 2465
rect 3786 2456 3792 2468
rect 3844 2496 3850 2508
rect 4632 2496 4660 2527
rect 5074 2524 5080 2536
rect 5132 2564 5138 2576
rect 6641 2567 6699 2573
rect 6641 2564 6653 2567
rect 5132 2536 6653 2564
rect 5132 2524 5138 2536
rect 6641 2533 6653 2536
rect 6687 2564 6699 2567
rect 6687 2536 7236 2564
rect 6687 2533 6699 2536
rect 6641 2527 6699 2533
rect 3844 2468 4660 2496
rect 5721 2499 5779 2505
rect 3844 2456 3850 2468
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6362 2496 6368 2508
rect 5767 2468 6368 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 7208 2505 7236 2536
rect 7466 2505 7472 2508
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2465 7251 2499
rect 7460 2496 7472 2505
rect 7193 2459 7251 2465
rect 7300 2468 7472 2496
rect 2958 2428 2964 2440
rect 2919 2400 2964 2428
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 6273 2431 6331 2437
rect 6273 2397 6285 2431
rect 6319 2428 6331 2431
rect 7300 2428 7328 2468
rect 7460 2459 7472 2468
rect 7466 2456 7472 2459
rect 7524 2456 7530 2508
rect 10060 2505 10088 2604
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11422 2632 11428 2644
rect 11383 2604 11428 2632
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 14274 2632 14280 2644
rect 12483 2604 14280 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 14274 2592 14280 2604
rect 14332 2632 14338 2644
rect 16853 2635 16911 2641
rect 16853 2632 16865 2635
rect 14332 2604 16865 2632
rect 14332 2592 14338 2604
rect 13262 2524 13268 2576
rect 13320 2564 13326 2576
rect 14476 2573 14504 2604
rect 16853 2601 16865 2604
rect 16899 2601 16911 2635
rect 16853 2595 16911 2601
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 19797 2635 19855 2641
rect 19797 2632 19809 2635
rect 19576 2604 19809 2632
rect 19576 2592 19582 2604
rect 19797 2601 19809 2604
rect 19843 2601 19855 2635
rect 22462 2632 22468 2644
rect 22423 2604 22468 2632
rect 19797 2595 19855 2601
rect 14369 2567 14427 2573
rect 14369 2564 14381 2567
rect 13320 2536 14381 2564
rect 13320 2524 13326 2536
rect 14369 2533 14381 2536
rect 14415 2533 14427 2567
rect 14369 2527 14427 2533
rect 14461 2567 14519 2573
rect 14461 2533 14473 2567
rect 14507 2533 14519 2567
rect 14461 2527 14519 2533
rect 14734 2524 14740 2576
rect 14792 2564 14798 2576
rect 14829 2567 14887 2573
rect 14829 2564 14841 2567
rect 14792 2536 14841 2564
rect 14792 2524 14798 2536
rect 14829 2533 14841 2536
rect 14875 2533 14887 2567
rect 14829 2527 14887 2533
rect 10318 2505 10324 2508
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2465 10103 2499
rect 10312 2496 10324 2505
rect 10045 2459 10103 2465
rect 10152 2468 10324 2496
rect 6319 2400 7328 2428
rect 9217 2431 9275 2437
rect 6319 2397 6331 2400
rect 6273 2391 6331 2397
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 10152 2428 10180 2468
rect 10312 2459 10324 2468
rect 10318 2456 10324 2459
rect 10376 2456 10382 2508
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11112 2468 11989 2496
rect 11112 2456 11118 2468
rect 11977 2465 11989 2468
rect 12023 2496 12035 2499
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 12023 2468 12725 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 12713 2459 12771 2465
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 9263 2400 10180 2428
rect 13648 2400 14289 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 1489 2363 1547 2369
rect 1489 2329 1501 2363
rect 1535 2360 1547 2363
rect 1854 2360 1860 2372
rect 1535 2332 1860 2360
rect 1535 2329 1547 2332
rect 1489 2323 1547 2329
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 4157 2363 4215 2369
rect 4157 2329 4169 2363
rect 4203 2360 4215 2363
rect 4246 2360 4252 2372
rect 4203 2332 4252 2360
rect 4203 2329 4215 2332
rect 4157 2323 4215 2329
rect 4246 2320 4252 2332
rect 4304 2320 4310 2372
rect 5902 2360 5908 2372
rect 5863 2332 5908 2360
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 13648 2304 13676 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14844 2428 14872 2527
rect 16758 2524 16764 2576
rect 16816 2564 16822 2576
rect 18049 2567 18107 2573
rect 18049 2564 18061 2567
rect 16816 2536 18061 2564
rect 16816 2524 16822 2536
rect 18049 2533 18061 2536
rect 18095 2564 18107 2567
rect 18693 2567 18751 2573
rect 18693 2564 18705 2567
rect 18095 2536 18705 2564
rect 18095 2533 18107 2536
rect 18049 2527 18107 2533
rect 18693 2533 18705 2536
rect 18739 2533 18751 2567
rect 18874 2564 18880 2576
rect 18835 2536 18880 2564
rect 18693 2527 18751 2533
rect 18874 2524 18880 2536
rect 18932 2524 18938 2576
rect 15746 2505 15752 2508
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2496 15347 2499
rect 15740 2496 15752 2505
rect 15335 2468 15752 2496
rect 15335 2465 15347 2468
rect 15289 2459 15347 2465
rect 15740 2459 15752 2468
rect 15746 2456 15752 2459
rect 15804 2456 15810 2508
rect 16666 2456 16672 2508
rect 16724 2496 16730 2508
rect 19521 2499 19579 2505
rect 19521 2496 19533 2499
rect 16724 2468 19533 2496
rect 16724 2456 16730 2468
rect 19521 2465 19533 2468
rect 19567 2496 19579 2499
rect 19812 2496 19840 2595
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 23658 2592 23664 2644
rect 23716 2632 23722 2644
rect 23753 2635 23811 2641
rect 23753 2632 23765 2635
rect 23716 2604 23765 2632
rect 23716 2592 23722 2604
rect 23753 2601 23765 2604
rect 23799 2632 23811 2635
rect 25130 2632 25136 2644
rect 23799 2604 24716 2632
rect 25091 2604 25136 2632
rect 23799 2601 23811 2604
rect 23753 2595 23811 2601
rect 20898 2524 20904 2576
rect 20956 2564 20962 2576
rect 24688 2573 24716 2604
rect 25130 2592 25136 2604
rect 25188 2592 25194 2644
rect 21729 2567 21787 2573
rect 21729 2564 21741 2567
rect 20956 2536 21741 2564
rect 20956 2524 20962 2536
rect 21729 2533 21741 2536
rect 21775 2533 21787 2567
rect 21729 2527 21787 2533
rect 24581 2567 24639 2573
rect 24581 2533 24593 2567
rect 24627 2533 24639 2567
rect 24581 2527 24639 2533
rect 24673 2567 24731 2573
rect 24673 2533 24685 2567
rect 24719 2533 24731 2567
rect 24673 2527 24731 2533
rect 19981 2499 20039 2505
rect 19981 2496 19993 2499
rect 19567 2468 19748 2496
rect 19812 2468 19993 2496
rect 19567 2465 19579 2468
rect 19521 2459 19579 2465
rect 15473 2431 15531 2437
rect 15473 2428 15485 2431
rect 14844 2400 15485 2428
rect 14277 2391 14335 2397
rect 15473 2397 15485 2400
rect 15519 2397 15531 2431
rect 18969 2431 19027 2437
rect 18969 2428 18981 2431
rect 15473 2391 15531 2397
rect 17696 2400 18981 2428
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 8260 2264 8585 2292
rect 8260 2252 8266 2264
rect 8573 2261 8585 2264
rect 8619 2292 8631 2295
rect 8938 2292 8944 2304
rect 8619 2264 8944 2292
rect 8619 2261 8631 2264
rect 8573 2255 8631 2261
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 12894 2292 12900 2304
rect 12855 2264 12900 2292
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 13262 2292 13268 2304
rect 13223 2264 13268 2292
rect 13262 2252 13268 2264
rect 13320 2252 13326 2304
rect 13630 2292 13636 2304
rect 13591 2264 13636 2292
rect 13630 2252 13636 2264
rect 13688 2252 13694 2304
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 14734 2292 14740 2304
rect 13955 2264 14740 2292
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17696 2301 17724 2400
rect 18969 2397 18981 2400
rect 19015 2428 19027 2431
rect 19058 2428 19064 2440
rect 19015 2400 19064 2428
rect 19015 2397 19027 2400
rect 18969 2391 19027 2397
rect 19058 2388 19064 2400
rect 19116 2388 19122 2440
rect 19720 2428 19748 2468
rect 19981 2465 19993 2468
rect 20027 2465 20039 2499
rect 21542 2496 21548 2508
rect 19981 2459 20039 2465
rect 20088 2468 21548 2496
rect 20088 2428 20116 2468
rect 21542 2456 21548 2468
rect 21600 2496 21606 2508
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 21600 2468 21833 2496
rect 21600 2456 21606 2468
rect 21821 2465 21833 2468
rect 21867 2465 21879 2499
rect 21821 2459 21879 2465
rect 21910 2456 21916 2508
rect 21968 2496 21974 2508
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 21968 2468 22753 2496
rect 21968 2456 21974 2468
rect 22741 2465 22753 2468
rect 22787 2496 22799 2499
rect 23293 2499 23351 2505
rect 23293 2496 23305 2499
rect 22787 2468 23305 2496
rect 22787 2465 22799 2468
rect 22741 2459 22799 2465
rect 23293 2465 23305 2468
rect 23339 2465 23351 2499
rect 23293 2459 23351 2465
rect 23750 2456 23756 2508
rect 23808 2496 23814 2508
rect 24596 2496 24624 2527
rect 26053 2499 26111 2505
rect 26053 2496 26065 2499
rect 23808 2468 26065 2496
rect 23808 2456 23814 2468
rect 26053 2465 26065 2468
rect 26099 2465 26111 2499
rect 26053 2459 26111 2465
rect 19720 2400 20116 2428
rect 20625 2431 20683 2437
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 21726 2428 21732 2440
rect 20671 2400 21732 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 20070 2320 20076 2372
rect 20128 2360 20134 2372
rect 20640 2360 20668 2391
rect 21726 2388 21732 2400
rect 21784 2388 21790 2440
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23532 2400 24593 2428
rect 23532 2388 23538 2400
rect 24581 2397 24593 2400
rect 24627 2428 24639 2431
rect 25406 2428 25412 2440
rect 24627 2400 25084 2428
rect 25367 2400 25412 2428
rect 24627 2397 24639 2400
rect 24581 2391 24639 2397
rect 20128 2332 20668 2360
rect 21269 2363 21327 2369
rect 20128 2320 20134 2332
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 21358 2360 21364 2372
rect 21315 2332 21364 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 21358 2320 21364 2332
rect 21416 2320 21422 2372
rect 22925 2363 22983 2369
rect 22925 2329 22937 2363
rect 22971 2360 22983 2363
rect 24026 2360 24032 2372
rect 22971 2332 24032 2360
rect 22971 2329 22983 2332
rect 22925 2323 22983 2329
rect 24026 2320 24032 2332
rect 24084 2320 24090 2372
rect 24121 2363 24179 2369
rect 24121 2329 24133 2363
rect 24167 2360 24179 2363
rect 24762 2360 24768 2372
rect 24167 2332 24768 2360
rect 24167 2329 24179 2332
rect 24121 2323 24179 2329
rect 24762 2320 24768 2332
rect 24820 2320 24826 2372
rect 25056 2360 25084 2400
rect 25406 2388 25412 2400
rect 25464 2388 25470 2440
rect 25590 2428 25596 2440
rect 25551 2400 25596 2428
rect 25590 2388 25596 2400
rect 25648 2388 25654 2440
rect 26421 2363 26479 2369
rect 26421 2360 26433 2363
rect 25056 2332 26433 2360
rect 26421 2329 26433 2332
rect 26467 2329 26479 2363
rect 26421 2323 26479 2329
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 18414 2292 18420 2304
rect 18375 2264 18420 2292
rect 17681 2255 17739 2261
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 20162 2292 20168 2304
rect 20123 2264 20168 2292
rect 20162 2252 20168 2264
rect 20220 2252 20226 2304
rect 20898 2292 20904 2304
rect 20859 2264 20904 2292
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 23658 2252 23664 2304
rect 23716 2292 23722 2304
rect 25222 2292 25228 2304
rect 23716 2264 25228 2292
rect 23716 2252 23722 2264
rect 25222 2252 25228 2264
rect 25280 2252 25286 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 14642 2048 14648 2100
rect 14700 2088 14706 2100
rect 15654 2088 15660 2100
rect 14700 2060 15660 2088
rect 14700 2048 14706 2060
rect 15654 2048 15660 2060
rect 15712 2048 15718 2100
rect 24118 2048 24124 2100
rect 24176 2088 24182 2100
rect 25774 2088 25780 2100
rect 24176 2060 25780 2088
rect 24176 2048 24182 2060
rect 25774 2048 25780 2060
rect 25832 2048 25838 2100
rect 11514 1980 11520 2032
rect 11572 2020 11578 2032
rect 18598 2020 18604 2032
rect 11572 1992 18604 2020
rect 11572 1980 11578 1992
rect 18598 1980 18604 1992
rect 18656 1980 18662 2032
<< via1 >>
rect 10784 26800 10836 26852
rect 17592 26800 17644 26852
rect 25228 26732 25280 26784
rect 7564 26664 7616 26716
rect 9588 26664 9640 26716
rect 12440 26596 12492 26648
rect 19432 26596 19484 26648
rect 7564 26528 7616 26580
rect 20812 26528 20864 26580
rect 11704 26460 11756 26512
rect 24768 26460 24820 26512
rect 13176 26392 13228 26444
rect 11520 26324 11572 26376
rect 13360 26324 13412 26376
rect 16028 26324 16080 26376
rect 4344 26256 4396 26308
rect 20444 26256 20496 26308
rect 1308 26188 1360 26240
rect 14464 26188 14516 26240
rect 25504 26188 25556 26240
rect 4712 26120 4764 26172
rect 9864 26120 9916 26172
rect 10048 26120 10100 26172
rect 21548 26120 21600 26172
rect 7748 26052 7800 26104
rect 17040 26052 17092 26104
rect 18880 26052 18932 26104
rect 24308 26052 24360 26104
rect 3056 25984 3108 26036
rect 8760 25984 8812 26036
rect 19800 25984 19852 26036
rect 26056 25984 26108 26036
rect 6920 25916 6972 25968
rect 13912 25916 13964 25968
rect 15660 25916 15712 25968
rect 17868 25916 17920 25968
rect 1952 25848 2004 25900
rect 7288 25848 7340 25900
rect 848 25644 900 25696
rect 14556 25780 14608 25832
rect 14740 25780 14792 25832
rect 23204 25848 23256 25900
rect 23756 25780 23808 25832
rect 18696 25712 18748 25764
rect 18788 25712 18840 25764
rect 27620 25712 27672 25764
rect 9956 25644 10008 25696
rect 11428 25644 11480 25696
rect 22100 25644 22152 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 7748 25440 7800 25492
rect 8760 25483 8812 25492
rect 8760 25449 8769 25483
rect 8769 25449 8803 25483
rect 8803 25449 8812 25483
rect 8760 25440 8812 25449
rect 10048 25483 10100 25492
rect 10048 25449 10057 25483
rect 10057 25449 10091 25483
rect 10091 25449 10100 25483
rect 10048 25440 10100 25449
rect 11060 25440 11112 25492
rect 13084 25440 13136 25492
rect 14096 25440 14148 25492
rect 14740 25440 14792 25492
rect 14924 25483 14976 25492
rect 14924 25449 14933 25483
rect 14933 25449 14967 25483
rect 14967 25449 14976 25483
rect 14924 25440 14976 25449
rect 15568 25440 15620 25492
rect 18788 25440 18840 25492
rect 20904 25440 20956 25492
rect 24768 25440 24820 25492
rect 6276 25372 6328 25424
rect 10784 25372 10836 25424
rect 13268 25372 13320 25424
rect 14832 25372 14884 25424
rect 15844 25415 15896 25424
rect 15844 25381 15853 25415
rect 15853 25381 15887 25415
rect 15887 25381 15896 25415
rect 15844 25372 15896 25381
rect 7748 25304 7800 25356
rect 9036 25304 9088 25356
rect 10968 25304 11020 25356
rect 11336 25347 11388 25356
rect 11336 25313 11345 25347
rect 11345 25313 11379 25347
rect 11379 25313 11388 25347
rect 11336 25304 11388 25313
rect 11796 25304 11848 25356
rect 12532 25304 12584 25356
rect 13360 25304 13412 25356
rect 14188 25304 14240 25356
rect 14372 25304 14424 25356
rect 15476 25304 15528 25356
rect 6460 25236 6512 25288
rect 8208 25168 8260 25220
rect 10048 25236 10100 25288
rect 10784 25236 10836 25288
rect 12808 25236 12860 25288
rect 16672 25236 16724 25288
rect 24860 25372 24912 25424
rect 6644 25143 6696 25152
rect 6644 25109 6653 25143
rect 6653 25109 6687 25143
rect 6687 25109 6696 25143
rect 6644 25100 6696 25109
rect 7840 25100 7892 25152
rect 8024 25143 8076 25152
rect 8024 25109 8033 25143
rect 8033 25109 8067 25143
rect 8067 25109 8076 25143
rect 8024 25100 8076 25109
rect 8392 25143 8444 25152
rect 8392 25109 8401 25143
rect 8401 25109 8435 25143
rect 8435 25109 8444 25143
rect 8392 25100 8444 25109
rect 9680 25100 9732 25152
rect 12532 25100 12584 25152
rect 12716 25143 12768 25152
rect 12716 25109 12725 25143
rect 12725 25109 12759 25143
rect 12759 25109 12768 25143
rect 12716 25100 12768 25109
rect 12992 25168 13044 25220
rect 18512 25304 18564 25356
rect 19524 25347 19576 25356
rect 19524 25313 19533 25347
rect 19533 25313 19567 25347
rect 19567 25313 19576 25347
rect 19524 25304 19576 25313
rect 21272 25304 21324 25356
rect 23020 25304 23072 25356
rect 24124 25304 24176 25356
rect 17500 25168 17552 25220
rect 25320 25236 25372 25288
rect 13820 25100 13872 25152
rect 14004 25143 14056 25152
rect 14004 25109 14013 25143
rect 14013 25109 14047 25143
rect 14047 25109 14056 25143
rect 14004 25100 14056 25109
rect 14372 25100 14424 25152
rect 16028 25100 16080 25152
rect 18236 25100 18288 25152
rect 22376 25168 22428 25220
rect 24676 25168 24728 25220
rect 19432 25100 19484 25152
rect 20076 25143 20128 25152
rect 20076 25109 20085 25143
rect 20085 25109 20119 25143
rect 20119 25109 20128 25143
rect 20076 25100 20128 25109
rect 20628 25100 20680 25152
rect 21640 25100 21692 25152
rect 22284 25143 22336 25152
rect 22284 25109 22293 25143
rect 22293 25109 22327 25143
rect 22327 25109 22336 25143
rect 22284 25100 22336 25109
rect 23664 25143 23716 25152
rect 23664 25109 23673 25143
rect 23673 25109 23707 25143
rect 23707 25109 23716 25143
rect 23664 25100 23716 25109
rect 24768 25143 24820 25152
rect 24768 25109 24777 25143
rect 24777 25109 24811 25143
rect 24811 25109 24820 25143
rect 24768 25100 24820 25109
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 6092 24896 6144 24948
rect 11428 24939 11480 24948
rect 1676 24828 1728 24880
rect 8944 24828 8996 24880
rect 11060 24871 11112 24880
rect 6920 24760 6972 24812
rect 11060 24837 11069 24871
rect 11069 24837 11103 24871
rect 11103 24837 11112 24871
rect 11060 24828 11112 24837
rect 11428 24905 11437 24939
rect 11437 24905 11471 24939
rect 11471 24905 11480 24939
rect 11428 24896 11480 24905
rect 15936 24896 15988 24948
rect 17500 24939 17552 24948
rect 17500 24905 17509 24939
rect 17509 24905 17543 24939
rect 17543 24905 17552 24939
rect 17500 24896 17552 24905
rect 19984 24896 20036 24948
rect 24216 24896 24268 24948
rect 11796 24828 11848 24880
rect 13636 24828 13688 24880
rect 13820 24828 13872 24880
rect 15568 24828 15620 24880
rect 15660 24828 15712 24880
rect 16120 24828 16172 24880
rect 20260 24828 20312 24880
rect 11336 24760 11388 24812
rect 13084 24760 13136 24812
rect 14096 24760 14148 24812
rect 6736 24692 6788 24744
rect 8024 24692 8076 24744
rect 7104 24624 7156 24676
rect 8484 24667 8536 24676
rect 8484 24633 8493 24667
rect 8493 24633 8527 24667
rect 8527 24633 8536 24667
rect 8484 24624 8536 24633
rect 14004 24735 14056 24744
rect 8760 24624 8812 24676
rect 9864 24667 9916 24676
rect 9864 24633 9873 24667
rect 9873 24633 9907 24667
rect 9907 24633 9916 24667
rect 9864 24624 9916 24633
rect 10140 24667 10192 24676
rect 10140 24633 10149 24667
rect 10149 24633 10183 24667
rect 10183 24633 10192 24667
rect 10140 24624 10192 24633
rect 14004 24701 14013 24735
rect 14013 24701 14047 24735
rect 14047 24701 14056 24735
rect 14004 24692 14056 24701
rect 15292 24760 15344 24812
rect 23020 24828 23072 24880
rect 25136 24828 25188 24880
rect 22192 24803 22244 24812
rect 22192 24769 22201 24803
rect 22201 24769 22235 24803
rect 22235 24769 22244 24803
rect 22192 24760 22244 24769
rect 15384 24692 15436 24744
rect 16396 24735 16448 24744
rect 16396 24701 16405 24735
rect 16405 24701 16439 24735
rect 16439 24701 16448 24735
rect 16396 24692 16448 24701
rect 18052 24692 18104 24744
rect 20076 24692 20128 24744
rect 23480 24692 23532 24744
rect 24124 24692 24176 24744
rect 25044 24692 25096 24744
rect 12992 24667 13044 24676
rect 12992 24633 13001 24667
rect 13001 24633 13035 24667
rect 13035 24633 13044 24667
rect 12992 24624 13044 24633
rect 13084 24667 13136 24676
rect 13084 24633 13093 24667
rect 13093 24633 13127 24667
rect 13127 24633 13136 24667
rect 13084 24624 13136 24633
rect 14280 24667 14332 24676
rect 14280 24633 14289 24667
rect 14289 24633 14323 24667
rect 14323 24633 14332 24667
rect 14280 24624 14332 24633
rect 15200 24624 15252 24676
rect 16856 24624 16908 24676
rect 17868 24624 17920 24676
rect 20628 24667 20680 24676
rect 4712 24556 4764 24608
rect 5264 24599 5316 24608
rect 5264 24565 5273 24599
rect 5273 24565 5307 24599
rect 5307 24565 5316 24599
rect 5264 24556 5316 24565
rect 5540 24599 5592 24608
rect 5540 24565 5549 24599
rect 5549 24565 5583 24599
rect 5583 24565 5592 24599
rect 5540 24556 5592 24565
rect 7012 24599 7064 24608
rect 7012 24565 7021 24599
rect 7021 24565 7055 24599
rect 7055 24565 7064 24599
rect 7012 24556 7064 24565
rect 7472 24556 7524 24608
rect 9036 24599 9088 24608
rect 9036 24565 9045 24599
rect 9045 24565 9079 24599
rect 9079 24565 9088 24599
rect 9036 24556 9088 24565
rect 9588 24599 9640 24608
rect 9588 24565 9621 24599
rect 9621 24565 9640 24599
rect 10048 24599 10100 24608
rect 9588 24556 9640 24565
rect 10048 24565 10057 24599
rect 10057 24565 10091 24599
rect 10091 24565 10100 24599
rect 10048 24556 10100 24565
rect 10968 24556 11020 24608
rect 11612 24556 11664 24608
rect 12532 24599 12584 24608
rect 12532 24565 12565 24599
rect 12565 24565 12584 24599
rect 12532 24556 12584 24565
rect 13360 24556 13412 24608
rect 14188 24556 14240 24608
rect 15660 24556 15712 24608
rect 18328 24556 18380 24608
rect 18512 24599 18564 24608
rect 18512 24565 18521 24599
rect 18521 24565 18555 24599
rect 18555 24565 18564 24599
rect 18512 24556 18564 24565
rect 19064 24599 19116 24608
rect 19064 24565 19073 24599
rect 19073 24565 19107 24599
rect 19107 24565 19116 24599
rect 19064 24556 19116 24565
rect 19432 24556 19484 24608
rect 20076 24599 20128 24608
rect 20076 24565 20109 24599
rect 20109 24565 20128 24599
rect 20628 24633 20637 24667
rect 20637 24633 20671 24667
rect 20671 24633 20680 24667
rect 20628 24624 20680 24633
rect 20076 24556 20128 24565
rect 21272 24556 21324 24608
rect 22008 24624 22060 24676
rect 22284 24667 22336 24676
rect 22284 24633 22293 24667
rect 22293 24633 22327 24667
rect 22327 24633 22336 24667
rect 22284 24624 22336 24633
rect 22928 24624 22980 24676
rect 23664 24624 23716 24676
rect 21824 24556 21876 24608
rect 23296 24556 23348 24608
rect 23480 24599 23532 24608
rect 23480 24565 23489 24599
rect 23489 24565 23523 24599
rect 23523 24565 23532 24599
rect 23480 24556 23532 24565
rect 23756 24599 23808 24608
rect 23756 24565 23789 24599
rect 23789 24565 23808 24599
rect 24308 24667 24360 24676
rect 24308 24633 24317 24667
rect 24317 24633 24351 24667
rect 24351 24633 24360 24667
rect 24308 24624 24360 24633
rect 23756 24556 23808 24565
rect 25412 24599 25464 24608
rect 25412 24565 25421 24599
rect 25421 24565 25455 24599
rect 25455 24565 25464 24599
rect 25412 24556 25464 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 6092 24352 6144 24404
rect 6460 24395 6512 24404
rect 6460 24361 6469 24395
rect 6469 24361 6503 24395
rect 6503 24361 6512 24395
rect 6460 24352 6512 24361
rect 7288 24352 7340 24404
rect 11244 24352 11296 24404
rect 12532 24352 12584 24404
rect 12716 24352 12768 24404
rect 15476 24395 15528 24404
rect 15476 24361 15485 24395
rect 15485 24361 15519 24395
rect 15519 24361 15528 24395
rect 15476 24352 15528 24361
rect 15844 24395 15896 24404
rect 15844 24361 15853 24395
rect 15853 24361 15887 24395
rect 15887 24361 15896 24395
rect 15844 24352 15896 24361
rect 16120 24352 16172 24404
rect 16856 24352 16908 24404
rect 18788 24395 18840 24404
rect 18788 24361 18797 24395
rect 18797 24361 18831 24395
rect 18831 24361 18840 24395
rect 18788 24352 18840 24361
rect 19984 24352 20036 24404
rect 20260 24395 20312 24404
rect 20260 24361 20269 24395
rect 20269 24361 20303 24395
rect 20303 24361 20312 24395
rect 20260 24352 20312 24361
rect 23020 24352 23072 24404
rect 2228 24216 2280 24268
rect 8852 24284 8904 24336
rect 13452 24284 13504 24336
rect 16948 24284 17000 24336
rect 18328 24327 18380 24336
rect 18328 24293 18337 24327
rect 18337 24293 18371 24327
rect 18371 24293 18380 24327
rect 18328 24284 18380 24293
rect 21088 24284 21140 24336
rect 22836 24284 22888 24336
rect 6920 24259 6972 24268
rect 6920 24225 6929 24259
rect 6929 24225 6963 24259
rect 6963 24225 6972 24259
rect 6920 24216 6972 24225
rect 7748 24216 7800 24268
rect 8024 24216 8076 24268
rect 8300 24216 8352 24268
rect 5172 24148 5224 24200
rect 6184 24148 6236 24200
rect 5356 24080 5408 24132
rect 11428 24216 11480 24268
rect 11980 24216 12032 24268
rect 10600 24191 10652 24200
rect 10600 24157 10609 24191
rect 10609 24157 10643 24191
rect 10643 24157 10652 24191
rect 10600 24148 10652 24157
rect 12440 24148 12492 24200
rect 12900 24148 12952 24200
rect 8208 24080 8260 24132
rect 12808 24080 12860 24132
rect 13268 24123 13320 24132
rect 13268 24089 13277 24123
rect 13277 24089 13311 24123
rect 13311 24089 13320 24123
rect 13268 24080 13320 24089
rect 14556 24259 14608 24268
rect 14556 24225 14565 24259
rect 14565 24225 14599 24259
rect 14599 24225 14608 24259
rect 14556 24216 14608 24225
rect 16580 24216 16632 24268
rect 19708 24259 19760 24268
rect 19708 24225 19717 24259
rect 19717 24225 19751 24259
rect 19751 24225 19760 24259
rect 19708 24216 19760 24225
rect 23296 24216 23348 24268
rect 24308 24216 24360 24268
rect 24952 24216 25004 24268
rect 13544 24080 13596 24132
rect 16212 24148 16264 24200
rect 18052 24148 18104 24200
rect 18236 24191 18288 24200
rect 18236 24157 18245 24191
rect 18245 24157 18279 24191
rect 18279 24157 18288 24191
rect 18236 24148 18288 24157
rect 18420 24191 18472 24200
rect 18420 24157 18429 24191
rect 18429 24157 18463 24191
rect 18463 24157 18472 24191
rect 18420 24148 18472 24157
rect 21916 24191 21968 24200
rect 21916 24157 21925 24191
rect 21925 24157 21959 24191
rect 21959 24157 21968 24191
rect 21916 24148 21968 24157
rect 22100 24191 22152 24200
rect 22100 24157 22109 24191
rect 22109 24157 22143 24191
rect 22143 24157 22152 24191
rect 22100 24148 22152 24157
rect 23388 24148 23440 24200
rect 6552 24012 6604 24064
rect 6828 24055 6880 24064
rect 6828 24021 6837 24055
rect 6837 24021 6871 24055
rect 6871 24021 6880 24055
rect 6828 24012 6880 24021
rect 7748 24012 7800 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 9496 24055 9548 24064
rect 9496 24021 9505 24055
rect 9505 24021 9539 24055
rect 9539 24021 9548 24055
rect 9496 24012 9548 24021
rect 9864 24055 9916 24064
rect 9864 24021 9873 24055
rect 9873 24021 9907 24055
rect 9907 24021 9916 24055
rect 9864 24012 9916 24021
rect 11980 24055 12032 24064
rect 11980 24021 11989 24055
rect 11989 24021 12023 24055
rect 12023 24021 12032 24055
rect 11980 24012 12032 24021
rect 14740 24080 14792 24132
rect 18696 24080 18748 24132
rect 21824 24080 21876 24132
rect 16304 24055 16356 24064
rect 16304 24021 16313 24055
rect 16313 24021 16347 24055
rect 16347 24021 16356 24055
rect 16304 24012 16356 24021
rect 17592 24055 17644 24064
rect 17592 24021 17601 24055
rect 17601 24021 17635 24055
rect 17635 24021 17644 24055
rect 17592 24012 17644 24021
rect 18236 24012 18288 24064
rect 19156 24055 19208 24064
rect 19156 24021 19165 24055
rect 19165 24021 19199 24055
rect 19199 24021 19208 24055
rect 19156 24012 19208 24021
rect 19524 24055 19576 24064
rect 19524 24021 19533 24055
rect 19533 24021 19567 24055
rect 19567 24021 19576 24055
rect 19524 24012 19576 24021
rect 20720 24055 20772 24064
rect 20720 24021 20729 24055
rect 20729 24021 20763 24055
rect 20763 24021 20772 24055
rect 20720 24012 20772 24021
rect 21548 24055 21600 24064
rect 21548 24021 21557 24055
rect 21557 24021 21591 24055
rect 21591 24021 21600 24055
rect 21548 24012 21600 24021
rect 22560 24055 22612 24064
rect 22560 24021 22569 24055
rect 22569 24021 22603 24055
rect 22603 24021 22612 24055
rect 22560 24012 22612 24021
rect 23204 24055 23256 24064
rect 23204 24021 23213 24055
rect 23213 24021 23247 24055
rect 23247 24021 23256 24055
rect 23204 24012 23256 24021
rect 24124 24055 24176 24064
rect 24124 24021 24133 24055
rect 24133 24021 24167 24055
rect 24167 24021 24176 24055
rect 24124 24012 24176 24021
rect 24768 24012 24820 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1400 23808 1452 23860
rect 6276 23808 6328 23860
rect 7564 23851 7616 23860
rect 7564 23817 7573 23851
rect 7573 23817 7607 23851
rect 7607 23817 7616 23851
rect 7564 23808 7616 23817
rect 8208 23808 8260 23860
rect 9036 23808 9088 23860
rect 12348 23808 12400 23860
rect 12532 23851 12584 23860
rect 12532 23817 12541 23851
rect 12541 23817 12575 23851
rect 12575 23817 12584 23851
rect 12532 23808 12584 23817
rect 14556 23808 14608 23860
rect 11428 23783 11480 23792
rect 11428 23749 11437 23783
rect 11437 23749 11471 23783
rect 11471 23749 11480 23783
rect 11428 23740 11480 23749
rect 12808 23740 12860 23792
rect 15752 23808 15804 23860
rect 18144 23851 18196 23860
rect 18144 23817 18153 23851
rect 18153 23817 18187 23851
rect 18187 23817 18196 23851
rect 18144 23808 18196 23817
rect 18972 23808 19024 23860
rect 8024 23715 8076 23724
rect 8024 23681 8033 23715
rect 8033 23681 8067 23715
rect 8067 23681 8076 23715
rect 8024 23672 8076 23681
rect 11980 23672 12032 23724
rect 13084 23715 13136 23724
rect 13084 23681 13093 23715
rect 13093 23681 13127 23715
rect 13127 23681 13136 23715
rect 13084 23672 13136 23681
rect 18420 23672 18472 23724
rect 4620 23604 4672 23656
rect 9036 23647 9088 23656
rect 3976 23536 4028 23588
rect 4804 23536 4856 23588
rect 6276 23536 6328 23588
rect 2228 23468 2280 23520
rect 2412 23511 2464 23520
rect 2412 23477 2421 23511
rect 2421 23477 2455 23511
rect 2455 23477 2464 23511
rect 2412 23468 2464 23477
rect 3240 23511 3292 23520
rect 3240 23477 3249 23511
rect 3249 23477 3283 23511
rect 3283 23477 3292 23511
rect 3240 23468 3292 23477
rect 3792 23468 3844 23520
rect 4896 23468 4948 23520
rect 9036 23613 9045 23647
rect 9045 23613 9079 23647
rect 9079 23613 9088 23647
rect 9036 23604 9088 23613
rect 9128 23604 9180 23656
rect 10140 23604 10192 23656
rect 10600 23604 10652 23656
rect 6920 23536 6972 23588
rect 7380 23536 7432 23588
rect 7748 23536 7800 23588
rect 6736 23468 6788 23520
rect 7564 23468 7616 23520
rect 8300 23468 8352 23520
rect 8852 23511 8904 23520
rect 8852 23477 8861 23511
rect 8861 23477 8895 23511
rect 8895 23477 8904 23511
rect 8852 23468 8904 23477
rect 9680 23468 9732 23520
rect 12348 23536 12400 23588
rect 11152 23468 11204 23520
rect 12624 23604 12676 23656
rect 13452 23647 13504 23656
rect 13452 23613 13461 23647
rect 13461 23613 13495 23647
rect 13495 23613 13504 23647
rect 13452 23604 13504 23613
rect 12716 23536 12768 23588
rect 13268 23536 13320 23588
rect 13544 23536 13596 23588
rect 13452 23468 13504 23520
rect 16488 23604 16540 23656
rect 17592 23604 17644 23656
rect 18328 23604 18380 23656
rect 18788 23672 18840 23724
rect 19064 23740 19116 23792
rect 19708 23808 19760 23860
rect 22100 23808 22152 23860
rect 22836 23851 22888 23860
rect 22836 23817 22845 23851
rect 22845 23817 22879 23851
rect 22879 23817 22888 23851
rect 22836 23808 22888 23817
rect 25688 23851 25740 23860
rect 25688 23817 25697 23851
rect 25697 23817 25731 23851
rect 25731 23817 25740 23851
rect 25688 23808 25740 23817
rect 20812 23740 20864 23792
rect 21364 23783 21416 23792
rect 21364 23749 21373 23783
rect 21373 23749 21407 23783
rect 21407 23749 21416 23783
rect 21364 23740 21416 23749
rect 23480 23740 23532 23792
rect 24032 23783 24084 23792
rect 24032 23749 24041 23783
rect 24041 23749 24075 23783
rect 24075 23749 24084 23783
rect 24032 23740 24084 23749
rect 18972 23604 19024 23656
rect 21640 23647 21692 23656
rect 21640 23613 21649 23647
rect 21649 23613 21683 23647
rect 21683 23613 21692 23647
rect 21640 23604 21692 23613
rect 14740 23536 14792 23588
rect 15292 23536 15344 23588
rect 15752 23536 15804 23588
rect 18144 23536 18196 23588
rect 18604 23579 18656 23588
rect 18604 23545 18613 23579
rect 18613 23545 18647 23579
rect 18647 23545 18656 23579
rect 18604 23536 18656 23545
rect 20352 23579 20404 23588
rect 20352 23545 20361 23579
rect 20361 23545 20395 23579
rect 20395 23545 20404 23579
rect 20352 23536 20404 23545
rect 16212 23511 16264 23520
rect 16212 23477 16221 23511
rect 16221 23477 16255 23511
rect 16255 23477 16264 23511
rect 16212 23468 16264 23477
rect 16672 23468 16724 23520
rect 19984 23468 20036 23520
rect 21088 23468 21140 23520
rect 21824 23672 21876 23724
rect 24216 23672 24268 23724
rect 22560 23604 22612 23656
rect 25504 23647 25556 23656
rect 25504 23613 25513 23647
rect 25513 23613 25547 23647
rect 25547 23613 25556 23647
rect 25504 23604 25556 23613
rect 22100 23536 22152 23588
rect 22836 23536 22888 23588
rect 23388 23536 23440 23588
rect 23480 23536 23532 23588
rect 24124 23536 24176 23588
rect 22192 23468 22244 23520
rect 23020 23468 23072 23520
rect 23940 23468 23992 23520
rect 24952 23511 25004 23520
rect 24952 23477 24961 23511
rect 24961 23477 24995 23511
rect 24995 23477 25004 23511
rect 24952 23468 25004 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1492 23264 1544 23316
rect 5632 23264 5684 23316
rect 6552 23196 6604 23248
rect 8392 23239 8444 23248
rect 8392 23205 8401 23239
rect 8401 23205 8435 23239
rect 8435 23205 8444 23239
rect 8392 23196 8444 23205
rect 8576 23239 8628 23248
rect 8576 23205 8585 23239
rect 8585 23205 8619 23239
rect 8619 23205 8628 23239
rect 8576 23196 8628 23205
rect 8760 23196 8812 23248
rect 9128 23196 9180 23248
rect 12440 23264 12492 23316
rect 13268 23307 13320 23316
rect 13268 23273 13277 23307
rect 13277 23273 13311 23307
rect 13311 23273 13320 23307
rect 13268 23264 13320 23273
rect 15936 23264 15988 23316
rect 16212 23264 16264 23316
rect 16580 23264 16632 23316
rect 18144 23307 18196 23316
rect 18144 23273 18153 23307
rect 18153 23273 18187 23307
rect 18187 23273 18196 23307
rect 18144 23264 18196 23273
rect 19340 23264 19392 23316
rect 20076 23264 20128 23316
rect 20352 23264 20404 23316
rect 20720 23264 20772 23316
rect 21456 23307 21508 23316
rect 21456 23273 21465 23307
rect 21465 23273 21499 23307
rect 21499 23273 21508 23307
rect 21456 23264 21508 23273
rect 21916 23307 21968 23316
rect 21916 23273 21925 23307
rect 21925 23273 21959 23307
rect 21959 23273 21968 23307
rect 21916 23264 21968 23273
rect 24860 23307 24912 23316
rect 11428 23196 11480 23248
rect 15476 23196 15528 23248
rect 15844 23239 15896 23248
rect 15844 23205 15853 23239
rect 15853 23205 15887 23239
rect 15887 23205 15896 23239
rect 15844 23196 15896 23205
rect 17408 23239 17460 23248
rect 17408 23205 17417 23239
rect 17417 23205 17451 23239
rect 17451 23205 17460 23239
rect 17408 23196 17460 23205
rect 17960 23196 18012 23248
rect 18880 23196 18932 23248
rect 18972 23239 19024 23248
rect 18972 23205 18981 23239
rect 18981 23205 19015 23239
rect 19015 23205 19024 23239
rect 18972 23196 19024 23205
rect 23572 23196 23624 23248
rect 24860 23273 24869 23307
rect 24869 23273 24903 23307
rect 24903 23273 24912 23307
rect 24860 23264 24912 23273
rect 2780 23128 2832 23180
rect 4988 23128 5040 23180
rect 6920 23128 6972 23180
rect 10232 23128 10284 23180
rect 11152 23128 11204 23180
rect 12164 23128 12216 23180
rect 13912 23171 13964 23180
rect 13912 23137 13921 23171
rect 13921 23137 13955 23171
rect 13955 23137 13964 23171
rect 13912 23128 13964 23137
rect 1768 23060 1820 23112
rect 5080 23060 5132 23112
rect 7012 23103 7064 23112
rect 7012 23069 7021 23103
rect 7021 23069 7055 23103
rect 7055 23069 7064 23103
rect 7012 23060 7064 23069
rect 9036 23060 9088 23112
rect 2964 22992 3016 23044
rect 6828 22992 6880 23044
rect 7288 22992 7340 23044
rect 7748 22992 7800 23044
rect 8116 23035 8168 23044
rect 1952 22967 2004 22976
rect 1952 22933 1961 22967
rect 1961 22933 1995 22967
rect 1995 22933 2004 22967
rect 1952 22924 2004 22933
rect 2320 22967 2372 22976
rect 2320 22933 2329 22967
rect 2329 22933 2363 22967
rect 2363 22933 2372 22967
rect 2320 22924 2372 22933
rect 2412 22924 2464 22976
rect 3056 22967 3108 22976
rect 3056 22933 3065 22967
rect 3065 22933 3099 22967
rect 3099 22933 3108 22967
rect 3056 22924 3108 22933
rect 3148 22924 3200 22976
rect 4528 22924 4580 22976
rect 5448 22924 5500 22976
rect 6092 22924 6144 22976
rect 6460 22924 6512 22976
rect 7564 22967 7616 22976
rect 7564 22933 7573 22967
rect 7573 22933 7607 22967
rect 7607 22933 7616 22967
rect 7564 22924 7616 22933
rect 8116 23001 8125 23035
rect 8125 23001 8159 23035
rect 8159 23001 8168 23035
rect 8116 22992 8168 23001
rect 9036 22924 9088 22976
rect 9128 22924 9180 22976
rect 9312 22924 9364 22976
rect 9588 22924 9640 22976
rect 12256 22992 12308 23044
rect 13820 23060 13872 23112
rect 15108 23035 15160 23044
rect 15108 23001 15117 23035
rect 15117 23001 15151 23035
rect 15151 23001 15160 23035
rect 15108 22992 15160 23001
rect 15384 23035 15436 23044
rect 15384 23001 15393 23035
rect 15393 23001 15427 23035
rect 15427 23001 15436 23035
rect 15384 22992 15436 23001
rect 10324 22924 10376 22976
rect 11336 22924 11388 22976
rect 11980 22967 12032 22976
rect 11980 22933 11989 22967
rect 11989 22933 12023 22967
rect 12023 22933 12032 22967
rect 11980 22924 12032 22933
rect 13728 22967 13780 22976
rect 13728 22933 13737 22967
rect 13737 22933 13771 22967
rect 13771 22933 13780 22967
rect 13728 22924 13780 22933
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 15936 22924 15988 22976
rect 18512 23128 18564 23180
rect 21824 23128 21876 23180
rect 22100 23128 22152 23180
rect 24860 23128 24912 23180
rect 17684 23060 17736 23112
rect 16948 23035 17000 23044
rect 16948 23001 16957 23035
rect 16957 23001 16991 23035
rect 16991 23001 17000 23035
rect 16948 22992 17000 23001
rect 21364 23103 21416 23112
rect 21364 23069 21373 23103
rect 21373 23069 21407 23103
rect 21407 23069 21416 23103
rect 21364 23060 21416 23069
rect 21548 23103 21600 23112
rect 21548 23069 21557 23103
rect 21557 23069 21591 23103
rect 21591 23069 21600 23103
rect 21548 23060 21600 23069
rect 22652 23060 22704 23112
rect 24952 23103 25004 23112
rect 19800 22992 19852 23044
rect 20352 22992 20404 23044
rect 18052 22924 18104 22976
rect 18144 22924 18196 22976
rect 19340 22924 19392 22976
rect 19432 22924 19484 22976
rect 19984 22924 20036 22976
rect 20536 22967 20588 22976
rect 20536 22933 20545 22967
rect 20545 22933 20579 22967
rect 20579 22933 20588 22967
rect 20536 22924 20588 22933
rect 21640 22992 21692 23044
rect 24952 23069 24961 23103
rect 24961 23069 24995 23103
rect 24995 23069 25004 23103
rect 24952 23060 25004 23069
rect 23756 22992 23808 23044
rect 24124 22992 24176 23044
rect 21180 22924 21232 22976
rect 22192 22924 22244 22976
rect 22744 22924 22796 22976
rect 23940 22967 23992 22976
rect 23940 22933 23949 22967
rect 23949 22933 23983 22967
rect 23983 22933 23992 22967
rect 23940 22924 23992 22933
rect 24676 22924 24728 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2688 22763 2740 22772
rect 2688 22729 2697 22763
rect 2697 22729 2731 22763
rect 2731 22729 2740 22763
rect 2688 22720 2740 22729
rect 6920 22720 6972 22772
rect 8392 22720 8444 22772
rect 8576 22720 8628 22772
rect 10048 22720 10100 22772
rect 11796 22720 11848 22772
rect 14740 22763 14792 22772
rect 14740 22729 14749 22763
rect 14749 22729 14783 22763
rect 14783 22729 14792 22763
rect 14740 22720 14792 22729
rect 15476 22720 15528 22772
rect 16488 22763 16540 22772
rect 16488 22729 16497 22763
rect 16497 22729 16531 22763
rect 16531 22729 16540 22763
rect 16488 22720 16540 22729
rect 17408 22763 17460 22772
rect 17408 22729 17417 22763
rect 17417 22729 17451 22763
rect 17451 22729 17460 22763
rect 17408 22720 17460 22729
rect 21548 22720 21600 22772
rect 23388 22763 23440 22772
rect 23388 22729 23397 22763
rect 23397 22729 23431 22763
rect 23431 22729 23440 22763
rect 23388 22720 23440 22729
rect 25136 22720 25188 22772
rect 1584 22695 1636 22704
rect 1584 22661 1593 22695
rect 1593 22661 1627 22695
rect 1627 22661 1636 22695
rect 1584 22652 1636 22661
rect 4068 22652 4120 22704
rect 8760 22695 8812 22704
rect 1400 22559 1452 22568
rect 1400 22525 1409 22559
rect 1409 22525 1443 22559
rect 1443 22525 1452 22559
rect 1400 22516 1452 22525
rect 2872 22448 2924 22500
rect 4988 22584 5040 22636
rect 5448 22584 5500 22636
rect 6460 22584 6512 22636
rect 5632 22516 5684 22568
rect 4160 22448 4212 22500
rect 6920 22516 6972 22568
rect 8760 22661 8769 22695
rect 8769 22661 8803 22695
rect 8803 22661 8812 22695
rect 8760 22652 8812 22661
rect 16764 22652 16816 22704
rect 17684 22652 17736 22704
rect 19340 22652 19392 22704
rect 19708 22652 19760 22704
rect 19800 22652 19852 22704
rect 23756 22695 23808 22704
rect 23756 22661 23765 22695
rect 23765 22661 23799 22695
rect 23799 22661 23808 22695
rect 23756 22652 23808 22661
rect 24768 22652 24820 22704
rect 7104 22584 7156 22636
rect 8024 22584 8076 22636
rect 10784 22584 10836 22636
rect 11244 22627 11296 22636
rect 11244 22593 11253 22627
rect 11253 22593 11287 22627
rect 11287 22593 11296 22627
rect 11244 22584 11296 22593
rect 11428 22627 11480 22636
rect 11428 22593 11437 22627
rect 11437 22593 11471 22627
rect 11471 22593 11480 22627
rect 11428 22584 11480 22593
rect 21272 22584 21324 22636
rect 22376 22627 22428 22636
rect 22376 22593 22385 22627
rect 22385 22593 22419 22627
rect 22419 22593 22428 22627
rect 22376 22584 22428 22593
rect 7748 22516 7800 22568
rect 8208 22516 8260 22568
rect 10232 22516 10284 22568
rect 12164 22559 12216 22568
rect 12164 22525 12173 22559
rect 12173 22525 12207 22559
rect 12207 22525 12216 22559
rect 12164 22516 12216 22525
rect 9772 22491 9824 22500
rect 9772 22457 9781 22491
rect 9781 22457 9815 22491
rect 9815 22457 9824 22491
rect 9772 22448 9824 22457
rect 10324 22491 10376 22500
rect 10324 22457 10333 22491
rect 10333 22457 10367 22491
rect 10367 22457 10376 22491
rect 13452 22516 13504 22568
rect 14832 22516 14884 22568
rect 10324 22448 10376 22457
rect 1768 22380 1820 22432
rect 2780 22380 2832 22432
rect 3516 22380 3568 22432
rect 5724 22423 5776 22432
rect 5724 22389 5733 22423
rect 5733 22389 5767 22423
rect 5767 22389 5776 22423
rect 5724 22380 5776 22389
rect 6552 22423 6604 22432
rect 6552 22389 6561 22423
rect 6561 22389 6595 22423
rect 6595 22389 6604 22423
rect 6552 22380 6604 22389
rect 7104 22423 7156 22432
rect 7104 22389 7113 22423
rect 7113 22389 7147 22423
rect 7147 22389 7156 22423
rect 7104 22380 7156 22389
rect 7840 22380 7892 22432
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 12440 22380 12492 22432
rect 13728 22448 13780 22500
rect 16488 22448 16540 22500
rect 16856 22448 16908 22500
rect 17500 22516 17552 22568
rect 19340 22516 19392 22568
rect 20536 22516 20588 22568
rect 22100 22559 22152 22568
rect 22100 22525 22109 22559
rect 22109 22525 22143 22559
rect 22143 22525 22152 22559
rect 24124 22584 24176 22636
rect 24952 22584 25004 22636
rect 22100 22516 22152 22525
rect 23848 22516 23900 22568
rect 25228 22559 25280 22568
rect 25228 22525 25237 22559
rect 25237 22525 25271 22559
rect 25271 22525 25280 22559
rect 25228 22516 25280 22525
rect 13268 22380 13320 22432
rect 15844 22380 15896 22432
rect 17224 22423 17276 22432
rect 17224 22389 17233 22423
rect 17233 22389 17267 22423
rect 17267 22389 17276 22423
rect 17224 22380 17276 22389
rect 17868 22380 17920 22432
rect 18236 22448 18288 22500
rect 20444 22448 20496 22500
rect 19340 22380 19392 22432
rect 21364 22448 21416 22500
rect 23664 22448 23716 22500
rect 25320 22448 25372 22500
rect 20720 22380 20772 22432
rect 22192 22380 22244 22432
rect 23388 22380 23440 22432
rect 23480 22380 23532 22432
rect 24860 22380 24912 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1400 22176 1452 22228
rect 2044 22176 2096 22228
rect 5448 22219 5500 22228
rect 5448 22185 5457 22219
rect 5457 22185 5491 22219
rect 5491 22185 5500 22219
rect 5448 22176 5500 22185
rect 7840 22176 7892 22228
rect 11060 22176 11112 22228
rect 12992 22176 13044 22228
rect 17224 22176 17276 22228
rect 18236 22176 18288 22228
rect 4160 22108 4212 22160
rect 7196 22108 7248 22160
rect 2504 22083 2556 22092
rect 2504 22049 2513 22083
rect 2513 22049 2547 22083
rect 2547 22049 2556 22083
rect 2504 22040 2556 22049
rect 3332 22040 3384 22092
rect 7288 22040 7340 22092
rect 8208 22040 8260 22092
rect 1860 21972 1912 22024
rect 3884 21972 3936 22024
rect 4712 21972 4764 22024
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 5540 21972 5592 21981
rect 7012 22015 7064 22024
rect 7012 21981 7021 22015
rect 7021 21981 7055 22015
rect 7055 21981 7064 22015
rect 7012 21972 7064 21981
rect 7840 21972 7892 22024
rect 9128 22108 9180 22160
rect 9404 22108 9456 22160
rect 10232 22151 10284 22160
rect 10232 22117 10241 22151
rect 10241 22117 10275 22151
rect 10275 22117 10284 22151
rect 10232 22108 10284 22117
rect 11428 22108 11480 22160
rect 12072 22108 12124 22160
rect 13912 22108 13964 22160
rect 8852 22040 8904 22092
rect 8944 22040 8996 22092
rect 9772 22040 9824 22092
rect 10876 22040 10928 22092
rect 11704 22040 11756 22092
rect 13544 22040 13596 22092
rect 17776 22108 17828 22160
rect 18880 22151 18932 22160
rect 18880 22117 18889 22151
rect 18889 22117 18923 22151
rect 18923 22117 18932 22151
rect 18880 22108 18932 22117
rect 15384 22040 15436 22092
rect 15568 22083 15620 22092
rect 15568 22049 15577 22083
rect 15577 22049 15611 22083
rect 15611 22049 15620 22083
rect 15568 22040 15620 22049
rect 17132 22040 17184 22092
rect 18052 22040 18104 22092
rect 18972 22040 19024 22092
rect 19156 22040 19208 22092
rect 20812 22176 20864 22228
rect 21456 22219 21508 22228
rect 21456 22185 21465 22219
rect 21465 22185 21499 22219
rect 21499 22185 21508 22219
rect 21456 22176 21508 22185
rect 19616 22151 19668 22160
rect 19616 22117 19625 22151
rect 19625 22117 19659 22151
rect 19659 22117 19668 22151
rect 19616 22108 19668 22117
rect 20996 22151 21048 22160
rect 20996 22117 21021 22151
rect 21021 22117 21048 22151
rect 20996 22108 21048 22117
rect 23388 22108 23440 22160
rect 23756 22176 23808 22228
rect 24216 22108 24268 22160
rect 25780 22176 25832 22228
rect 24768 22108 24820 22160
rect 8576 21972 8628 22024
rect 2596 21904 2648 21956
rect 3516 21904 3568 21956
rect 3700 21904 3752 21956
rect 1584 21879 1636 21888
rect 1584 21845 1593 21879
rect 1593 21845 1627 21879
rect 1627 21845 1636 21879
rect 1584 21836 1636 21845
rect 2412 21879 2464 21888
rect 2412 21845 2421 21879
rect 2421 21845 2455 21879
rect 2455 21845 2464 21879
rect 2412 21836 2464 21845
rect 3056 21879 3108 21888
rect 3056 21845 3065 21879
rect 3065 21845 3099 21879
rect 3099 21845 3108 21879
rect 3056 21836 3108 21845
rect 4160 21904 4212 21956
rect 4988 21947 5040 21956
rect 4988 21913 4997 21947
rect 4997 21913 5031 21947
rect 5031 21913 5040 21947
rect 4988 21904 5040 21913
rect 5632 21904 5684 21956
rect 6368 21904 6420 21956
rect 4252 21879 4304 21888
rect 4252 21845 4261 21879
rect 4261 21845 4295 21879
rect 4295 21845 4304 21879
rect 4252 21836 4304 21845
rect 4436 21836 4488 21888
rect 6000 21879 6052 21888
rect 6000 21845 6009 21879
rect 6009 21845 6043 21879
rect 6043 21845 6052 21879
rect 6000 21836 6052 21845
rect 6184 21836 6236 21888
rect 8392 21836 8444 21888
rect 9404 21972 9456 22024
rect 10508 21972 10560 22024
rect 11796 21972 11848 22024
rect 12256 22015 12308 22024
rect 12256 21981 12265 22015
rect 12265 21981 12299 22015
rect 12299 21981 12308 22015
rect 12256 21972 12308 21981
rect 13728 22015 13780 22024
rect 13728 21981 13737 22015
rect 13737 21981 13771 22015
rect 13771 21981 13780 22015
rect 13728 21972 13780 21981
rect 14004 21972 14056 22024
rect 15108 22015 15160 22024
rect 15108 21981 15117 22015
rect 15117 21981 15151 22015
rect 15151 21981 15160 22015
rect 15108 21972 15160 21981
rect 9864 21904 9916 21956
rect 11336 21904 11388 21956
rect 16488 21904 16540 21956
rect 9220 21836 9272 21888
rect 10784 21879 10836 21888
rect 10784 21845 10793 21879
rect 10793 21845 10827 21879
rect 10827 21845 10836 21879
rect 10784 21836 10836 21845
rect 11060 21836 11112 21888
rect 12716 21879 12768 21888
rect 12716 21845 12725 21879
rect 12725 21845 12759 21879
rect 12759 21845 12768 21879
rect 12716 21836 12768 21845
rect 14280 21879 14332 21888
rect 14280 21845 14289 21879
rect 14289 21845 14323 21879
rect 14323 21845 14332 21879
rect 14280 21836 14332 21845
rect 15568 21836 15620 21888
rect 15936 21836 15988 21888
rect 17684 21972 17736 22024
rect 18788 21972 18840 22024
rect 19524 22015 19576 22024
rect 19524 21981 19533 22015
rect 19533 21981 19567 22015
rect 19567 21981 19576 22015
rect 19524 21972 19576 21981
rect 20720 22040 20772 22092
rect 21088 22040 21140 22092
rect 22652 22040 22704 22092
rect 20904 21972 20956 22024
rect 17224 21836 17276 21888
rect 17316 21836 17368 21888
rect 21088 21904 21140 21956
rect 22744 21972 22796 22024
rect 24124 22040 24176 22092
rect 22560 21947 22612 21956
rect 22560 21913 22569 21947
rect 22569 21913 22603 21947
rect 22603 21913 22612 21947
rect 22560 21904 22612 21913
rect 23480 21972 23532 22024
rect 23572 21904 23624 21956
rect 24768 21904 24820 21956
rect 24952 21972 25004 22024
rect 25320 21904 25372 21956
rect 20352 21836 20404 21888
rect 21548 21836 21600 21888
rect 22284 21836 22336 21888
rect 22836 21836 22888 21888
rect 23020 21836 23072 21888
rect 23664 21879 23716 21888
rect 23664 21845 23673 21879
rect 23673 21845 23707 21879
rect 23707 21845 23716 21879
rect 23664 21836 23716 21845
rect 25228 21836 25280 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1308 21632 1360 21684
rect 1676 21632 1728 21684
rect 2688 21632 2740 21684
rect 4068 21632 4120 21684
rect 5448 21632 5500 21684
rect 7748 21632 7800 21684
rect 1216 21564 1268 21616
rect 1492 21564 1544 21616
rect 3700 21607 3752 21616
rect 3700 21573 3709 21607
rect 3709 21573 3743 21607
rect 3743 21573 3752 21607
rect 3700 21564 3752 21573
rect 5540 21564 5592 21616
rect 8024 21564 8076 21616
rect 10968 21632 11020 21684
rect 12716 21632 12768 21684
rect 13360 21632 13412 21684
rect 13636 21632 13688 21684
rect 13820 21675 13872 21684
rect 13820 21641 13829 21675
rect 13829 21641 13863 21675
rect 13863 21641 13872 21675
rect 13820 21632 13872 21641
rect 15384 21632 15436 21684
rect 15660 21632 15712 21684
rect 16488 21675 16540 21684
rect 16488 21641 16497 21675
rect 16497 21641 16531 21675
rect 16531 21641 16540 21675
rect 16488 21632 16540 21641
rect 16948 21632 17000 21684
rect 17132 21632 17184 21684
rect 17224 21632 17276 21684
rect 17500 21632 17552 21684
rect 17868 21632 17920 21684
rect 11428 21564 11480 21616
rect 15936 21564 15988 21616
rect 16120 21564 16172 21616
rect 2044 21539 2096 21548
rect 2044 21505 2053 21539
rect 2053 21505 2087 21539
rect 2087 21505 2096 21539
rect 2044 21496 2096 21505
rect 2228 21496 2280 21548
rect 5632 21496 5684 21548
rect 2412 21428 2464 21480
rect 6920 21471 6972 21480
rect 4068 21360 4120 21412
rect 6920 21437 6929 21471
rect 6929 21437 6963 21471
rect 6963 21437 6972 21471
rect 6920 21428 6972 21437
rect 8208 21471 8260 21480
rect 4528 21360 4580 21412
rect 5172 21360 5224 21412
rect 5540 21403 5592 21412
rect 5540 21369 5549 21403
rect 5549 21369 5583 21403
rect 5583 21369 5592 21403
rect 5540 21360 5592 21369
rect 5816 21403 5868 21412
rect 5816 21369 5825 21403
rect 5825 21369 5859 21403
rect 5859 21369 5868 21403
rect 5816 21360 5868 21369
rect 6000 21360 6052 21412
rect 7012 21360 7064 21412
rect 7196 21403 7248 21412
rect 7196 21369 7205 21403
rect 7205 21369 7239 21403
rect 7239 21369 7248 21403
rect 7196 21360 7248 21369
rect 7840 21360 7892 21412
rect 1860 21292 1912 21344
rect 2596 21335 2648 21344
rect 2596 21301 2605 21335
rect 2605 21301 2639 21335
rect 2639 21301 2648 21335
rect 2596 21292 2648 21301
rect 4160 21335 4212 21344
rect 4160 21301 4169 21335
rect 4169 21301 4203 21335
rect 4203 21301 4212 21335
rect 4160 21292 4212 21301
rect 5356 21292 5408 21344
rect 6644 21292 6696 21344
rect 8208 21437 8217 21471
rect 8217 21437 8251 21471
rect 8251 21437 8260 21471
rect 8208 21428 8260 21437
rect 10968 21496 11020 21548
rect 11980 21496 12032 21548
rect 18144 21496 18196 21548
rect 21824 21632 21876 21684
rect 22100 21632 22152 21684
rect 22652 21632 22704 21684
rect 24768 21632 24820 21684
rect 26332 21675 26384 21684
rect 26332 21641 26341 21675
rect 26341 21641 26375 21675
rect 26375 21641 26384 21675
rect 26332 21632 26384 21641
rect 22836 21564 22888 21616
rect 21824 21539 21876 21548
rect 10232 21428 10284 21480
rect 12348 21428 12400 21480
rect 12716 21471 12768 21480
rect 12716 21437 12750 21471
rect 12750 21437 12768 21471
rect 12716 21428 12768 21437
rect 13452 21428 13504 21480
rect 14832 21471 14884 21480
rect 14832 21437 14841 21471
rect 14841 21437 14875 21471
rect 14875 21437 14884 21471
rect 14832 21428 14884 21437
rect 9864 21360 9916 21412
rect 10508 21403 10560 21412
rect 10508 21369 10517 21403
rect 10517 21369 10551 21403
rect 10551 21369 10560 21403
rect 10508 21360 10560 21369
rect 11336 21403 11388 21412
rect 11336 21369 11345 21403
rect 11345 21369 11379 21403
rect 11379 21369 11388 21403
rect 11336 21360 11388 21369
rect 9496 21292 9548 21344
rect 10048 21335 10100 21344
rect 10048 21301 10057 21335
rect 10057 21301 10091 21335
rect 10091 21301 10100 21335
rect 10048 21292 10100 21301
rect 10784 21292 10836 21344
rect 11980 21292 12032 21344
rect 16580 21428 16632 21480
rect 16948 21428 17000 21480
rect 17500 21428 17552 21480
rect 18236 21428 18288 21480
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 22100 21496 22152 21548
rect 23756 21496 23808 21548
rect 24032 21496 24084 21548
rect 25044 21496 25096 21548
rect 16764 21360 16816 21412
rect 17132 21360 17184 21412
rect 19340 21428 19392 21480
rect 21548 21428 21600 21480
rect 22376 21428 22428 21480
rect 24124 21428 24176 21480
rect 25228 21471 25280 21480
rect 20904 21360 20956 21412
rect 22928 21360 22980 21412
rect 24032 21360 24084 21412
rect 25228 21437 25237 21471
rect 25237 21437 25271 21471
rect 25271 21437 25280 21471
rect 25228 21428 25280 21437
rect 26148 21428 26200 21480
rect 25504 21403 25556 21412
rect 25504 21369 25513 21403
rect 25513 21369 25547 21403
rect 25547 21369 25556 21403
rect 25504 21360 25556 21369
rect 16120 21292 16172 21344
rect 17040 21292 17092 21344
rect 19984 21292 20036 21344
rect 20352 21292 20404 21344
rect 21548 21292 21600 21344
rect 22100 21292 22152 21344
rect 22652 21292 22704 21344
rect 25320 21292 25372 21344
rect 25964 21335 26016 21344
rect 25964 21301 25973 21335
rect 25973 21301 26007 21335
rect 26007 21301 26016 21335
rect 25964 21292 26016 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1768 21088 1820 21140
rect 2044 21088 2096 21140
rect 2780 21063 2832 21072
rect 2780 21029 2789 21063
rect 2789 21029 2823 21063
rect 2823 21029 2832 21063
rect 2780 21020 2832 21029
rect 1952 20952 2004 21004
rect 2228 20952 2280 21004
rect 3332 21020 3384 21072
rect 1768 20791 1820 20800
rect 1768 20757 1777 20791
rect 1777 20757 1811 20791
rect 1811 20757 1820 20791
rect 1768 20748 1820 20757
rect 1952 20748 2004 20800
rect 3332 20884 3384 20936
rect 4988 21088 5040 21140
rect 6460 21088 6512 21140
rect 7104 21088 7156 21140
rect 7748 21088 7800 21140
rect 8024 21131 8076 21140
rect 8024 21097 8033 21131
rect 8033 21097 8067 21131
rect 8067 21097 8076 21131
rect 8024 21088 8076 21097
rect 9772 21088 9824 21140
rect 11060 21131 11112 21140
rect 11060 21097 11069 21131
rect 11069 21097 11103 21131
rect 11103 21097 11112 21131
rect 11060 21088 11112 21097
rect 12256 21088 12308 21140
rect 13912 21131 13964 21140
rect 13912 21097 13921 21131
rect 13921 21097 13955 21131
rect 13955 21097 13964 21131
rect 13912 21088 13964 21097
rect 14372 21088 14424 21140
rect 15016 21131 15068 21140
rect 15016 21097 15025 21131
rect 15025 21097 15059 21131
rect 15059 21097 15068 21131
rect 15016 21088 15068 21097
rect 15844 21131 15896 21140
rect 15844 21097 15853 21131
rect 15853 21097 15887 21131
rect 15887 21097 15896 21131
rect 15844 21088 15896 21097
rect 16764 21088 16816 21140
rect 20352 21088 20404 21140
rect 21364 21088 21416 21140
rect 22928 21088 22980 21140
rect 23204 21088 23256 21140
rect 24860 21088 24912 21140
rect 25780 21088 25832 21140
rect 5264 21020 5316 21072
rect 5448 21020 5500 21072
rect 8576 21063 8628 21072
rect 8576 21029 8585 21063
rect 8585 21029 8619 21063
rect 8619 21029 8628 21063
rect 8576 21020 8628 21029
rect 9680 21020 9732 21072
rect 14832 21020 14884 21072
rect 15752 21020 15804 21072
rect 16304 21020 16356 21072
rect 17316 21020 17368 21072
rect 17500 21063 17552 21072
rect 17500 21029 17509 21063
rect 17509 21029 17543 21063
rect 17543 21029 17552 21063
rect 17500 21020 17552 21029
rect 18972 21063 19024 21072
rect 18972 21029 18981 21063
rect 18981 21029 19015 21063
rect 19015 21029 19024 21063
rect 18972 21020 19024 21029
rect 20536 21020 20588 21072
rect 21088 21020 21140 21072
rect 21548 21063 21600 21072
rect 21548 21029 21557 21063
rect 21557 21029 21591 21063
rect 21591 21029 21600 21063
rect 21548 21020 21600 21029
rect 23756 21020 23808 21072
rect 24676 21020 24728 21072
rect 25044 21063 25096 21072
rect 25044 21029 25053 21063
rect 25053 21029 25087 21063
rect 25087 21029 25096 21063
rect 25044 21020 25096 21029
rect 4252 20952 4304 21004
rect 5816 20952 5868 21004
rect 7288 20952 7340 21004
rect 12440 20952 12492 21004
rect 13544 20952 13596 21004
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 5448 20884 5500 20936
rect 2688 20748 2740 20800
rect 3056 20748 3108 20800
rect 3332 20748 3384 20800
rect 4068 20748 4120 20800
rect 4436 20748 4488 20800
rect 6000 20884 6052 20936
rect 6644 20927 6696 20936
rect 6644 20893 6653 20927
rect 6653 20893 6687 20927
rect 6687 20893 6696 20927
rect 6644 20884 6696 20893
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 11704 20927 11756 20936
rect 9680 20884 9732 20893
rect 11704 20893 11713 20927
rect 11713 20893 11747 20927
rect 11747 20893 11756 20927
rect 11704 20884 11756 20893
rect 12256 20816 12308 20868
rect 12532 20884 12584 20936
rect 14280 20952 14332 21004
rect 19248 20952 19300 21004
rect 22836 20995 22888 21004
rect 22836 20961 22845 20995
rect 22845 20961 22879 20995
rect 22879 20961 22888 20995
rect 22836 20952 22888 20961
rect 23296 20952 23348 21004
rect 24124 20952 24176 21004
rect 6368 20748 6420 20800
rect 8944 20748 8996 20800
rect 11060 20748 11112 20800
rect 11244 20748 11296 20800
rect 12624 20791 12676 20800
rect 12624 20757 12633 20791
rect 12633 20757 12667 20791
rect 12667 20757 12676 20791
rect 12624 20748 12676 20757
rect 14648 20884 14700 20936
rect 15752 20884 15804 20936
rect 19064 20927 19116 20936
rect 19064 20893 19073 20927
rect 19073 20893 19107 20927
rect 19107 20893 19116 20927
rect 19064 20884 19116 20893
rect 21088 20884 21140 20936
rect 23112 20927 23164 20936
rect 23112 20893 23121 20927
rect 23121 20893 23155 20927
rect 23155 20893 23164 20927
rect 23112 20884 23164 20893
rect 25780 20927 25832 20936
rect 13912 20816 13964 20868
rect 16856 20816 16908 20868
rect 18788 20816 18840 20868
rect 20996 20859 21048 20868
rect 20996 20825 21005 20859
rect 21005 20825 21039 20859
rect 21039 20825 21048 20859
rect 20996 20816 21048 20825
rect 22560 20859 22612 20868
rect 22560 20825 22569 20859
rect 22569 20825 22603 20859
rect 22603 20825 22612 20859
rect 22560 20816 22612 20825
rect 23020 20816 23072 20868
rect 25780 20893 25789 20927
rect 25789 20893 25823 20927
rect 25823 20893 25832 20927
rect 25780 20884 25832 20893
rect 25044 20816 25096 20868
rect 25320 20816 25372 20868
rect 25964 20816 26016 20868
rect 14004 20748 14056 20800
rect 18512 20791 18564 20800
rect 18512 20757 18521 20791
rect 18521 20757 18555 20791
rect 18555 20757 18564 20791
rect 18512 20748 18564 20757
rect 20352 20791 20404 20800
rect 20352 20757 20361 20791
rect 20361 20757 20395 20791
rect 20395 20757 20404 20791
rect 20352 20748 20404 20757
rect 22008 20791 22060 20800
rect 22008 20757 22017 20791
rect 22017 20757 22051 20791
rect 22051 20757 22060 20791
rect 22008 20748 22060 20757
rect 22376 20791 22428 20800
rect 22376 20757 22385 20791
rect 22385 20757 22419 20791
rect 22419 20757 22428 20791
rect 22376 20748 22428 20757
rect 22836 20748 22888 20800
rect 24032 20748 24084 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2780 20544 2832 20596
rect 3056 20544 3108 20596
rect 3884 20544 3936 20596
rect 4160 20544 4212 20596
rect 5448 20544 5500 20596
rect 7656 20544 7708 20596
rect 9312 20587 9364 20596
rect 9312 20553 9321 20587
rect 9321 20553 9355 20587
rect 9355 20553 9364 20587
rect 9312 20544 9364 20553
rect 10968 20544 11020 20596
rect 12072 20544 12124 20596
rect 12440 20544 12492 20596
rect 14832 20587 14884 20596
rect 14832 20553 14841 20587
rect 14841 20553 14875 20587
rect 14875 20553 14884 20587
rect 14832 20544 14884 20553
rect 15844 20544 15896 20596
rect 16764 20587 16816 20596
rect 16764 20553 16773 20587
rect 16773 20553 16807 20587
rect 16807 20553 16816 20587
rect 16764 20544 16816 20553
rect 17684 20544 17736 20596
rect 17868 20587 17920 20596
rect 17868 20553 17877 20587
rect 17877 20553 17911 20587
rect 17911 20553 17920 20587
rect 17868 20544 17920 20553
rect 18144 20544 18196 20596
rect 19064 20544 19116 20596
rect 19524 20544 19576 20596
rect 20904 20544 20956 20596
rect 21548 20544 21600 20596
rect 21824 20544 21876 20596
rect 22100 20544 22152 20596
rect 1768 20476 1820 20528
rect 2596 20476 2648 20528
rect 1952 20408 2004 20460
rect 1124 20340 1176 20392
rect 1860 20272 1912 20324
rect 3240 20340 3292 20392
rect 4068 20476 4120 20528
rect 5356 20476 5408 20528
rect 4252 20451 4304 20460
rect 4252 20417 4261 20451
rect 4261 20417 4295 20451
rect 4295 20417 4304 20451
rect 4252 20408 4304 20417
rect 6000 20408 6052 20460
rect 6460 20408 6512 20460
rect 9680 20476 9732 20528
rect 12348 20476 12400 20528
rect 13820 20476 13872 20528
rect 8392 20408 8444 20460
rect 9956 20408 10008 20460
rect 5264 20340 5316 20392
rect 10784 20408 10836 20460
rect 11336 20451 11388 20460
rect 11336 20417 11345 20451
rect 11345 20417 11379 20451
rect 11379 20417 11388 20451
rect 11336 20408 11388 20417
rect 14740 20408 14792 20460
rect 16856 20476 16908 20528
rect 18604 20476 18656 20528
rect 18880 20519 18932 20528
rect 18880 20485 18889 20519
rect 18889 20485 18923 20519
rect 18923 20485 18932 20519
rect 18880 20476 18932 20485
rect 22468 20476 22520 20528
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 15568 20408 15620 20460
rect 16212 20408 16264 20460
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 20076 20408 20128 20460
rect 20904 20451 20956 20460
rect 20904 20417 20913 20451
rect 20913 20417 20947 20451
rect 20947 20417 20956 20451
rect 20904 20408 20956 20417
rect 22376 20408 22428 20460
rect 12440 20383 12492 20392
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 12440 20340 12492 20349
rect 12532 20340 12584 20392
rect 16856 20383 16908 20392
rect 16856 20349 16871 20383
rect 16871 20349 16905 20383
rect 16905 20349 16908 20383
rect 16856 20340 16908 20349
rect 20352 20340 20404 20392
rect 23480 20544 23532 20596
rect 5356 20272 5408 20324
rect 5908 20272 5960 20324
rect 6644 20272 6696 20324
rect 9772 20315 9824 20324
rect 9772 20281 9781 20315
rect 9781 20281 9815 20315
rect 9815 20281 9824 20315
rect 9772 20272 9824 20281
rect 11244 20272 11296 20324
rect 15476 20315 15528 20324
rect 15476 20281 15485 20315
rect 15485 20281 15519 20315
rect 15519 20281 15528 20315
rect 15476 20272 15528 20281
rect 19432 20315 19484 20324
rect 1308 20204 1360 20256
rect 1584 20204 1636 20256
rect 2136 20204 2188 20256
rect 3240 20204 3292 20256
rect 3976 20204 4028 20256
rect 4252 20204 4304 20256
rect 4988 20247 5040 20256
rect 4988 20213 4997 20247
rect 4997 20213 5031 20247
rect 5031 20213 5040 20247
rect 4988 20204 5040 20213
rect 6184 20204 6236 20256
rect 6460 20204 6512 20256
rect 8024 20204 8076 20256
rect 8392 20204 8444 20256
rect 9680 20204 9732 20256
rect 12348 20204 12400 20256
rect 13452 20204 13504 20256
rect 14372 20247 14424 20256
rect 14372 20213 14381 20247
rect 14381 20213 14415 20247
rect 14415 20213 14424 20247
rect 19432 20281 19441 20315
rect 19441 20281 19475 20315
rect 19475 20281 19484 20315
rect 19432 20272 19484 20281
rect 22100 20272 22152 20324
rect 23388 20340 23440 20392
rect 25228 20383 25280 20392
rect 25228 20349 25237 20383
rect 25237 20349 25271 20383
rect 25271 20349 25280 20383
rect 25228 20340 25280 20349
rect 24032 20315 24084 20324
rect 24032 20281 24041 20315
rect 24041 20281 24075 20315
rect 24075 20281 24084 20315
rect 24032 20272 24084 20281
rect 24124 20272 24176 20324
rect 24308 20315 24360 20324
rect 24308 20281 24317 20315
rect 24317 20281 24351 20315
rect 24351 20281 24360 20315
rect 24308 20272 24360 20281
rect 25780 20272 25832 20324
rect 14372 20204 14424 20213
rect 15752 20204 15804 20256
rect 16672 20204 16724 20256
rect 19340 20247 19392 20256
rect 19340 20213 19349 20247
rect 19349 20213 19383 20247
rect 19383 20213 19392 20247
rect 19340 20204 19392 20213
rect 19524 20204 19576 20256
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 21364 20247 21416 20256
rect 21364 20213 21373 20247
rect 21373 20213 21407 20247
rect 21407 20213 21416 20247
rect 21364 20204 21416 20213
rect 22560 20204 22612 20256
rect 23480 20247 23532 20256
rect 23480 20213 23489 20247
rect 23489 20213 23523 20247
rect 23523 20213 23532 20247
rect 23480 20204 23532 20213
rect 24676 20247 24728 20256
rect 24676 20213 24685 20247
rect 24685 20213 24719 20247
rect 24719 20213 24728 20247
rect 24676 20204 24728 20213
rect 25044 20247 25096 20256
rect 25044 20213 25053 20247
rect 25053 20213 25087 20247
rect 25087 20213 25096 20247
rect 25044 20204 25096 20213
rect 26332 20247 26384 20256
rect 26332 20213 26341 20247
rect 26341 20213 26375 20247
rect 26375 20213 26384 20247
rect 26332 20204 26384 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1952 20000 2004 20052
rect 2136 20043 2188 20052
rect 2136 20009 2145 20043
rect 2145 20009 2179 20043
rect 2179 20009 2188 20043
rect 2136 20000 2188 20009
rect 2872 20000 2924 20052
rect 3516 20000 3568 20052
rect 3792 20000 3844 20052
rect 5264 20000 5316 20052
rect 7288 20043 7340 20052
rect 7288 20009 7297 20043
rect 7297 20009 7331 20043
rect 7331 20009 7340 20043
rect 7288 20000 7340 20009
rect 8300 20043 8352 20052
rect 5172 19932 5224 19984
rect 6092 19932 6144 19984
rect 8300 20009 8309 20043
rect 8309 20009 8343 20043
rect 8343 20009 8352 20043
rect 8300 20000 8352 20009
rect 9588 20000 9640 20052
rect 12900 20000 12952 20052
rect 13452 20000 13504 20052
rect 14372 20000 14424 20052
rect 14648 20043 14700 20052
rect 14648 20009 14657 20043
rect 14657 20009 14691 20043
rect 14691 20009 14700 20043
rect 14648 20000 14700 20009
rect 15476 20000 15528 20052
rect 15752 20043 15804 20052
rect 15752 20009 15761 20043
rect 15761 20009 15795 20043
rect 15795 20009 15804 20043
rect 15752 20000 15804 20009
rect 16948 20000 17000 20052
rect 19432 20000 19484 20052
rect 24124 20000 24176 20052
rect 9680 19932 9732 19984
rect 11336 19932 11388 19984
rect 12348 19932 12400 19984
rect 15292 19975 15344 19984
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 5540 19864 5592 19916
rect 5908 19907 5960 19916
rect 5908 19873 5917 19907
rect 5917 19873 5951 19907
rect 5951 19873 5960 19907
rect 5908 19864 5960 19873
rect 3240 19796 3292 19848
rect 4988 19839 5040 19848
rect 4988 19805 4997 19839
rect 4997 19805 5031 19839
rect 5031 19805 5040 19839
rect 6460 19864 6512 19916
rect 6644 19864 6696 19916
rect 10600 19864 10652 19916
rect 12900 19864 12952 19916
rect 15292 19941 15301 19975
rect 15301 19941 15335 19975
rect 15335 19941 15344 19975
rect 15292 19932 15344 19941
rect 16488 19932 16540 19984
rect 19984 19932 20036 19984
rect 21456 19932 21508 19984
rect 21548 19932 21600 19984
rect 16396 19864 16448 19916
rect 19156 19864 19208 19916
rect 20904 19864 20956 19916
rect 21364 19907 21416 19916
rect 21364 19873 21373 19907
rect 21373 19873 21407 19907
rect 21407 19873 21416 19907
rect 21364 19864 21416 19873
rect 22100 19864 22152 19916
rect 23112 19932 23164 19984
rect 23572 19932 23624 19984
rect 22836 19864 22888 19916
rect 23296 19864 23348 19916
rect 4988 19796 5040 19805
rect 9864 19796 9916 19848
rect 10784 19796 10836 19848
rect 11612 19796 11664 19848
rect 12348 19796 12400 19848
rect 13636 19839 13688 19848
rect 13636 19805 13645 19839
rect 13645 19805 13679 19839
rect 13679 19805 13688 19839
rect 13636 19796 13688 19805
rect 15936 19796 15988 19848
rect 17868 19796 17920 19848
rect 18328 19796 18380 19848
rect 2504 19771 2556 19780
rect 2504 19737 2513 19771
rect 2513 19737 2547 19771
rect 2547 19737 2556 19771
rect 2504 19728 2556 19737
rect 5448 19728 5500 19780
rect 10876 19728 10928 19780
rect 11704 19728 11756 19780
rect 12440 19728 12492 19780
rect 13728 19728 13780 19780
rect 19248 19728 19300 19780
rect 20352 19796 20404 19848
rect 23480 19796 23532 19848
rect 24032 19796 24084 19848
rect 3884 19660 3936 19712
rect 7840 19660 7892 19712
rect 9772 19703 9824 19712
rect 9772 19669 9781 19703
rect 9781 19669 9815 19703
rect 9815 19669 9824 19703
rect 9772 19660 9824 19669
rect 10968 19660 11020 19712
rect 12256 19660 12308 19712
rect 13176 19703 13228 19712
rect 13176 19669 13185 19703
rect 13185 19669 13219 19703
rect 13219 19669 13228 19703
rect 13176 19660 13228 19669
rect 16120 19703 16172 19712
rect 16120 19669 16129 19703
rect 16129 19669 16163 19703
rect 16163 19669 16172 19703
rect 16120 19660 16172 19669
rect 18328 19703 18380 19712
rect 18328 19669 18337 19703
rect 18337 19669 18371 19703
rect 18371 19669 18380 19703
rect 18328 19660 18380 19669
rect 20076 19660 20128 19712
rect 20904 19660 20956 19712
rect 21088 19703 21140 19712
rect 21088 19669 21097 19703
rect 21097 19669 21131 19703
rect 21131 19669 21140 19703
rect 21088 19660 21140 19669
rect 23296 19728 23348 19780
rect 24308 19728 24360 19780
rect 24768 19796 24820 19848
rect 24676 19728 24728 19780
rect 25228 19771 25280 19780
rect 25228 19737 25237 19771
rect 25237 19737 25271 19771
rect 25271 19737 25280 19771
rect 25228 19728 25280 19737
rect 22744 19703 22796 19712
rect 22744 19669 22753 19703
rect 22753 19669 22787 19703
rect 22787 19669 22796 19703
rect 22744 19660 22796 19669
rect 24124 19660 24176 19712
rect 25964 19660 26016 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 4068 19456 4120 19508
rect 5264 19499 5316 19508
rect 5264 19465 5273 19499
rect 5273 19465 5307 19499
rect 5307 19465 5316 19499
rect 5264 19456 5316 19465
rect 5356 19456 5408 19508
rect 6460 19456 6512 19508
rect 7012 19499 7064 19508
rect 7012 19465 7021 19499
rect 7021 19465 7055 19499
rect 7055 19465 7064 19499
rect 7012 19456 7064 19465
rect 10600 19499 10652 19508
rect 10600 19465 10609 19499
rect 10609 19465 10643 19499
rect 10643 19465 10652 19499
rect 10600 19456 10652 19465
rect 13452 19499 13504 19508
rect 13452 19465 13461 19499
rect 13461 19465 13495 19499
rect 13495 19465 13504 19499
rect 13452 19456 13504 19465
rect 14556 19456 14608 19508
rect 15936 19456 15988 19508
rect 16212 19499 16264 19508
rect 3056 19388 3108 19440
rect 3792 19388 3844 19440
rect 4988 19320 5040 19372
rect 2412 19295 2464 19304
rect 2412 19261 2421 19295
rect 2421 19261 2455 19295
rect 2455 19261 2464 19295
rect 2412 19252 2464 19261
rect 3056 19252 3108 19304
rect 4160 19252 4212 19304
rect 6920 19388 6972 19440
rect 9496 19388 9548 19440
rect 11060 19388 11112 19440
rect 11704 19388 11756 19440
rect 11796 19388 11848 19440
rect 6092 19320 6144 19372
rect 6184 19320 6236 19372
rect 5540 19295 5592 19304
rect 2596 19227 2648 19236
rect 2228 19116 2280 19168
rect 2596 19193 2605 19227
rect 2605 19193 2639 19227
rect 2639 19193 2648 19227
rect 2596 19184 2648 19193
rect 5540 19261 5549 19295
rect 5549 19261 5583 19295
rect 5583 19261 5592 19295
rect 5540 19252 5592 19261
rect 2504 19116 2556 19168
rect 3240 19116 3292 19168
rect 4068 19116 4120 19168
rect 5172 19184 5224 19236
rect 6368 19184 6420 19236
rect 5908 19116 5960 19168
rect 9956 19252 10008 19304
rect 11796 19252 11848 19304
rect 6644 19227 6696 19236
rect 6644 19193 6653 19227
rect 6653 19193 6687 19227
rect 6687 19193 6696 19227
rect 6644 19184 6696 19193
rect 7656 19116 7708 19168
rect 8392 19184 8444 19236
rect 10876 19227 10928 19236
rect 10876 19193 10885 19227
rect 10885 19193 10919 19227
rect 10919 19193 10928 19227
rect 10876 19184 10928 19193
rect 12900 19388 12952 19440
rect 14648 19388 14700 19440
rect 15384 19388 15436 19440
rect 16212 19465 16221 19499
rect 16221 19465 16255 19499
rect 16255 19465 16264 19499
rect 16212 19456 16264 19465
rect 19432 19456 19484 19508
rect 12256 19320 12308 19372
rect 16120 19320 16172 19372
rect 19340 19320 19392 19372
rect 19616 19320 19668 19372
rect 21364 19456 21416 19508
rect 22100 19499 22152 19508
rect 22100 19465 22109 19499
rect 22109 19465 22143 19499
rect 22143 19465 22152 19499
rect 22100 19456 22152 19465
rect 23756 19499 23808 19508
rect 23756 19465 23765 19499
rect 23765 19465 23799 19499
rect 23799 19465 23808 19499
rect 23756 19456 23808 19465
rect 24768 19456 24820 19508
rect 22744 19388 22796 19440
rect 12716 19252 12768 19304
rect 12900 19252 12952 19304
rect 14372 19252 14424 19304
rect 15936 19252 15988 19304
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 23572 19320 23624 19372
rect 23848 19320 23900 19372
rect 24032 19320 24084 19372
rect 24308 19320 24360 19372
rect 24492 19320 24544 19372
rect 25044 19388 25096 19440
rect 21456 19252 21508 19304
rect 23020 19252 23072 19304
rect 25228 19295 25280 19304
rect 25228 19261 25237 19295
rect 25237 19261 25271 19295
rect 25271 19261 25280 19295
rect 25228 19252 25280 19261
rect 13728 19184 13780 19236
rect 14556 19184 14608 19236
rect 18328 19184 18380 19236
rect 19432 19184 19484 19236
rect 23112 19184 23164 19236
rect 23848 19184 23900 19236
rect 24032 19227 24084 19236
rect 24032 19193 24041 19227
rect 24041 19193 24075 19227
rect 24075 19193 24084 19227
rect 24032 19184 24084 19193
rect 24216 19227 24268 19236
rect 24216 19193 24225 19227
rect 24225 19193 24259 19227
rect 24259 19193 24268 19227
rect 24216 19184 24268 19193
rect 24676 19227 24728 19236
rect 10784 19116 10836 19168
rect 11060 19159 11112 19168
rect 11060 19125 11069 19159
rect 11069 19125 11103 19159
rect 11103 19125 11112 19159
rect 11060 19116 11112 19125
rect 11244 19116 11296 19168
rect 11336 19116 11388 19168
rect 11612 19116 11664 19168
rect 12808 19116 12860 19168
rect 13636 19116 13688 19168
rect 14004 19116 14056 19168
rect 15200 19116 15252 19168
rect 16856 19116 16908 19168
rect 20076 19116 20128 19168
rect 23480 19159 23532 19168
rect 23480 19125 23489 19159
rect 23489 19125 23523 19159
rect 23523 19125 23532 19159
rect 23480 19116 23532 19125
rect 23664 19116 23716 19168
rect 24676 19193 24685 19227
rect 24685 19193 24719 19227
rect 24719 19193 24728 19227
rect 24676 19184 24728 19193
rect 25412 19159 25464 19168
rect 25412 19125 25421 19159
rect 25421 19125 25455 19159
rect 25455 19125 25464 19159
rect 25412 19116 25464 19125
rect 26332 19116 26384 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1400 18912 1452 18964
rect 3884 18912 3936 18964
rect 4988 18912 5040 18964
rect 6000 18955 6052 18964
rect 6000 18921 6009 18955
rect 6009 18921 6043 18955
rect 6043 18921 6052 18955
rect 6000 18912 6052 18921
rect 2872 18844 2924 18896
rect 3056 18844 3108 18896
rect 4068 18844 4120 18896
rect 5264 18887 5316 18896
rect 5264 18853 5273 18887
rect 5273 18853 5307 18887
rect 5307 18853 5316 18887
rect 5264 18844 5316 18853
rect 5448 18887 5500 18896
rect 5448 18853 5457 18887
rect 5457 18853 5491 18887
rect 5491 18853 5500 18887
rect 5448 18844 5500 18853
rect 6276 18844 6328 18896
rect 6460 18844 6512 18896
rect 7288 18844 7340 18896
rect 8116 18844 8168 18896
rect 8576 18887 8628 18896
rect 8576 18853 8585 18887
rect 8585 18853 8619 18887
rect 8619 18853 8628 18887
rect 8576 18844 8628 18853
rect 4436 18776 4488 18828
rect 4988 18776 5040 18828
rect 2044 18708 2096 18760
rect 2872 18751 2924 18760
rect 2872 18717 2881 18751
rect 2881 18717 2915 18751
rect 2915 18717 2924 18751
rect 2872 18708 2924 18717
rect 3424 18708 3476 18760
rect 5908 18776 5960 18828
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 7196 18776 7248 18828
rect 4436 18572 4488 18624
rect 4804 18640 4856 18692
rect 6276 18640 6328 18692
rect 7472 18708 7524 18760
rect 8484 18751 8536 18760
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 9588 18912 9640 18964
rect 11796 18955 11848 18964
rect 11796 18921 11805 18955
rect 11805 18921 11839 18955
rect 11839 18921 11848 18955
rect 11796 18912 11848 18921
rect 13728 18912 13780 18964
rect 16488 18912 16540 18964
rect 18144 18955 18196 18964
rect 18144 18921 18153 18955
rect 18153 18921 18187 18955
rect 18187 18921 18196 18955
rect 18144 18912 18196 18921
rect 10876 18844 10928 18896
rect 13452 18887 13504 18896
rect 13452 18853 13461 18887
rect 13461 18853 13495 18887
rect 13495 18853 13504 18887
rect 13452 18844 13504 18853
rect 16212 18844 16264 18896
rect 17408 18887 17460 18896
rect 17408 18853 17417 18887
rect 17417 18853 17451 18887
rect 17451 18853 17460 18887
rect 17408 18844 17460 18853
rect 18972 18887 19024 18896
rect 18972 18853 18981 18887
rect 18981 18853 19015 18887
rect 19015 18853 19024 18887
rect 18972 18844 19024 18853
rect 19432 18912 19484 18964
rect 19984 18912 20036 18964
rect 21548 18912 21600 18964
rect 22100 18912 22152 18964
rect 24032 18912 24084 18964
rect 19524 18844 19576 18896
rect 20076 18844 20128 18896
rect 11796 18776 11848 18828
rect 12256 18776 12308 18828
rect 15108 18819 15160 18828
rect 15108 18785 15117 18819
rect 15117 18785 15151 18819
rect 15151 18785 15160 18819
rect 15108 18776 15160 18785
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 15936 18819 15988 18828
rect 15936 18785 15945 18819
rect 15945 18785 15979 18819
rect 15979 18785 15988 18819
rect 15936 18776 15988 18785
rect 18512 18776 18564 18828
rect 20536 18844 20588 18896
rect 21456 18887 21508 18896
rect 21456 18853 21465 18887
rect 21465 18853 21499 18887
rect 21499 18853 21508 18887
rect 21456 18844 21508 18853
rect 22284 18844 22336 18896
rect 22744 18844 22796 18896
rect 23020 18887 23072 18896
rect 23020 18853 23029 18887
rect 23029 18853 23063 18887
rect 23063 18853 23072 18887
rect 23020 18844 23072 18853
rect 24676 18844 24728 18896
rect 25044 18887 25096 18896
rect 25044 18853 25053 18887
rect 25053 18853 25087 18887
rect 25087 18853 25096 18887
rect 25044 18844 25096 18853
rect 22376 18776 22428 18828
rect 9496 18708 9548 18760
rect 9772 18708 9824 18760
rect 10140 18708 10192 18760
rect 10232 18708 10284 18760
rect 13912 18708 13964 18760
rect 17316 18751 17368 18760
rect 17316 18717 17325 18751
rect 17325 18717 17359 18751
rect 17359 18717 17368 18751
rect 17316 18708 17368 18717
rect 17776 18708 17828 18760
rect 20904 18708 20956 18760
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 22008 18708 22060 18760
rect 24216 18708 24268 18760
rect 12900 18640 12952 18692
rect 15384 18683 15436 18692
rect 6644 18572 6696 18624
rect 7472 18615 7524 18624
rect 7472 18581 7481 18615
rect 7481 18581 7515 18615
rect 7515 18581 7524 18615
rect 7472 18572 7524 18581
rect 7840 18615 7892 18624
rect 7840 18581 7849 18615
rect 7849 18581 7883 18615
rect 7883 18581 7892 18615
rect 7840 18572 7892 18581
rect 9956 18615 10008 18624
rect 9956 18581 9965 18615
rect 9965 18581 9999 18615
rect 9999 18581 10008 18615
rect 9956 18572 10008 18581
rect 10140 18572 10192 18624
rect 12256 18572 12308 18624
rect 12440 18615 12492 18624
rect 12440 18581 12449 18615
rect 12449 18581 12483 18615
rect 12483 18581 12492 18615
rect 12440 18572 12492 18581
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 13728 18572 13780 18624
rect 14004 18572 14056 18624
rect 15384 18649 15393 18683
rect 15393 18649 15427 18683
rect 15427 18649 15436 18683
rect 15384 18640 15436 18649
rect 16948 18683 17000 18692
rect 16948 18649 16957 18683
rect 16957 18649 16991 18683
rect 16991 18649 17000 18683
rect 16948 18640 17000 18649
rect 19248 18640 19300 18692
rect 20996 18683 21048 18692
rect 20996 18649 21005 18683
rect 21005 18649 21039 18683
rect 21039 18649 21048 18683
rect 20996 18640 21048 18649
rect 22836 18640 22888 18692
rect 24032 18640 24084 18692
rect 24308 18640 24360 18692
rect 24400 18640 24452 18692
rect 24860 18708 24912 18760
rect 25044 18708 25096 18760
rect 26424 18640 26476 18692
rect 15476 18572 15528 18624
rect 19984 18572 20036 18624
rect 20352 18572 20404 18624
rect 22376 18615 22428 18624
rect 22376 18581 22385 18615
rect 22385 18581 22419 18615
rect 22419 18581 22428 18615
rect 22376 18572 22428 18581
rect 23664 18615 23716 18624
rect 23664 18581 23673 18615
rect 23673 18581 23707 18615
rect 23707 18581 23716 18615
rect 23664 18572 23716 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 3056 18368 3108 18420
rect 3792 18411 3844 18420
rect 3792 18377 3801 18411
rect 3801 18377 3835 18411
rect 3835 18377 3844 18411
rect 3792 18368 3844 18377
rect 2780 18343 2832 18352
rect 2780 18309 2789 18343
rect 2789 18309 2823 18343
rect 2823 18309 2832 18343
rect 2780 18300 2832 18309
rect 1584 18232 1636 18284
rect 3240 18275 3292 18284
rect 3240 18241 3249 18275
rect 3249 18241 3283 18275
rect 3283 18241 3292 18275
rect 3240 18232 3292 18241
rect 5172 18368 5224 18420
rect 6460 18368 6512 18420
rect 8116 18411 8168 18420
rect 8116 18377 8125 18411
rect 8125 18377 8159 18411
rect 8159 18377 8168 18411
rect 8116 18368 8168 18377
rect 8300 18368 8352 18420
rect 5448 18300 5500 18352
rect 5264 18232 5316 18284
rect 7656 18300 7708 18352
rect 7472 18275 7524 18284
rect 7472 18241 7481 18275
rect 7481 18241 7515 18275
rect 7515 18241 7524 18275
rect 7472 18232 7524 18241
rect 10232 18368 10284 18420
rect 11060 18368 11112 18420
rect 13452 18411 13504 18420
rect 13452 18377 13461 18411
rect 13461 18377 13495 18411
rect 13495 18377 13504 18411
rect 13452 18368 13504 18377
rect 10876 18300 10928 18352
rect 12624 18300 12676 18352
rect 13084 18300 13136 18352
rect 14556 18368 14608 18420
rect 15292 18368 15344 18420
rect 15936 18368 15988 18420
rect 17040 18411 17092 18420
rect 17040 18377 17049 18411
rect 17049 18377 17083 18411
rect 17083 18377 17092 18411
rect 17040 18368 17092 18377
rect 18972 18368 19024 18420
rect 19432 18411 19484 18420
rect 19432 18377 19441 18411
rect 19441 18377 19475 18411
rect 19475 18377 19484 18411
rect 19432 18368 19484 18377
rect 21364 18411 21416 18420
rect 18144 18343 18196 18352
rect 18144 18309 18153 18343
rect 18153 18309 18187 18343
rect 18187 18309 18196 18343
rect 18144 18300 18196 18309
rect 18696 18300 18748 18352
rect 21364 18377 21373 18411
rect 21373 18377 21407 18411
rect 21407 18377 21416 18411
rect 21364 18368 21416 18377
rect 21456 18368 21508 18420
rect 22008 18368 22060 18420
rect 22652 18411 22704 18420
rect 22652 18377 22661 18411
rect 22661 18377 22695 18411
rect 22695 18377 22704 18411
rect 22652 18368 22704 18377
rect 23664 18368 23716 18420
rect 24216 18368 24268 18420
rect 25044 18411 25096 18420
rect 25044 18377 25053 18411
rect 25053 18377 25087 18411
rect 25087 18377 25096 18411
rect 25044 18368 25096 18377
rect 25596 18368 25648 18420
rect 25780 18411 25832 18420
rect 25780 18377 25789 18411
rect 25789 18377 25823 18411
rect 25823 18377 25832 18411
rect 25780 18368 25832 18377
rect 26240 18343 26292 18352
rect 26240 18309 26249 18343
rect 26249 18309 26283 18343
rect 26283 18309 26292 18343
rect 26240 18300 26292 18309
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 6368 18164 6420 18216
rect 1584 18096 1636 18148
rect 3056 18096 3108 18148
rect 3608 18028 3660 18080
rect 4436 18028 4488 18080
rect 5448 18096 5500 18148
rect 6828 18096 6880 18148
rect 7380 18139 7432 18148
rect 7380 18105 7389 18139
rect 7389 18105 7423 18139
rect 7423 18105 7432 18139
rect 7380 18096 7432 18105
rect 5540 18028 5592 18080
rect 9312 18028 9364 18080
rect 9496 18028 9548 18080
rect 9588 18028 9640 18080
rect 11060 18232 11112 18284
rect 11428 18232 11480 18284
rect 13360 18232 13412 18284
rect 14280 18275 14332 18284
rect 14280 18241 14289 18275
rect 14289 18241 14323 18275
rect 14323 18241 14332 18275
rect 14280 18232 14332 18241
rect 16120 18232 16172 18284
rect 16304 18232 16356 18284
rect 17408 18232 17460 18284
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 23848 18232 23900 18284
rect 24860 18232 24912 18284
rect 10600 18164 10652 18216
rect 10876 18164 10928 18216
rect 9956 18096 10008 18148
rect 10692 18096 10744 18148
rect 14556 18139 14608 18148
rect 14556 18105 14590 18139
rect 14590 18105 14608 18139
rect 14556 18096 14608 18105
rect 10784 18028 10836 18080
rect 11152 18028 11204 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 15384 18028 15436 18080
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 18236 18164 18288 18216
rect 17408 18071 17460 18080
rect 17408 18037 17417 18071
rect 17417 18037 17451 18071
rect 17451 18037 17460 18071
rect 17408 18028 17460 18037
rect 18788 18028 18840 18080
rect 20076 18164 20128 18216
rect 22376 18164 22428 18216
rect 24032 18207 24084 18216
rect 24032 18173 24041 18207
rect 24041 18173 24075 18207
rect 24075 18173 24084 18207
rect 24032 18164 24084 18173
rect 25044 18164 25096 18216
rect 25780 18164 25832 18216
rect 20904 18096 20956 18148
rect 21548 18096 21600 18148
rect 22100 18096 22152 18148
rect 23020 18139 23072 18148
rect 23020 18105 23029 18139
rect 23029 18105 23063 18139
rect 23063 18105 23072 18139
rect 23020 18096 23072 18105
rect 24124 18096 24176 18148
rect 22192 18071 22244 18080
rect 22192 18037 22201 18071
rect 22201 18037 22235 18071
rect 22235 18037 22244 18071
rect 22192 18028 22244 18037
rect 23848 18028 23900 18080
rect 24676 18071 24728 18080
rect 24676 18037 24685 18071
rect 24685 18037 24719 18071
rect 24719 18037 24728 18071
rect 24676 18028 24728 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2688 17824 2740 17876
rect 2780 17824 2832 17876
rect 3516 17867 3568 17876
rect 3516 17833 3525 17867
rect 3525 17833 3559 17867
rect 3559 17833 3568 17867
rect 3516 17824 3568 17833
rect 3608 17824 3660 17876
rect 2596 17756 2648 17808
rect 2872 17756 2924 17808
rect 2688 17688 2740 17740
rect 6828 17824 6880 17876
rect 7104 17824 7156 17876
rect 7380 17824 7432 17876
rect 8484 17867 8536 17876
rect 8484 17833 8493 17867
rect 8493 17833 8527 17867
rect 8527 17833 8536 17867
rect 8484 17824 8536 17833
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 3608 17620 3660 17672
rect 4436 17620 4488 17672
rect 4712 17620 4764 17672
rect 5172 17756 5224 17808
rect 6184 17756 6236 17808
rect 5540 17688 5592 17740
rect 7012 17688 7064 17740
rect 7564 17688 7616 17740
rect 7748 17688 7800 17740
rect 10324 17799 10376 17808
rect 10324 17765 10333 17799
rect 10333 17765 10367 17799
rect 10367 17765 10376 17799
rect 10324 17756 10376 17765
rect 12072 17756 12124 17808
rect 9404 17688 9456 17740
rect 9864 17688 9916 17740
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 3700 17552 3752 17604
rect 6000 17552 6052 17604
rect 8116 17663 8168 17672
rect 8116 17629 8125 17663
rect 8125 17629 8159 17663
rect 8159 17629 8168 17663
rect 8116 17620 8168 17629
rect 8944 17620 8996 17672
rect 9588 17620 9640 17672
rect 2136 17484 2188 17536
rect 4712 17484 4764 17536
rect 6184 17484 6236 17536
rect 8208 17552 8260 17604
rect 7656 17484 7708 17536
rect 9680 17552 9732 17604
rect 9588 17484 9640 17536
rect 10692 17620 10744 17672
rect 11060 17552 11112 17604
rect 10784 17527 10836 17536
rect 10784 17493 10793 17527
rect 10793 17493 10827 17527
rect 10827 17493 10836 17527
rect 10784 17484 10836 17493
rect 10968 17484 11020 17536
rect 11796 17688 11848 17740
rect 12900 17824 12952 17876
rect 13360 17824 13412 17876
rect 13544 17824 13596 17876
rect 15108 17867 15160 17876
rect 15108 17833 15117 17867
rect 15117 17833 15151 17867
rect 15151 17833 15160 17867
rect 15108 17824 15160 17833
rect 16028 17824 16080 17876
rect 18052 17867 18104 17876
rect 18052 17833 18061 17867
rect 18061 17833 18095 17867
rect 18095 17833 18104 17867
rect 18052 17824 18104 17833
rect 18512 17824 18564 17876
rect 20904 17824 20956 17876
rect 12808 17756 12860 17808
rect 13268 17799 13320 17808
rect 13268 17765 13277 17799
rect 13277 17765 13311 17799
rect 13311 17765 13320 17799
rect 13268 17756 13320 17765
rect 14280 17688 14332 17740
rect 14556 17688 14608 17740
rect 17868 17756 17920 17808
rect 19800 17799 19852 17808
rect 19800 17765 19809 17799
rect 19809 17765 19843 17799
rect 19843 17765 19852 17799
rect 19800 17756 19852 17765
rect 20812 17756 20864 17808
rect 22284 17867 22336 17876
rect 22284 17833 22293 17867
rect 22293 17833 22327 17867
rect 22327 17833 22336 17867
rect 22284 17824 22336 17833
rect 23664 17867 23716 17876
rect 23664 17833 23673 17867
rect 23673 17833 23707 17867
rect 23707 17833 23716 17867
rect 23664 17824 23716 17833
rect 23756 17824 23808 17876
rect 16212 17688 16264 17740
rect 16580 17688 16632 17740
rect 17224 17688 17276 17740
rect 19432 17688 19484 17740
rect 20444 17688 20496 17740
rect 21548 17756 21600 17808
rect 22836 17799 22888 17808
rect 22836 17765 22845 17799
rect 22845 17765 22879 17799
rect 22879 17765 22888 17799
rect 22836 17756 22888 17765
rect 23112 17756 23164 17808
rect 24860 17824 24912 17876
rect 24400 17731 24452 17740
rect 24400 17697 24409 17731
rect 24409 17697 24443 17731
rect 24443 17697 24452 17731
rect 24400 17688 24452 17697
rect 24860 17688 24912 17740
rect 25044 17688 25096 17740
rect 13452 17620 13504 17672
rect 12164 17552 12216 17604
rect 12992 17527 13044 17536
rect 12992 17493 13001 17527
rect 13001 17493 13035 17527
rect 13035 17493 13044 17527
rect 12992 17484 13044 17493
rect 14188 17484 14240 17536
rect 15660 17620 15712 17672
rect 15936 17552 15988 17604
rect 18880 17620 18932 17672
rect 20904 17620 20956 17672
rect 21180 17620 21232 17672
rect 21548 17663 21600 17672
rect 21548 17629 21557 17663
rect 21557 17629 21591 17663
rect 21591 17629 21600 17663
rect 21548 17620 21600 17629
rect 24676 17663 24728 17672
rect 14648 17527 14700 17536
rect 14648 17493 14657 17527
rect 14657 17493 14691 17527
rect 14691 17493 14700 17527
rect 14648 17484 14700 17493
rect 16580 17527 16632 17536
rect 16580 17493 16589 17527
rect 16589 17493 16623 17527
rect 16623 17493 16632 17527
rect 16580 17484 16632 17493
rect 19616 17552 19668 17604
rect 21088 17552 21140 17604
rect 24676 17629 24685 17663
rect 24685 17629 24719 17663
rect 24719 17629 24728 17663
rect 24676 17620 24728 17629
rect 24124 17595 24176 17604
rect 24124 17561 24133 17595
rect 24133 17561 24167 17595
rect 24167 17561 24176 17595
rect 24124 17552 24176 17561
rect 18972 17484 19024 17536
rect 20536 17484 20588 17536
rect 20720 17484 20772 17536
rect 22560 17527 22612 17536
rect 22560 17493 22569 17527
rect 22569 17493 22603 17527
rect 22603 17493 22612 17527
rect 22560 17484 22612 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2412 17280 2464 17332
rect 3608 17280 3660 17332
rect 4344 17323 4396 17332
rect 4344 17289 4353 17323
rect 4353 17289 4387 17323
rect 4387 17289 4396 17323
rect 4344 17280 4396 17289
rect 5172 17280 5224 17332
rect 6920 17323 6972 17332
rect 6920 17289 6929 17323
rect 6929 17289 6963 17323
rect 6963 17289 6972 17323
rect 6920 17280 6972 17289
rect 7012 17280 7064 17332
rect 7932 17280 7984 17332
rect 3240 17212 3292 17264
rect 3884 17144 3936 17196
rect 1768 17076 1820 17128
rect 2872 17076 2924 17128
rect 3516 17076 3568 17128
rect 2780 17008 2832 17060
rect 3056 17051 3108 17060
rect 3056 17017 3065 17051
rect 3065 17017 3099 17051
rect 3099 17017 3108 17051
rect 3056 17008 3108 17017
rect 3608 17008 3660 17060
rect 5632 17212 5684 17264
rect 7196 17212 7248 17264
rect 8944 17280 8996 17332
rect 12532 17323 12584 17332
rect 12532 17289 12541 17323
rect 12541 17289 12575 17323
rect 12575 17289 12584 17323
rect 12532 17280 12584 17289
rect 13544 17323 13596 17332
rect 13544 17289 13553 17323
rect 13553 17289 13587 17323
rect 13587 17289 13596 17323
rect 13544 17280 13596 17289
rect 14188 17280 14240 17332
rect 14372 17280 14424 17332
rect 14832 17280 14884 17332
rect 16212 17323 16264 17332
rect 16212 17289 16221 17323
rect 16221 17289 16255 17323
rect 16255 17289 16264 17323
rect 16212 17280 16264 17289
rect 17592 17280 17644 17332
rect 4804 17187 4856 17196
rect 4804 17153 4813 17187
rect 4813 17153 4847 17187
rect 4847 17153 4856 17187
rect 4804 17144 4856 17153
rect 5448 17144 5500 17196
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 10968 17212 11020 17264
rect 12164 17255 12216 17264
rect 12164 17221 12173 17255
rect 12173 17221 12207 17255
rect 12207 17221 12216 17255
rect 12164 17212 12216 17221
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 12072 17187 12124 17196
rect 12072 17153 12081 17187
rect 12081 17153 12115 17187
rect 12115 17153 12124 17187
rect 12072 17144 12124 17153
rect 12716 17144 12768 17196
rect 13176 17144 13228 17196
rect 15936 17212 15988 17264
rect 17224 17212 17276 17264
rect 17868 17212 17920 17264
rect 19800 17280 19852 17332
rect 20720 17280 20772 17332
rect 20812 17280 20864 17332
rect 21272 17280 21324 17332
rect 18788 17187 18840 17196
rect 4712 17076 4764 17128
rect 9956 17076 10008 17128
rect 4804 17051 4856 17060
rect 4804 17017 4813 17051
rect 4813 17017 4847 17051
rect 4847 17017 4856 17051
rect 4804 17008 4856 17017
rect 6920 17008 6972 17060
rect 7380 17051 7432 17060
rect 7380 17017 7389 17051
rect 7389 17017 7423 17051
rect 7423 17017 7432 17051
rect 7380 17008 7432 17017
rect 8116 17008 8168 17060
rect 9128 17008 9180 17060
rect 12348 17008 12400 17060
rect 12440 17008 12492 17060
rect 12992 17051 13044 17060
rect 12992 17017 13001 17051
rect 13001 17017 13035 17051
rect 13035 17017 13044 17051
rect 12992 17008 13044 17017
rect 13084 17051 13136 17060
rect 13084 17017 13093 17051
rect 13093 17017 13127 17051
rect 13127 17017 13136 17051
rect 13084 17008 13136 17017
rect 13544 17008 13596 17060
rect 16672 17076 16724 17128
rect 17040 17076 17092 17128
rect 18788 17153 18797 17187
rect 18797 17153 18831 17187
rect 18831 17153 18840 17187
rect 18788 17144 18840 17153
rect 19524 17187 19576 17196
rect 19524 17153 19533 17187
rect 19533 17153 19567 17187
rect 19567 17153 19576 17187
rect 19524 17144 19576 17153
rect 19616 17187 19668 17196
rect 19616 17153 19625 17187
rect 19625 17153 19659 17187
rect 19659 17153 19668 17187
rect 19616 17144 19668 17153
rect 20352 17144 20404 17196
rect 14372 17008 14424 17060
rect 16948 17008 17000 17060
rect 19892 17076 19944 17128
rect 3700 16983 3752 16992
rect 3700 16949 3709 16983
rect 3709 16949 3743 16983
rect 3743 16949 3752 16983
rect 3700 16940 3752 16949
rect 4252 16940 4304 16992
rect 4712 16940 4764 16992
rect 5540 16940 5592 16992
rect 11060 16940 11112 16992
rect 11244 16940 11296 16992
rect 14188 16940 14240 16992
rect 17776 16940 17828 16992
rect 18236 16940 18288 16992
rect 19248 16940 19300 16992
rect 19984 16940 20036 16992
rect 20536 17212 20588 17264
rect 20996 17212 21048 17264
rect 22560 17280 22612 17332
rect 22836 17280 22888 17332
rect 23756 17323 23808 17332
rect 23756 17289 23765 17323
rect 23765 17289 23799 17323
rect 23799 17289 23808 17323
rect 23756 17280 23808 17289
rect 25688 17280 25740 17332
rect 22192 17212 22244 17264
rect 24676 17255 24728 17264
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 22376 17144 22428 17196
rect 21180 17119 21232 17128
rect 21180 17085 21189 17119
rect 21189 17085 21223 17119
rect 21223 17085 21232 17119
rect 21180 17076 21232 17085
rect 21456 17076 21508 17128
rect 22284 17119 22336 17128
rect 22284 17085 22293 17119
rect 22293 17085 22327 17119
rect 22327 17085 22336 17119
rect 22284 17076 22336 17085
rect 24676 17221 24685 17255
rect 24685 17221 24719 17255
rect 24719 17221 24728 17255
rect 24676 17212 24728 17221
rect 25320 17212 25372 17264
rect 25872 17212 25924 17264
rect 23664 17144 23716 17196
rect 20536 16940 20588 16992
rect 21548 16983 21600 16992
rect 21548 16949 21557 16983
rect 21557 16949 21591 16983
rect 21591 16949 21600 16983
rect 24676 17008 24728 17060
rect 21548 16940 21600 16949
rect 23020 16940 23072 16992
rect 24216 16983 24268 16992
rect 24216 16949 24225 16983
rect 24225 16949 24259 16983
rect 24259 16949 24268 16983
rect 24216 16940 24268 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2412 16736 2464 16788
rect 3056 16736 3108 16788
rect 3424 16779 3476 16788
rect 3424 16745 3433 16779
rect 3433 16745 3467 16779
rect 3467 16745 3476 16779
rect 3424 16736 3476 16745
rect 3884 16779 3936 16788
rect 3884 16745 3893 16779
rect 3893 16745 3927 16779
rect 3927 16745 3936 16779
rect 5448 16779 5500 16788
rect 3884 16736 3936 16745
rect 2596 16668 2648 16720
rect 3976 16668 4028 16720
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 9864 16779 9916 16788
rect 6000 16668 6052 16720
rect 6184 16668 6236 16720
rect 9864 16745 9873 16779
rect 9873 16745 9907 16779
rect 9907 16745 9916 16779
rect 9864 16736 9916 16745
rect 10692 16779 10744 16788
rect 10692 16745 10701 16779
rect 10701 16745 10735 16779
rect 10735 16745 10744 16779
rect 10692 16736 10744 16745
rect 11060 16736 11112 16788
rect 13084 16736 13136 16788
rect 13176 16736 13228 16788
rect 14648 16736 14700 16788
rect 15016 16779 15068 16788
rect 15016 16745 15025 16779
rect 15025 16745 15059 16779
rect 15059 16745 15068 16779
rect 15844 16779 15896 16788
rect 15016 16736 15068 16745
rect 8852 16668 8904 16720
rect 1768 16600 1820 16652
rect 2504 16532 2556 16584
rect 4344 16643 4396 16652
rect 4344 16609 4378 16643
rect 4378 16609 4396 16643
rect 4344 16600 4396 16609
rect 6828 16600 6880 16652
rect 7196 16600 7248 16652
rect 8208 16600 8260 16652
rect 10232 16600 10284 16652
rect 2136 16464 2188 16516
rect 2688 16464 2740 16516
rect 1952 16439 2004 16448
rect 1952 16405 1961 16439
rect 1961 16405 1995 16439
rect 1995 16405 2004 16439
rect 1952 16396 2004 16405
rect 2872 16396 2924 16448
rect 9864 16532 9916 16584
rect 4252 16396 4304 16448
rect 5172 16396 5224 16448
rect 6000 16439 6052 16448
rect 6000 16405 6009 16439
rect 6009 16405 6043 16439
rect 6043 16405 6052 16439
rect 6000 16396 6052 16405
rect 10968 16668 11020 16720
rect 13452 16711 13504 16720
rect 13452 16677 13461 16711
rect 13461 16677 13495 16711
rect 13495 16677 13504 16711
rect 13452 16668 13504 16677
rect 13820 16668 13872 16720
rect 15844 16745 15853 16779
rect 15853 16745 15887 16779
rect 15887 16745 15896 16779
rect 15844 16736 15896 16745
rect 18420 16736 18472 16788
rect 19432 16779 19484 16788
rect 19432 16745 19441 16779
rect 19441 16745 19475 16779
rect 19475 16745 19484 16779
rect 19432 16736 19484 16745
rect 20536 16779 20588 16788
rect 20536 16745 20545 16779
rect 20545 16745 20579 16779
rect 20579 16745 20588 16779
rect 20536 16736 20588 16745
rect 17224 16668 17276 16720
rect 18052 16668 18104 16720
rect 20444 16668 20496 16720
rect 12716 16600 12768 16652
rect 10784 16532 10836 16584
rect 10876 16396 10928 16448
rect 13084 16532 13136 16584
rect 13636 16532 13688 16584
rect 14924 16600 14976 16652
rect 14096 16464 14148 16516
rect 16488 16600 16540 16652
rect 17316 16600 17368 16652
rect 18328 16600 18380 16652
rect 19984 16600 20036 16652
rect 21180 16736 21232 16788
rect 22008 16736 22060 16788
rect 22284 16736 22336 16788
rect 23940 16779 23992 16788
rect 23940 16745 23949 16779
rect 23949 16745 23983 16779
rect 23983 16745 23992 16779
rect 23940 16736 23992 16745
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 25136 16779 25188 16788
rect 25136 16745 25145 16779
rect 25145 16745 25179 16779
rect 25179 16745 25188 16779
rect 25136 16736 25188 16745
rect 20996 16668 21048 16720
rect 21548 16668 21600 16720
rect 22376 16668 22428 16720
rect 23388 16668 23440 16720
rect 21180 16643 21232 16652
rect 21180 16609 21214 16643
rect 21214 16609 21232 16643
rect 21180 16600 21232 16609
rect 22560 16600 22612 16652
rect 24952 16643 25004 16652
rect 24952 16609 24961 16643
rect 24961 16609 24995 16643
rect 24995 16609 25004 16643
rect 24952 16600 25004 16609
rect 16396 16532 16448 16584
rect 20444 16532 20496 16584
rect 22836 16532 22888 16584
rect 23296 16532 23348 16584
rect 15660 16464 15712 16516
rect 19524 16464 19576 16516
rect 20536 16464 20588 16516
rect 24216 16464 24268 16516
rect 11428 16396 11480 16448
rect 14372 16396 14424 16448
rect 16028 16396 16080 16448
rect 21180 16396 21232 16448
rect 23204 16439 23256 16448
rect 23204 16405 23213 16439
rect 23213 16405 23247 16439
rect 23247 16405 23256 16439
rect 23204 16396 23256 16405
rect 23296 16396 23348 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1676 16192 1728 16244
rect 2504 16235 2556 16244
rect 2504 16201 2513 16235
rect 2513 16201 2547 16235
rect 2547 16201 2556 16235
rect 2504 16192 2556 16201
rect 4252 16192 4304 16244
rect 4804 16192 4856 16244
rect 6184 16192 6236 16244
rect 9128 16235 9180 16244
rect 9128 16201 9137 16235
rect 9137 16201 9171 16235
rect 9171 16201 9180 16235
rect 9128 16192 9180 16201
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 13084 16192 13136 16244
rect 13820 16192 13872 16244
rect 14188 16192 14240 16244
rect 14372 16192 14424 16244
rect 16028 16235 16080 16244
rect 2596 16124 2648 16176
rect 8760 16124 8812 16176
rect 12532 16167 12584 16176
rect 12532 16133 12541 16167
rect 12541 16133 12575 16167
rect 12575 16133 12584 16167
rect 12532 16124 12584 16133
rect 16028 16201 16037 16235
rect 16037 16201 16071 16235
rect 16071 16201 16080 16235
rect 16028 16192 16080 16201
rect 17224 16235 17276 16244
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 17316 16192 17368 16244
rect 19156 16192 19208 16244
rect 4804 16056 4856 16108
rect 4988 16056 5040 16108
rect 5540 16056 5592 16108
rect 9772 16056 9824 16108
rect 10876 16099 10928 16108
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 1584 15988 1636 16040
rect 2596 16031 2648 16040
rect 2596 15997 2605 16031
rect 2605 15997 2639 16031
rect 2639 15997 2648 16031
rect 2596 15988 2648 15997
rect 4160 15988 4212 16040
rect 4620 15988 4672 16040
rect 1952 15920 2004 15972
rect 3884 15852 3936 15904
rect 4344 15920 4396 15972
rect 5540 15920 5592 15972
rect 6092 15920 6144 15972
rect 4988 15895 5040 15904
rect 4988 15861 4997 15895
rect 4997 15861 5031 15895
rect 5031 15861 5040 15895
rect 4988 15852 5040 15861
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 8576 15988 8628 16040
rect 9128 15988 9180 16040
rect 10324 15988 10376 16040
rect 10876 16065 10885 16099
rect 10885 16065 10919 16099
rect 10919 16065 10928 16099
rect 10876 16056 10928 16065
rect 13452 16056 13504 16108
rect 7656 15920 7708 15972
rect 10232 15920 10284 15972
rect 10692 15988 10744 16040
rect 7196 15852 7248 15861
rect 9588 15852 9640 15904
rect 10876 15852 10928 15904
rect 11428 15852 11480 15904
rect 11704 15852 11756 15904
rect 11888 15920 11940 15972
rect 12164 15852 12216 15904
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 15384 15988 15436 16040
rect 18328 16031 18380 16040
rect 18328 15997 18337 16031
rect 18337 15997 18371 16031
rect 18371 15997 18380 16031
rect 18328 15988 18380 15997
rect 21180 16031 21232 16040
rect 21180 15997 21214 16031
rect 21214 15997 21232 16031
rect 14924 15963 14976 15972
rect 14924 15929 14958 15963
rect 14958 15929 14976 15963
rect 14924 15920 14976 15929
rect 18788 15920 18840 15972
rect 19248 15920 19300 15972
rect 20444 15963 20496 15972
rect 15200 15852 15252 15904
rect 15660 15852 15712 15904
rect 16396 15852 16448 15904
rect 18420 15852 18472 15904
rect 19340 15852 19392 15904
rect 20444 15929 20453 15963
rect 20453 15929 20487 15963
rect 20487 15929 20496 15963
rect 20444 15920 20496 15929
rect 21180 15988 21232 15997
rect 22100 16192 22152 16244
rect 22560 16192 22612 16244
rect 23480 16235 23532 16244
rect 23480 16201 23489 16235
rect 23489 16201 23523 16235
rect 23523 16201 23532 16235
rect 23480 16192 23532 16201
rect 24952 16235 25004 16244
rect 24952 16201 24961 16235
rect 24961 16201 24995 16235
rect 24995 16201 25004 16235
rect 24952 16192 25004 16201
rect 25504 16192 25556 16244
rect 23388 16124 23440 16176
rect 24400 16124 24452 16176
rect 25228 16124 25280 16176
rect 24216 16056 24268 16108
rect 24952 15988 25004 16040
rect 26148 15988 26200 16040
rect 21456 15920 21508 15972
rect 23572 15920 23624 15972
rect 22100 15852 22152 15904
rect 23020 15852 23072 15904
rect 23480 15852 23532 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 3884 15691 3936 15700
rect 3884 15657 3893 15691
rect 3893 15657 3927 15691
rect 3927 15657 3936 15691
rect 3884 15648 3936 15657
rect 4252 15691 4304 15700
rect 4252 15657 4261 15691
rect 4261 15657 4295 15691
rect 4295 15657 4304 15691
rect 4252 15648 4304 15657
rect 4896 15648 4948 15700
rect 3148 15580 3200 15632
rect 4160 15580 4212 15632
rect 4344 15580 4396 15632
rect 5448 15648 5500 15700
rect 6460 15648 6512 15700
rect 6736 15691 6788 15700
rect 6736 15657 6745 15691
rect 6745 15657 6779 15691
rect 6779 15657 6788 15691
rect 6736 15648 6788 15657
rect 8760 15648 8812 15700
rect 9772 15648 9824 15700
rect 10692 15648 10744 15700
rect 10968 15691 11020 15700
rect 10968 15657 10977 15691
rect 10977 15657 11011 15691
rect 11011 15657 11020 15691
rect 10968 15648 11020 15657
rect 13452 15691 13504 15700
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 14740 15648 14792 15700
rect 17868 15691 17920 15700
rect 17868 15657 17877 15691
rect 17877 15657 17911 15691
rect 17911 15657 17920 15691
rect 17868 15648 17920 15657
rect 18420 15691 18472 15700
rect 18420 15657 18429 15691
rect 18429 15657 18463 15691
rect 18463 15657 18472 15691
rect 18420 15648 18472 15657
rect 20352 15648 20404 15700
rect 21180 15648 21232 15700
rect 6368 15580 6420 15632
rect 6644 15580 6696 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 3056 15555 3108 15564
rect 3056 15521 3065 15555
rect 3065 15521 3099 15555
rect 3099 15521 3108 15555
rect 3056 15512 3108 15521
rect 3976 15512 4028 15564
rect 6184 15512 6236 15564
rect 2688 15444 2740 15496
rect 5264 15444 5316 15496
rect 2504 15419 2556 15428
rect 2504 15385 2513 15419
rect 2513 15385 2547 15419
rect 2547 15385 2556 15419
rect 2504 15376 2556 15385
rect 4620 15376 4672 15428
rect 10692 15512 10744 15564
rect 11152 15512 11204 15564
rect 13820 15580 13872 15632
rect 14556 15580 14608 15632
rect 15200 15580 15252 15632
rect 15660 15623 15712 15632
rect 15660 15589 15669 15623
rect 15669 15589 15703 15623
rect 15703 15589 15712 15623
rect 15660 15580 15712 15589
rect 15844 15623 15896 15632
rect 15844 15589 15853 15623
rect 15853 15589 15887 15623
rect 15887 15589 15896 15623
rect 15844 15580 15896 15589
rect 17592 15580 17644 15632
rect 19432 15623 19484 15632
rect 19432 15589 19441 15623
rect 19441 15589 19475 15623
rect 19475 15589 19484 15623
rect 19432 15580 19484 15589
rect 21272 15580 21324 15632
rect 23204 15648 23256 15700
rect 23940 15648 23992 15700
rect 24400 15648 24452 15700
rect 23756 15580 23808 15632
rect 14924 15512 14976 15564
rect 15384 15512 15436 15564
rect 16396 15512 16448 15564
rect 6736 15444 6788 15496
rect 7840 15444 7892 15496
rect 8484 15444 8536 15496
rect 6092 15351 6144 15360
rect 6092 15317 6101 15351
rect 6101 15317 6135 15351
rect 6135 15317 6144 15351
rect 6092 15308 6144 15317
rect 7380 15308 7432 15360
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 7840 15351 7892 15360
rect 7840 15317 7849 15351
rect 7849 15317 7883 15351
rect 7883 15317 7892 15351
rect 7840 15308 7892 15317
rect 13636 15419 13688 15428
rect 13636 15385 13645 15419
rect 13645 15385 13679 15419
rect 13679 15385 13688 15419
rect 13636 15376 13688 15385
rect 14648 15444 14700 15496
rect 16672 15444 16724 15496
rect 18052 15444 18104 15496
rect 18512 15444 18564 15496
rect 20444 15512 20496 15564
rect 24584 15512 24636 15564
rect 20996 15444 21048 15496
rect 21456 15444 21508 15496
rect 24676 15487 24728 15496
rect 24676 15453 24685 15487
rect 24685 15453 24719 15487
rect 24719 15453 24728 15487
rect 24676 15444 24728 15453
rect 25136 15444 25188 15496
rect 16488 15376 16540 15428
rect 19248 15376 19300 15428
rect 24216 15419 24268 15428
rect 11428 15308 11480 15360
rect 12440 15351 12492 15360
rect 12440 15317 12449 15351
rect 12449 15317 12483 15351
rect 12483 15317 12492 15351
rect 12440 15308 12492 15317
rect 16672 15308 16724 15360
rect 16856 15308 16908 15360
rect 17868 15308 17920 15360
rect 18972 15351 19024 15360
rect 18972 15317 18981 15351
rect 18981 15317 19015 15351
rect 19015 15317 19024 15351
rect 18972 15308 19024 15317
rect 21272 15308 21324 15360
rect 24216 15385 24225 15419
rect 24225 15385 24259 15419
rect 24259 15385 24268 15419
rect 24216 15376 24268 15385
rect 22008 15308 22060 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1768 15147 1820 15156
rect 1768 15113 1777 15147
rect 1777 15113 1811 15147
rect 1811 15113 1820 15147
rect 1768 15104 1820 15113
rect 2688 15104 2740 15156
rect 3056 15104 3108 15156
rect 4344 15147 4396 15156
rect 4344 15113 4353 15147
rect 4353 15113 4387 15147
rect 4387 15113 4396 15147
rect 4344 15104 4396 15113
rect 5448 15104 5500 15156
rect 6368 15104 6420 15156
rect 6460 15104 6512 15156
rect 6920 15104 6972 15156
rect 4712 15079 4764 15088
rect 1952 14968 2004 15020
rect 2872 14968 2924 15020
rect 2320 14943 2372 14952
rect 2320 14909 2329 14943
rect 2329 14909 2363 14943
rect 2363 14909 2372 14943
rect 2320 14900 2372 14909
rect 4712 15045 4721 15079
rect 4721 15045 4755 15079
rect 4755 15045 4764 15079
rect 4712 15036 4764 15045
rect 5264 15036 5316 15088
rect 3792 14968 3844 15020
rect 5356 14968 5408 15020
rect 5080 14900 5132 14952
rect 6460 14900 6512 14952
rect 7932 15104 7984 15156
rect 10140 15104 10192 15156
rect 10784 15104 10836 15156
rect 12532 15079 12584 15088
rect 12532 15045 12541 15079
rect 12541 15045 12575 15079
rect 12575 15045 12584 15079
rect 12532 15036 12584 15045
rect 13820 15104 13872 15156
rect 14096 15147 14148 15156
rect 14096 15113 14105 15147
rect 14105 15113 14139 15147
rect 14139 15113 14148 15147
rect 14096 15104 14148 15113
rect 16948 15104 17000 15156
rect 17592 15104 17644 15156
rect 17776 15147 17828 15156
rect 17776 15113 17785 15147
rect 17785 15113 17819 15147
rect 17819 15113 17828 15147
rect 17776 15104 17828 15113
rect 19064 15104 19116 15156
rect 20720 15104 20772 15156
rect 20996 15147 21048 15156
rect 20996 15113 21005 15147
rect 21005 15113 21039 15147
rect 21039 15113 21048 15147
rect 20996 15104 21048 15113
rect 21088 15104 21140 15156
rect 23020 15147 23072 15156
rect 23020 15113 23029 15147
rect 23029 15113 23063 15147
rect 23063 15113 23072 15147
rect 23020 15104 23072 15113
rect 23204 15104 23256 15156
rect 18512 15079 18564 15088
rect 18512 15045 18521 15079
rect 18521 15045 18555 15079
rect 18555 15045 18564 15079
rect 18512 15036 18564 15045
rect 23572 15104 23624 15156
rect 25136 15104 25188 15156
rect 2228 14832 2280 14884
rect 3792 14875 3844 14884
rect 3792 14841 3801 14875
rect 3801 14841 3835 14875
rect 3835 14841 3844 14875
rect 3792 14832 3844 14841
rect 3884 14832 3936 14884
rect 3148 14764 3200 14816
rect 5172 14764 5224 14816
rect 6736 14832 6788 14884
rect 11060 15011 11112 15020
rect 11060 14977 11069 15011
rect 11069 14977 11103 15011
rect 11103 14977 11112 15011
rect 11060 14968 11112 14977
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 13452 14968 13504 15020
rect 15660 14968 15712 15020
rect 16672 14968 16724 15020
rect 17040 14968 17092 15020
rect 17960 14968 18012 15020
rect 20444 14968 20496 15020
rect 21640 14968 21692 15020
rect 23388 14968 23440 15020
rect 9588 14900 9640 14952
rect 9864 14900 9916 14952
rect 8484 14832 8536 14884
rect 10784 14875 10836 14884
rect 10784 14841 10793 14875
rect 10793 14841 10827 14875
rect 10827 14841 10836 14875
rect 10784 14832 10836 14841
rect 12072 14900 12124 14952
rect 12256 14875 12308 14884
rect 12256 14841 12265 14875
rect 12265 14841 12299 14875
rect 12299 14841 12308 14875
rect 12256 14832 12308 14841
rect 14372 14875 14424 14884
rect 14372 14841 14381 14875
rect 14381 14841 14415 14875
rect 14415 14841 14424 14875
rect 14372 14832 14424 14841
rect 14648 14875 14700 14884
rect 14648 14841 14657 14875
rect 14657 14841 14691 14875
rect 14691 14841 14700 14875
rect 14648 14832 14700 14841
rect 16672 14832 16724 14884
rect 16948 14875 17000 14884
rect 16948 14841 16957 14875
rect 16957 14841 16991 14875
rect 16991 14841 17000 14875
rect 16948 14832 17000 14841
rect 18788 14900 18840 14952
rect 21180 14900 21232 14952
rect 17224 14832 17276 14884
rect 19432 14832 19484 14884
rect 19892 14832 19944 14884
rect 22008 14832 22060 14884
rect 23296 14900 23348 14952
rect 25136 14900 25188 14952
rect 23020 14832 23072 14884
rect 24032 14875 24084 14884
rect 7196 14764 7248 14816
rect 7932 14764 7984 14816
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 11428 14764 11480 14816
rect 11888 14764 11940 14816
rect 14280 14764 14332 14816
rect 15384 14807 15436 14816
rect 15384 14773 15393 14807
rect 15393 14773 15427 14807
rect 15427 14773 15436 14807
rect 15384 14764 15436 14773
rect 20076 14764 20128 14816
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 22652 14764 22704 14816
rect 22744 14764 22796 14816
rect 23296 14764 23348 14816
rect 24032 14841 24041 14875
rect 24041 14841 24075 14875
rect 24075 14841 24084 14875
rect 24032 14832 24084 14841
rect 25504 14875 25556 14884
rect 25504 14841 25513 14875
rect 25513 14841 25547 14875
rect 25547 14841 25556 14875
rect 25504 14832 25556 14841
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2872 14603 2924 14612
rect 2872 14569 2881 14603
rect 2881 14569 2915 14603
rect 2915 14569 2924 14603
rect 2872 14560 2924 14569
rect 4712 14560 4764 14612
rect 5172 14560 5224 14612
rect 6644 14603 6696 14612
rect 6644 14569 6653 14603
rect 6653 14569 6687 14603
rect 6687 14569 6696 14603
rect 6644 14560 6696 14569
rect 6920 14603 6972 14612
rect 6920 14569 6929 14603
rect 6929 14569 6963 14603
rect 6963 14569 6972 14603
rect 6920 14560 6972 14569
rect 8852 14603 8904 14612
rect 8852 14569 8861 14603
rect 8861 14569 8895 14603
rect 8895 14569 8904 14603
rect 8852 14560 8904 14569
rect 9772 14560 9824 14612
rect 11152 14603 11204 14612
rect 11152 14569 11161 14603
rect 11161 14569 11195 14603
rect 11195 14569 11204 14603
rect 11152 14560 11204 14569
rect 11428 14560 11480 14612
rect 11704 14560 11756 14612
rect 1676 14492 1728 14544
rect 2596 14492 2648 14544
rect 4344 14492 4396 14544
rect 5448 14492 5500 14544
rect 8300 14492 8352 14544
rect 10048 14492 10100 14544
rect 12072 14560 12124 14612
rect 16764 14560 16816 14612
rect 17960 14560 18012 14612
rect 19248 14560 19300 14612
rect 19432 14603 19484 14612
rect 19432 14569 19441 14603
rect 19441 14569 19475 14603
rect 19475 14569 19484 14603
rect 19432 14560 19484 14569
rect 19984 14560 20036 14612
rect 20260 14603 20312 14612
rect 20260 14569 20269 14603
rect 20269 14569 20303 14603
rect 20303 14569 20312 14603
rect 20260 14560 20312 14569
rect 20720 14603 20772 14612
rect 20720 14569 20729 14603
rect 20729 14569 20763 14603
rect 20763 14569 20772 14603
rect 20720 14560 20772 14569
rect 15200 14492 15252 14544
rect 15660 14492 15712 14544
rect 17868 14492 17920 14544
rect 21364 14492 21416 14544
rect 21732 14560 21784 14612
rect 22008 14560 22060 14612
rect 23388 14560 23440 14612
rect 21640 14492 21692 14544
rect 3056 14424 3108 14476
rect 4712 14424 4764 14476
rect 6092 14424 6144 14476
rect 6644 14424 6696 14476
rect 7656 14424 7708 14476
rect 9312 14424 9364 14476
rect 3148 14356 3200 14408
rect 4160 14288 4212 14340
rect 3056 14220 3108 14272
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4252 14220 4304 14229
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 4988 14356 5040 14408
rect 6184 14356 6236 14408
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 8484 14399 8536 14408
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 11152 14424 11204 14476
rect 12440 14424 12492 14476
rect 14740 14424 14792 14476
rect 15384 14424 15436 14476
rect 19708 14467 19760 14476
rect 19708 14433 19717 14467
rect 19717 14433 19751 14467
rect 19751 14433 19760 14467
rect 19708 14424 19760 14433
rect 20168 14424 20220 14476
rect 20444 14424 20496 14476
rect 20720 14424 20772 14476
rect 23388 14424 23440 14476
rect 8484 14356 8536 14365
rect 4896 14288 4948 14340
rect 10508 14356 10560 14408
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 18420 14399 18472 14408
rect 18420 14365 18429 14399
rect 18429 14365 18463 14399
rect 18463 14365 18472 14399
rect 18420 14356 18472 14365
rect 21732 14356 21784 14408
rect 22652 14356 22704 14408
rect 14372 14288 14424 14340
rect 15200 14288 15252 14340
rect 18052 14288 18104 14340
rect 18972 14288 19024 14340
rect 20996 14331 21048 14340
rect 20996 14297 21005 14331
rect 21005 14297 21039 14331
rect 21039 14297 21048 14331
rect 20996 14288 21048 14297
rect 7196 14220 7248 14272
rect 7840 14220 7892 14272
rect 8484 14220 8536 14272
rect 9680 14220 9732 14272
rect 10968 14220 11020 14272
rect 11336 14220 11388 14272
rect 12072 14220 12124 14272
rect 13176 14220 13228 14272
rect 13452 14220 13504 14272
rect 14280 14220 14332 14272
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 16764 14220 16816 14272
rect 18788 14220 18840 14272
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 22744 14220 22796 14272
rect 25228 14263 25280 14272
rect 25228 14229 25237 14263
rect 25237 14229 25271 14263
rect 25271 14229 25280 14263
rect 25228 14220 25280 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 3056 14059 3108 14068
rect 3056 14025 3065 14059
rect 3065 14025 3099 14059
rect 3099 14025 3108 14059
rect 3056 14016 3108 14025
rect 3976 14016 4028 14068
rect 4896 14016 4948 14068
rect 5264 14016 5316 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 8208 14016 8260 14068
rect 8484 14016 8536 14068
rect 10048 14016 10100 14068
rect 10508 14059 10560 14068
rect 10508 14025 10517 14059
rect 10517 14025 10551 14059
rect 10551 14025 10560 14059
rect 10508 14016 10560 14025
rect 12900 14016 12952 14068
rect 13084 14016 13136 14068
rect 14556 14016 14608 14068
rect 16488 14059 16540 14068
rect 16488 14025 16497 14059
rect 16497 14025 16531 14059
rect 16531 14025 16540 14059
rect 16488 14016 16540 14025
rect 18512 14059 18564 14068
rect 18512 14025 18521 14059
rect 18521 14025 18555 14059
rect 18555 14025 18564 14059
rect 18512 14016 18564 14025
rect 18788 14016 18840 14068
rect 19708 14016 19760 14068
rect 21088 14016 21140 14068
rect 21456 14016 21508 14068
rect 22284 14016 22336 14068
rect 23020 14059 23072 14068
rect 23020 14025 23029 14059
rect 23029 14025 23063 14059
rect 23063 14025 23072 14059
rect 23020 14016 23072 14025
rect 24676 14016 24728 14068
rect 25228 14016 25280 14068
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 5908 13948 5960 14000
rect 8024 13948 8076 14000
rect 8392 13948 8444 14000
rect 16212 13948 16264 14000
rect 21364 13948 21416 14000
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 7656 13923 7708 13932
rect 6644 13812 6696 13864
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 16304 13923 16356 13932
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16948 13923 17000 13932
rect 16304 13880 16356 13889
rect 16948 13889 16957 13923
rect 16957 13889 16991 13923
rect 16991 13889 17000 13923
rect 16948 13880 17000 13889
rect 1952 13787 2004 13796
rect 1952 13753 1986 13787
rect 1986 13753 2004 13787
rect 1952 13744 2004 13753
rect 2044 13744 2096 13796
rect 2412 13744 2464 13796
rect 3976 13744 4028 13796
rect 4620 13744 4672 13796
rect 4988 13744 5040 13796
rect 7932 13812 7984 13864
rect 8852 13855 8904 13864
rect 8852 13821 8886 13855
rect 8886 13821 8904 13855
rect 8852 13812 8904 13821
rect 7564 13787 7616 13796
rect 7564 13753 7573 13787
rect 7573 13753 7607 13787
rect 7607 13753 7616 13787
rect 7564 13744 7616 13753
rect 7656 13744 7708 13796
rect 12256 13812 12308 13864
rect 17224 13880 17276 13932
rect 18420 13880 18472 13932
rect 11520 13744 11572 13796
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 6092 13719 6144 13728
rect 6092 13685 6101 13719
rect 6101 13685 6135 13719
rect 6135 13685 6144 13719
rect 6092 13676 6144 13685
rect 6828 13676 6880 13728
rect 7104 13676 7156 13728
rect 8116 13676 8168 13728
rect 9588 13676 9640 13728
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 11888 13676 11940 13728
rect 18512 13812 18564 13864
rect 21548 13923 21600 13932
rect 21548 13889 21557 13923
rect 21557 13889 21591 13923
rect 21591 13889 21600 13923
rect 21548 13880 21600 13889
rect 21640 13880 21692 13932
rect 13176 13744 13228 13796
rect 16488 13744 16540 13796
rect 17132 13744 17184 13796
rect 18972 13744 19024 13796
rect 15384 13719 15436 13728
rect 15384 13685 15393 13719
rect 15393 13685 15427 13719
rect 15427 13685 15436 13719
rect 15384 13676 15436 13685
rect 15844 13676 15896 13728
rect 16856 13676 16908 13728
rect 21088 13812 21140 13864
rect 21824 13812 21876 13864
rect 22652 13855 22704 13864
rect 22652 13821 22661 13855
rect 22661 13821 22695 13855
rect 22695 13821 22704 13855
rect 22652 13812 22704 13821
rect 23940 13812 23992 13864
rect 24676 13812 24728 13864
rect 25780 13855 25832 13864
rect 25780 13821 25789 13855
rect 25789 13821 25823 13855
rect 25823 13821 25832 13855
rect 25780 13812 25832 13821
rect 22192 13744 22244 13796
rect 22928 13744 22980 13796
rect 20168 13676 20220 13728
rect 22560 13676 22612 13728
rect 23480 13719 23532 13728
rect 23480 13685 23489 13719
rect 23489 13685 23523 13719
rect 23523 13685 23532 13719
rect 23480 13676 23532 13685
rect 24584 13676 24636 13728
rect 24768 13676 24820 13728
rect 25964 13676 26016 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1676 13472 1728 13524
rect 2596 13472 2648 13524
rect 2688 13472 2740 13524
rect 3332 13472 3384 13524
rect 5448 13472 5500 13524
rect 3056 13447 3108 13456
rect 3056 13413 3065 13447
rect 3065 13413 3099 13447
rect 3099 13413 3108 13447
rect 5908 13447 5960 13456
rect 3056 13404 3108 13413
rect 5908 13413 5917 13447
rect 5917 13413 5951 13447
rect 5951 13413 5960 13447
rect 5908 13404 5960 13413
rect 6368 13404 6420 13456
rect 1952 13336 2004 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 3148 13268 3200 13320
rect 3332 13336 3384 13388
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 5540 13336 5592 13388
rect 6460 13336 6512 13388
rect 7104 13336 7156 13388
rect 7472 13472 7524 13524
rect 8116 13472 8168 13524
rect 8852 13472 8904 13524
rect 9036 13472 9088 13524
rect 10048 13472 10100 13524
rect 11428 13472 11480 13524
rect 13176 13515 13228 13524
rect 13176 13481 13185 13515
rect 13185 13481 13219 13515
rect 13219 13481 13228 13515
rect 13176 13472 13228 13481
rect 14004 13472 14056 13524
rect 16488 13515 16540 13524
rect 8760 13404 8812 13456
rect 9588 13404 9640 13456
rect 10324 13404 10376 13456
rect 4344 13311 4396 13320
rect 4344 13277 4353 13311
rect 4353 13277 4387 13311
rect 4387 13277 4396 13311
rect 4344 13268 4396 13277
rect 5080 13268 5132 13320
rect 2320 13200 2372 13252
rect 5356 13200 5408 13252
rect 6184 13268 6236 13320
rect 7472 13268 7524 13320
rect 8024 13268 8076 13320
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 11060 13404 11112 13456
rect 11244 13404 11296 13456
rect 9680 13336 9732 13345
rect 10600 13336 10652 13388
rect 14096 13404 14148 13456
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 16764 13515 16816 13524
rect 16764 13481 16773 13515
rect 16773 13481 16807 13515
rect 16807 13481 16816 13515
rect 16764 13472 16816 13481
rect 19432 13515 19484 13524
rect 19432 13481 19441 13515
rect 19441 13481 19475 13515
rect 19475 13481 19484 13515
rect 19432 13472 19484 13481
rect 21456 13515 21508 13524
rect 21456 13481 21465 13515
rect 21465 13481 21499 13515
rect 21499 13481 21508 13515
rect 21456 13472 21508 13481
rect 22284 13515 22336 13524
rect 22284 13481 22293 13515
rect 22293 13481 22327 13515
rect 22327 13481 22336 13515
rect 22284 13472 22336 13481
rect 22652 13472 22704 13524
rect 23388 13472 23440 13524
rect 24584 13472 24636 13524
rect 24860 13472 24912 13524
rect 15936 13447 15988 13456
rect 15936 13413 15945 13447
rect 15945 13413 15979 13447
rect 15979 13413 15988 13447
rect 15936 13404 15988 13413
rect 17224 13447 17276 13456
rect 17224 13413 17258 13447
rect 17258 13413 17276 13447
rect 17224 13404 17276 13413
rect 18972 13447 19024 13456
rect 18972 13413 18981 13447
rect 18981 13413 19015 13447
rect 19015 13413 19024 13447
rect 18972 13404 19024 13413
rect 20076 13404 20128 13456
rect 21180 13404 21232 13456
rect 12348 13336 12400 13388
rect 14740 13336 14792 13388
rect 15660 13336 15712 13388
rect 16488 13336 16540 13388
rect 16856 13336 16908 13388
rect 17500 13336 17552 13388
rect 18512 13336 18564 13388
rect 19248 13336 19300 13388
rect 19432 13336 19484 13388
rect 22560 13336 22612 13388
rect 22928 13447 22980 13456
rect 22928 13413 22962 13447
rect 22962 13413 22980 13447
rect 22928 13404 22980 13413
rect 23940 13336 23992 13388
rect 25044 13336 25096 13388
rect 11612 13268 11664 13320
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 13084 13268 13136 13320
rect 13912 13268 13964 13320
rect 5908 13200 5960 13252
rect 6092 13200 6144 13252
rect 6828 13200 6880 13252
rect 3976 13132 4028 13184
rect 5080 13132 5132 13184
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 7564 13175 7616 13184
rect 7564 13141 7573 13175
rect 7573 13141 7607 13175
rect 7607 13141 7616 13175
rect 7564 13132 7616 13141
rect 7840 13175 7892 13184
rect 7840 13141 7849 13175
rect 7849 13141 7883 13175
rect 7883 13141 7892 13175
rect 7840 13132 7892 13141
rect 8208 13200 8260 13252
rect 11244 13243 11296 13252
rect 11244 13209 11253 13243
rect 11253 13209 11287 13243
rect 11287 13209 11296 13243
rect 11244 13200 11296 13209
rect 13728 13243 13780 13252
rect 13728 13209 13737 13243
rect 13737 13209 13771 13243
rect 13771 13209 13780 13243
rect 13728 13200 13780 13209
rect 14556 13268 14608 13320
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 21456 13268 21508 13320
rect 24952 13311 25004 13320
rect 24952 13277 24961 13311
rect 24961 13277 24995 13311
rect 24995 13277 25004 13311
rect 24952 13268 25004 13277
rect 14740 13200 14792 13252
rect 15752 13200 15804 13252
rect 20536 13200 20588 13252
rect 9312 13132 9364 13184
rect 10508 13175 10560 13184
rect 10508 13141 10517 13175
rect 10517 13141 10551 13175
rect 10551 13141 10560 13175
rect 10508 13132 10560 13141
rect 11428 13132 11480 13184
rect 13544 13175 13596 13184
rect 13544 13141 13553 13175
rect 13553 13141 13587 13175
rect 13587 13141 13596 13175
rect 13544 13132 13596 13141
rect 18328 13175 18380 13184
rect 18328 13141 18337 13175
rect 18337 13141 18371 13175
rect 18371 13141 18380 13175
rect 18328 13132 18380 13141
rect 19340 13175 19392 13184
rect 19340 13141 19349 13175
rect 19349 13141 19383 13175
rect 19383 13141 19392 13175
rect 19340 13132 19392 13141
rect 20168 13132 20220 13184
rect 21272 13132 21324 13184
rect 21732 13132 21784 13184
rect 24124 13132 24176 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2228 12928 2280 12980
rect 4160 12928 4212 12980
rect 6184 12928 6236 12980
rect 6460 12928 6512 12980
rect 6644 12928 6696 12980
rect 6920 12928 6972 12980
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 8576 12971 8628 12980
rect 8576 12937 8585 12971
rect 8585 12937 8619 12971
rect 8619 12937 8628 12971
rect 8576 12928 8628 12937
rect 9220 12928 9272 12980
rect 9588 12928 9640 12980
rect 11796 12928 11848 12980
rect 11888 12928 11940 12980
rect 3148 12860 3200 12912
rect 5080 12903 5132 12912
rect 5080 12869 5089 12903
rect 5089 12869 5123 12903
rect 5123 12869 5132 12903
rect 5080 12860 5132 12869
rect 2320 12792 2372 12844
rect 3056 12792 3108 12844
rect 3608 12792 3660 12844
rect 3884 12835 3936 12844
rect 3884 12801 3893 12835
rect 3893 12801 3927 12835
rect 3927 12801 3936 12835
rect 3884 12792 3936 12801
rect 7840 12860 7892 12912
rect 8760 12903 8812 12912
rect 8760 12869 8769 12903
rect 8769 12869 8803 12903
rect 8803 12869 8812 12903
rect 8760 12860 8812 12869
rect 9036 12860 9088 12912
rect 10876 12903 10928 12912
rect 6460 12792 6512 12844
rect 7196 12792 7248 12844
rect 7564 12792 7616 12844
rect 8576 12792 8628 12844
rect 9128 12792 9180 12844
rect 2780 12724 2832 12776
rect 2320 12699 2372 12708
rect 2320 12665 2329 12699
rect 2329 12665 2363 12699
rect 2363 12665 2372 12699
rect 2320 12656 2372 12665
rect 4068 12656 4120 12708
rect 4252 12656 4304 12708
rect 5264 12656 5316 12708
rect 6828 12724 6880 12776
rect 7288 12724 7340 12776
rect 8668 12724 8720 12776
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 9588 12724 9640 12776
rect 10324 12724 10376 12776
rect 6000 12699 6052 12708
rect 6000 12665 6009 12699
rect 6009 12665 6043 12699
rect 6043 12665 6052 12699
rect 6000 12656 6052 12665
rect 7104 12656 7156 12708
rect 7656 12699 7708 12708
rect 7656 12665 7665 12699
rect 7665 12665 7699 12699
rect 7699 12665 7708 12699
rect 7656 12656 7708 12665
rect 9128 12656 9180 12708
rect 9864 12656 9916 12708
rect 2412 12588 2464 12640
rect 3792 12631 3844 12640
rect 3792 12597 3801 12631
rect 3801 12597 3835 12631
rect 3835 12597 3844 12631
rect 3792 12588 3844 12597
rect 5080 12588 5132 12640
rect 7932 12588 7984 12640
rect 8852 12588 8904 12640
rect 10876 12869 10885 12903
rect 10885 12869 10919 12903
rect 10919 12869 10928 12903
rect 10876 12860 10928 12869
rect 11244 12835 11296 12844
rect 11244 12801 11253 12835
rect 11253 12801 11287 12835
rect 11287 12801 11296 12835
rect 11244 12792 11296 12801
rect 11612 12792 11664 12844
rect 12992 12928 13044 12980
rect 13544 12928 13596 12980
rect 15752 12928 15804 12980
rect 16028 12928 16080 12980
rect 16488 12971 16540 12980
rect 16488 12937 16497 12971
rect 16497 12937 16531 12971
rect 16531 12937 16540 12971
rect 16488 12928 16540 12937
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 19524 12928 19576 12980
rect 20720 12928 20772 12980
rect 23756 12971 23808 12980
rect 23756 12937 23765 12971
rect 23765 12937 23799 12971
rect 23799 12937 23808 12971
rect 23756 12928 23808 12937
rect 24676 12971 24728 12980
rect 13912 12903 13964 12912
rect 13912 12869 13921 12903
rect 13921 12869 13955 12903
rect 13955 12869 13964 12903
rect 13912 12860 13964 12869
rect 17224 12860 17276 12912
rect 18420 12860 18472 12912
rect 19156 12860 19208 12912
rect 21180 12860 21232 12912
rect 14556 12792 14608 12844
rect 15660 12792 15712 12844
rect 18328 12792 18380 12844
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 11428 12767 11480 12776
rect 11428 12733 11437 12767
rect 11437 12733 11471 12767
rect 11471 12733 11480 12767
rect 11428 12724 11480 12733
rect 10508 12656 10560 12708
rect 13544 12724 13596 12776
rect 14280 12724 14332 12776
rect 16764 12767 16816 12776
rect 16764 12733 16773 12767
rect 16773 12733 16807 12767
rect 16807 12733 16816 12767
rect 16764 12724 16816 12733
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 19248 12792 19300 12844
rect 20168 12792 20220 12844
rect 22284 12792 22336 12844
rect 24676 12937 24685 12971
rect 24685 12937 24719 12971
rect 24719 12937 24728 12971
rect 24676 12928 24728 12937
rect 25596 12928 25648 12980
rect 25044 12860 25096 12912
rect 17868 12724 17920 12733
rect 24216 12724 24268 12776
rect 24676 12724 24728 12776
rect 25504 12724 25556 12776
rect 13084 12699 13136 12708
rect 13084 12665 13093 12699
rect 13093 12665 13127 12699
rect 13127 12665 13136 12699
rect 13084 12656 13136 12665
rect 13912 12656 13964 12708
rect 18052 12656 18104 12708
rect 19800 12656 19852 12708
rect 21548 12656 21600 12708
rect 11244 12588 11296 12640
rect 13268 12588 13320 12640
rect 13544 12588 13596 12640
rect 16580 12588 16632 12640
rect 18972 12631 19024 12640
rect 18972 12597 18981 12631
rect 18981 12597 19015 12631
rect 19015 12597 19024 12631
rect 18972 12588 19024 12597
rect 19340 12588 19392 12640
rect 20536 12631 20588 12640
rect 20536 12597 20545 12631
rect 20545 12597 20579 12631
rect 20579 12597 20588 12631
rect 20536 12588 20588 12597
rect 21364 12631 21416 12640
rect 21364 12597 21373 12631
rect 21373 12597 21407 12631
rect 21407 12597 21416 12631
rect 21364 12588 21416 12597
rect 22652 12631 22704 12640
rect 22652 12597 22661 12631
rect 22661 12597 22695 12631
rect 22695 12597 22704 12631
rect 22652 12588 22704 12597
rect 23296 12588 23348 12640
rect 24216 12631 24268 12640
rect 24216 12597 24225 12631
rect 24225 12597 24259 12631
rect 24259 12597 24268 12631
rect 24216 12588 24268 12597
rect 25044 12631 25096 12640
rect 25044 12597 25053 12631
rect 25053 12597 25087 12631
rect 25087 12597 25096 12631
rect 25044 12588 25096 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1400 12427 1452 12436
rect 1400 12393 1409 12427
rect 1409 12393 1443 12427
rect 1443 12393 1452 12427
rect 1400 12384 1452 12393
rect 2320 12427 2372 12436
rect 2320 12393 2329 12427
rect 2329 12393 2363 12427
rect 2363 12393 2372 12427
rect 2320 12384 2372 12393
rect 3240 12384 3292 12436
rect 3608 12384 3660 12436
rect 4344 12384 4396 12436
rect 5264 12427 5316 12436
rect 5264 12393 5273 12427
rect 5273 12393 5307 12427
rect 5307 12393 5316 12427
rect 5264 12384 5316 12393
rect 6000 12384 6052 12436
rect 7656 12384 7708 12436
rect 8668 12427 8720 12436
rect 8668 12393 8677 12427
rect 8677 12393 8711 12427
rect 8711 12393 8720 12427
rect 8668 12384 8720 12393
rect 8852 12384 8904 12436
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 15752 12384 15804 12436
rect 16488 12384 16540 12436
rect 2504 12316 2556 12368
rect 2964 12359 3016 12368
rect 2964 12325 2973 12359
rect 2973 12325 3007 12359
rect 3007 12325 3016 12359
rect 2964 12316 3016 12325
rect 4620 12359 4672 12368
rect 4620 12325 4629 12359
rect 4629 12325 4663 12359
rect 4663 12325 4672 12359
rect 4620 12316 4672 12325
rect 4804 12359 4856 12368
rect 4804 12325 4813 12359
rect 4813 12325 4847 12359
rect 4847 12325 4856 12359
rect 4804 12316 4856 12325
rect 3332 12180 3384 12232
rect 5540 12316 5592 12368
rect 5448 12248 5500 12300
rect 6000 12248 6052 12300
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 6184 12248 6236 12257
rect 6460 12316 6512 12368
rect 8208 12359 8260 12368
rect 8208 12325 8217 12359
rect 8217 12325 8251 12359
rect 8251 12325 8260 12359
rect 8208 12316 8260 12325
rect 9680 12359 9732 12368
rect 9680 12325 9689 12359
rect 9689 12325 9723 12359
rect 9723 12325 9732 12359
rect 9680 12316 9732 12325
rect 13728 12359 13780 12368
rect 13728 12325 13737 12359
rect 13737 12325 13771 12359
rect 13771 12325 13780 12359
rect 13728 12316 13780 12325
rect 16396 12316 16448 12368
rect 18972 12384 19024 12436
rect 21088 12384 21140 12436
rect 22928 12384 22980 12436
rect 18420 12316 18472 12368
rect 20260 12359 20312 12368
rect 20260 12325 20269 12359
rect 20269 12325 20303 12359
rect 20303 12325 20312 12359
rect 20260 12316 20312 12325
rect 21456 12316 21508 12368
rect 6552 12248 6604 12300
rect 7380 12248 7432 12300
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 9036 12248 9088 12300
rect 9496 12248 9548 12300
rect 9956 12248 10008 12300
rect 10784 12248 10836 12300
rect 11428 12248 11480 12300
rect 13084 12291 13136 12300
rect 13084 12257 13093 12291
rect 13093 12257 13127 12291
rect 13127 12257 13136 12291
rect 13084 12248 13136 12257
rect 8300 12223 8352 12232
rect 2688 12112 2740 12164
rect 4436 12112 4488 12164
rect 4620 12112 4672 12164
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 10508 12180 10560 12232
rect 12072 12180 12124 12232
rect 12256 12180 12308 12232
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 14464 12248 14516 12300
rect 18052 12248 18104 12300
rect 18696 12248 18748 12300
rect 22652 12316 22704 12368
rect 25504 12316 25556 12368
rect 14004 12180 14056 12232
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 19156 12223 19208 12232
rect 19156 12189 19165 12223
rect 19165 12189 19199 12223
rect 19199 12189 19208 12223
rect 19156 12180 19208 12189
rect 20720 12180 20772 12232
rect 22560 12248 22612 12300
rect 23388 12248 23440 12300
rect 23848 12248 23900 12300
rect 24308 12223 24360 12232
rect 24308 12189 24317 12223
rect 24317 12189 24351 12223
rect 24351 12189 24360 12223
rect 24308 12180 24360 12189
rect 24952 12223 25004 12232
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 25228 12180 25280 12232
rect 8668 12112 8720 12164
rect 18972 12112 19024 12164
rect 21364 12112 21416 12164
rect 3792 12087 3844 12096
rect 3792 12053 3801 12087
rect 3801 12053 3835 12087
rect 3835 12053 3844 12087
rect 3792 12044 3844 12053
rect 5448 12044 5500 12096
rect 6552 12044 6604 12096
rect 7196 12044 7248 12096
rect 7656 12044 7708 12096
rect 7840 12044 7892 12096
rect 9496 12044 9548 12096
rect 10692 12044 10744 12096
rect 12072 12087 12124 12096
rect 12072 12053 12081 12087
rect 12081 12053 12115 12087
rect 12115 12053 12124 12087
rect 12072 12044 12124 12053
rect 13084 12044 13136 12096
rect 14280 12087 14332 12096
rect 14280 12053 14289 12087
rect 14289 12053 14323 12087
rect 14323 12053 14332 12087
rect 14280 12044 14332 12053
rect 17776 12087 17828 12096
rect 17776 12053 17785 12087
rect 17785 12053 17819 12087
rect 17819 12053 17828 12087
rect 17776 12044 17828 12053
rect 19248 12044 19300 12096
rect 20628 12044 20680 12096
rect 21548 12087 21600 12096
rect 21548 12053 21557 12087
rect 21557 12053 21591 12087
rect 21591 12053 21600 12087
rect 21548 12044 21600 12053
rect 23756 12044 23808 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2780 11883 2832 11892
rect 2780 11849 2789 11883
rect 2789 11849 2823 11883
rect 2823 11849 2832 11883
rect 2780 11840 2832 11849
rect 4436 11840 4488 11892
rect 6368 11883 6420 11892
rect 6368 11849 6377 11883
rect 6377 11849 6411 11883
rect 6411 11849 6420 11883
rect 6368 11840 6420 11849
rect 7196 11840 7248 11892
rect 8208 11840 8260 11892
rect 8484 11883 8536 11892
rect 8484 11849 8493 11883
rect 8493 11849 8527 11883
rect 8527 11849 8536 11883
rect 8484 11840 8536 11849
rect 9128 11840 9180 11892
rect 9588 11840 9640 11892
rect 10140 11840 10192 11892
rect 10508 11883 10560 11892
rect 10508 11849 10517 11883
rect 10517 11849 10551 11883
rect 10551 11849 10560 11883
rect 10508 11840 10560 11849
rect 11336 11840 11388 11892
rect 14004 11840 14056 11892
rect 19432 11883 19484 11892
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 21640 11840 21692 11892
rect 22652 11840 22704 11892
rect 25044 11883 25096 11892
rect 2596 11772 2648 11824
rect 2780 11704 2832 11756
rect 4068 11704 4120 11756
rect 5448 11772 5500 11824
rect 7012 11772 7064 11824
rect 7104 11772 7156 11824
rect 7840 11772 7892 11824
rect 1584 11636 1636 11688
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 5264 11704 5316 11756
rect 10692 11815 10744 11824
rect 10692 11781 10701 11815
rect 10701 11781 10735 11815
rect 10735 11781 10744 11815
rect 10692 11772 10744 11781
rect 15384 11772 15436 11824
rect 18788 11772 18840 11824
rect 19984 11815 20036 11824
rect 19984 11781 19993 11815
rect 19993 11781 20027 11815
rect 20027 11781 20036 11815
rect 19984 11772 20036 11781
rect 20076 11772 20128 11824
rect 23296 11772 23348 11824
rect 9588 11704 9640 11756
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 11612 11704 11664 11756
rect 12072 11704 12124 11756
rect 16304 11704 16356 11756
rect 19064 11704 19116 11756
rect 22284 11704 22336 11756
rect 22744 11704 22796 11756
rect 25044 11849 25053 11883
rect 25053 11849 25087 11883
rect 25087 11849 25096 11883
rect 25044 11840 25096 11849
rect 25964 11840 26016 11892
rect 4344 11636 4396 11688
rect 6460 11636 6512 11688
rect 8300 11636 8352 11688
rect 9220 11636 9272 11688
rect 10876 11636 10928 11688
rect 1676 11611 1728 11620
rect 1676 11577 1685 11611
rect 1685 11577 1719 11611
rect 1719 11577 1728 11611
rect 1676 11568 1728 11577
rect 3424 11568 3476 11620
rect 5448 11568 5500 11620
rect 8944 11611 8996 11620
rect 8944 11577 8953 11611
rect 8953 11577 8987 11611
rect 8987 11577 8996 11611
rect 8944 11568 8996 11577
rect 11060 11568 11112 11620
rect 11428 11568 11480 11620
rect 11980 11568 12032 11620
rect 6276 11500 6328 11552
rect 6828 11500 6880 11552
rect 6920 11500 6972 11552
rect 10876 11500 10928 11552
rect 11796 11500 11848 11552
rect 13176 11636 13228 11688
rect 15752 11636 15804 11688
rect 18696 11636 18748 11688
rect 19432 11636 19484 11688
rect 14280 11568 14332 11620
rect 14556 11568 14608 11620
rect 15568 11568 15620 11620
rect 12808 11500 12860 11552
rect 16672 11568 16724 11620
rect 18880 11611 18932 11620
rect 18880 11577 18889 11611
rect 18889 11577 18923 11611
rect 18923 11577 18932 11611
rect 18880 11568 18932 11577
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 19340 11500 19392 11552
rect 20352 11568 20404 11620
rect 20628 11568 20680 11620
rect 21272 11636 21324 11688
rect 25596 11679 25648 11688
rect 22008 11611 22060 11620
rect 20168 11500 20220 11552
rect 22008 11577 22017 11611
rect 22017 11577 22051 11611
rect 22051 11577 22060 11611
rect 22008 11568 22060 11577
rect 24768 11568 24820 11620
rect 25596 11645 25605 11679
rect 25605 11645 25639 11679
rect 25639 11645 25648 11679
rect 25596 11636 25648 11645
rect 26332 11568 26384 11620
rect 25504 11500 25556 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 3240 11296 3292 11348
rect 3332 11296 3384 11348
rect 4344 11296 4396 11348
rect 5908 11296 5960 11348
rect 6184 11296 6236 11348
rect 7564 11296 7616 11348
rect 11060 11296 11112 11348
rect 11888 11296 11940 11348
rect 2964 11271 3016 11280
rect 2964 11237 2973 11271
rect 2973 11237 3007 11271
rect 3007 11237 3016 11271
rect 2964 11228 3016 11237
rect 7104 11271 7156 11280
rect 3240 11160 3292 11212
rect 7104 11237 7113 11271
rect 7113 11237 7147 11271
rect 7147 11237 7156 11271
rect 7104 11228 7156 11237
rect 4804 11160 4856 11212
rect 8484 11228 8536 11280
rect 10140 11228 10192 11280
rect 10968 11228 11020 11280
rect 12624 11228 12676 11280
rect 8116 11203 8168 11212
rect 8116 11169 8125 11203
rect 8125 11169 8159 11203
rect 8159 11169 8168 11203
rect 8116 11160 8168 11169
rect 3056 11092 3108 11144
rect 3332 11092 3384 11144
rect 2412 11024 2464 11076
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 5172 10956 5224 11008
rect 6552 11092 6604 11144
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 6644 11067 6696 11076
rect 6644 11033 6653 11067
rect 6653 11033 6687 11067
rect 6687 11033 6696 11067
rect 6644 11024 6696 11033
rect 6460 10999 6512 11008
rect 6460 10965 6469 10999
rect 6469 10965 6503 10999
rect 6503 10965 6512 10999
rect 6460 10956 6512 10965
rect 6920 10956 6972 11008
rect 8300 10956 8352 11008
rect 8760 11160 8812 11212
rect 11336 11160 11388 11212
rect 13176 11296 13228 11348
rect 15844 11339 15896 11348
rect 15844 11305 15853 11339
rect 15853 11305 15887 11339
rect 15887 11305 15896 11339
rect 15844 11296 15896 11305
rect 19064 11296 19116 11348
rect 12992 11228 13044 11280
rect 13084 11160 13136 11212
rect 16488 11271 16540 11280
rect 16488 11237 16522 11271
rect 16522 11237 16540 11271
rect 16488 11228 16540 11237
rect 18696 11271 18748 11280
rect 18696 11237 18705 11271
rect 18705 11237 18739 11271
rect 18739 11237 18748 11271
rect 20720 11339 20772 11348
rect 18696 11228 18748 11237
rect 19708 11271 19760 11280
rect 19708 11237 19717 11271
rect 19717 11237 19751 11271
rect 19751 11237 19760 11271
rect 20720 11305 20729 11339
rect 20729 11305 20763 11339
rect 20763 11305 20772 11339
rect 20720 11296 20772 11305
rect 21640 11296 21692 11348
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 19708 11228 19760 11237
rect 20628 11228 20680 11280
rect 22008 11228 22060 11280
rect 22836 11271 22888 11280
rect 22836 11237 22845 11271
rect 22845 11237 22879 11271
rect 22879 11237 22888 11271
rect 22836 11228 22888 11237
rect 23020 11271 23072 11280
rect 23020 11237 23029 11271
rect 23029 11237 23063 11271
rect 23063 11237 23072 11271
rect 23020 11228 23072 11237
rect 23480 11296 23532 11348
rect 24584 11339 24636 11348
rect 24584 11305 24593 11339
rect 24593 11305 24627 11339
rect 24627 11305 24636 11339
rect 24584 11296 24636 11305
rect 19432 11160 19484 11212
rect 8484 11092 8536 11144
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 15476 11135 15528 11144
rect 12440 11092 12492 11101
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 18512 11092 18564 11144
rect 20352 11092 20404 11144
rect 21456 11135 21508 11144
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 23480 11160 23532 11212
rect 24216 11160 24268 11212
rect 24768 11228 24820 11280
rect 25320 11296 25372 11348
rect 25596 11296 25648 11348
rect 26516 11228 26568 11280
rect 23112 11135 23164 11144
rect 21456 11092 21508 11101
rect 8760 11024 8812 11076
rect 9312 10956 9364 11008
rect 14924 11024 14976 11076
rect 17224 11024 17276 11076
rect 19156 11024 19208 11076
rect 22560 11067 22612 11076
rect 22560 11033 22569 11067
rect 22569 11033 22603 11067
rect 22603 11033 22612 11067
rect 22560 11024 22612 11033
rect 23112 11101 23121 11135
rect 23121 11101 23155 11135
rect 23155 11101 23164 11135
rect 23112 11092 23164 11101
rect 25044 11135 25096 11144
rect 25044 11101 25053 11135
rect 25053 11101 25087 11135
rect 25087 11101 25096 11135
rect 25044 11092 25096 11101
rect 25228 11092 25280 11144
rect 24124 11067 24176 11076
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 12072 10956 12124 10965
rect 13268 10956 13320 11008
rect 14556 10956 14608 11008
rect 15568 10956 15620 11008
rect 22468 10956 22520 11008
rect 23664 10999 23716 11008
rect 23664 10965 23673 10999
rect 23673 10965 23707 10999
rect 23707 10965 23716 10999
rect 23664 10956 23716 10965
rect 24124 11033 24133 11067
rect 24133 11033 24167 11067
rect 24167 11033 24176 11067
rect 24124 11024 24176 11033
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2688 10752 2740 10804
rect 3240 10795 3292 10804
rect 3240 10761 3249 10795
rect 3249 10761 3283 10795
rect 3283 10761 3292 10795
rect 3240 10752 3292 10761
rect 5540 10752 5592 10804
rect 9220 10752 9272 10804
rect 9864 10752 9916 10804
rect 2320 10616 2372 10668
rect 7564 10616 7616 10668
rect 10968 10752 11020 10804
rect 11428 10752 11480 10804
rect 11612 10795 11664 10804
rect 11612 10761 11621 10795
rect 11621 10761 11655 10795
rect 11655 10761 11664 10795
rect 11612 10752 11664 10761
rect 12992 10752 13044 10804
rect 14648 10752 14700 10804
rect 15844 10795 15896 10804
rect 15844 10761 15853 10795
rect 15853 10761 15887 10795
rect 15887 10761 15896 10795
rect 15844 10752 15896 10761
rect 16396 10752 16448 10804
rect 16580 10752 16632 10804
rect 18512 10752 18564 10804
rect 19064 10752 19116 10804
rect 21456 10795 21508 10804
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 10324 10727 10376 10736
rect 10324 10693 10333 10727
rect 10333 10693 10367 10727
rect 10367 10693 10376 10727
rect 10324 10684 10376 10693
rect 11336 10727 11388 10736
rect 11336 10693 11345 10727
rect 11345 10693 11379 10727
rect 11379 10693 11388 10727
rect 11336 10684 11388 10693
rect 12348 10684 12400 10736
rect 13176 10684 13228 10736
rect 13820 10684 13872 10736
rect 19340 10684 19392 10736
rect 19616 10684 19668 10736
rect 20168 10727 20220 10736
rect 20168 10693 20177 10727
rect 20177 10693 20211 10727
rect 20211 10693 20220 10727
rect 20168 10684 20220 10693
rect 21640 10684 21692 10736
rect 1952 10480 2004 10532
rect 2228 10480 2280 10532
rect 5632 10548 5684 10600
rect 4620 10480 4672 10532
rect 7196 10480 7248 10532
rect 12992 10616 13044 10668
rect 12440 10548 12492 10600
rect 13452 10591 13504 10600
rect 13452 10557 13461 10591
rect 13461 10557 13495 10591
rect 13495 10557 13504 10591
rect 13452 10548 13504 10557
rect 15384 10616 15436 10668
rect 16856 10616 16908 10668
rect 17868 10616 17920 10668
rect 22008 10752 22060 10804
rect 23020 10752 23072 10804
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 23480 10752 23532 10761
rect 24124 10752 24176 10804
rect 24768 10684 24820 10736
rect 10968 10480 11020 10532
rect 12072 10480 12124 10532
rect 13176 10523 13228 10532
rect 13176 10489 13201 10523
rect 13201 10489 13228 10523
rect 14556 10548 14608 10600
rect 16672 10548 16724 10600
rect 19984 10548 20036 10600
rect 22744 10616 22796 10668
rect 22836 10616 22888 10668
rect 13176 10480 13228 10489
rect 14832 10480 14884 10532
rect 15568 10480 15620 10532
rect 4804 10412 4856 10464
rect 5908 10412 5960 10464
rect 7012 10455 7064 10464
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 7564 10455 7616 10464
rect 7564 10421 7573 10455
rect 7573 10421 7607 10455
rect 7607 10421 7616 10455
rect 7564 10412 7616 10421
rect 11336 10412 11388 10464
rect 14648 10412 14700 10464
rect 16396 10480 16448 10532
rect 18972 10480 19024 10532
rect 20076 10480 20128 10532
rect 20720 10523 20772 10532
rect 20720 10489 20729 10523
rect 20729 10489 20763 10523
rect 20763 10489 20772 10523
rect 20720 10480 20772 10489
rect 22008 10480 22060 10532
rect 22468 10480 22520 10532
rect 22836 10480 22888 10532
rect 23204 10616 23256 10668
rect 23940 10616 23992 10668
rect 23664 10548 23716 10600
rect 24216 10548 24268 10600
rect 23204 10480 23256 10532
rect 19248 10412 19300 10464
rect 22100 10412 22152 10464
rect 23940 10480 23992 10532
rect 24676 10616 24728 10668
rect 25780 10616 25832 10668
rect 25228 10591 25280 10600
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25228 10548 25280 10557
rect 26240 10480 26292 10532
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 2504 10208 2556 10260
rect 2964 10183 3016 10192
rect 2964 10149 2973 10183
rect 2973 10149 3007 10183
rect 3007 10149 3016 10183
rect 2964 10140 3016 10149
rect 4068 10208 4120 10260
rect 4344 10251 4396 10260
rect 4344 10217 4353 10251
rect 4353 10217 4387 10251
rect 4387 10217 4396 10251
rect 4344 10208 4396 10217
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 5632 10208 5684 10260
rect 5172 10140 5224 10192
rect 6920 10140 6972 10192
rect 7196 10208 7248 10260
rect 9312 10208 9364 10260
rect 4620 10072 4672 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2688 10004 2740 10056
rect 3424 9936 3476 9988
rect 3056 9868 3108 9920
rect 4160 9868 4212 9920
rect 4344 10004 4396 10056
rect 5172 10004 5224 10056
rect 7564 10072 7616 10124
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 5908 10004 5960 10056
rect 6092 10004 6144 10056
rect 10140 10140 10192 10192
rect 10968 10208 11020 10260
rect 13176 10208 13228 10260
rect 16396 10251 16448 10260
rect 16396 10217 16405 10251
rect 16405 10217 16439 10251
rect 16439 10217 16448 10251
rect 16396 10208 16448 10217
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 19524 10251 19576 10260
rect 19524 10217 19533 10251
rect 19533 10217 19567 10251
rect 19567 10217 19576 10251
rect 19524 10208 19576 10217
rect 8300 10072 8352 10124
rect 12348 10140 12400 10192
rect 13268 10140 13320 10192
rect 13820 10140 13872 10192
rect 15568 10140 15620 10192
rect 15752 10140 15804 10192
rect 17500 10183 17552 10192
rect 17500 10149 17509 10183
rect 17509 10149 17543 10183
rect 17543 10149 17552 10183
rect 17500 10140 17552 10149
rect 17960 10183 18012 10192
rect 17960 10149 17969 10183
rect 17969 10149 18003 10183
rect 18003 10149 18012 10183
rect 17960 10140 18012 10149
rect 19064 10183 19116 10192
rect 19064 10149 19073 10183
rect 19073 10149 19107 10183
rect 19107 10149 19116 10183
rect 19064 10140 19116 10149
rect 20076 10183 20128 10192
rect 20076 10149 20085 10183
rect 20085 10149 20119 10183
rect 20119 10149 20128 10183
rect 20076 10140 20128 10149
rect 22008 10208 22060 10260
rect 23112 10208 23164 10260
rect 23940 10208 23992 10260
rect 25412 10208 25464 10260
rect 20720 10140 20772 10192
rect 21364 10140 21416 10192
rect 22468 10140 22520 10192
rect 10508 10072 10560 10124
rect 10232 10047 10284 10056
rect 4896 9936 4948 9988
rect 9220 9936 9272 9988
rect 7196 9868 7248 9920
rect 7748 9868 7800 9920
rect 9404 9868 9456 9920
rect 9680 9936 9732 9988
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 10416 10004 10468 10056
rect 10692 10004 10744 10056
rect 11060 9936 11112 9988
rect 11152 9936 11204 9988
rect 10416 9868 10468 9920
rect 10600 9868 10652 9920
rect 11428 9868 11480 9920
rect 11888 9911 11940 9920
rect 11888 9877 11897 9911
rect 11897 9877 11931 9911
rect 11931 9877 11940 9911
rect 11888 9868 11940 9877
rect 12992 10072 13044 10124
rect 13084 10004 13136 10056
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 15384 10072 15436 10124
rect 16488 10072 16540 10124
rect 23940 10072 23992 10124
rect 14556 10004 14608 10056
rect 17408 10047 17460 10056
rect 13728 9979 13780 9988
rect 13728 9945 13737 9979
rect 13737 9945 13771 9979
rect 13771 9945 13780 9979
rect 13728 9936 13780 9945
rect 14096 9936 14148 9988
rect 15476 9979 15528 9988
rect 14832 9868 14884 9920
rect 15476 9945 15485 9979
rect 15485 9945 15519 9979
rect 15519 9945 15528 9979
rect 15476 9936 15528 9945
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 17592 10004 17644 10013
rect 18604 9979 18656 9988
rect 18604 9945 18613 9979
rect 18613 9945 18647 9979
rect 18647 9945 18656 9979
rect 18604 9936 18656 9945
rect 19156 10047 19208 10056
rect 19156 10013 19165 10047
rect 19165 10013 19199 10047
rect 19199 10013 19208 10047
rect 20904 10047 20956 10056
rect 19156 10004 19208 10013
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 20904 10004 20956 10013
rect 22744 10004 22796 10056
rect 19248 9936 19300 9988
rect 23020 9936 23072 9988
rect 15568 9868 15620 9920
rect 17040 9911 17092 9920
rect 17040 9877 17049 9911
rect 17049 9877 17083 9911
rect 17083 9877 17092 9911
rect 17040 9868 17092 9877
rect 22008 9868 22060 9920
rect 23204 9911 23256 9920
rect 23204 9877 23213 9911
rect 23213 9877 23247 9911
rect 23247 9877 23256 9911
rect 23204 9868 23256 9877
rect 24676 9936 24728 9988
rect 25412 9936 25464 9988
rect 25964 9936 26016 9988
rect 24952 9868 25004 9920
rect 25228 9868 25280 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2688 9664 2740 9716
rect 4620 9707 4672 9716
rect 4620 9673 4629 9707
rect 4629 9673 4663 9707
rect 4663 9673 4672 9707
rect 4620 9664 4672 9673
rect 6276 9664 6328 9716
rect 7564 9664 7616 9716
rect 10600 9664 10652 9716
rect 2136 9639 2188 9648
rect 2136 9605 2145 9639
rect 2145 9605 2179 9639
rect 2179 9605 2188 9639
rect 2136 9596 2188 9605
rect 3148 9596 3200 9648
rect 4712 9596 4764 9648
rect 4896 9596 4948 9648
rect 5264 9639 5316 9648
rect 5264 9605 5273 9639
rect 5273 9605 5307 9639
rect 5307 9605 5316 9639
rect 5264 9596 5316 9605
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 3792 9528 3844 9580
rect 4160 9528 4212 9580
rect 4344 9528 4396 9580
rect 6184 9528 6236 9580
rect 2504 9460 2556 9512
rect 3884 9460 3936 9512
rect 5172 9460 5224 9512
rect 5632 9460 5684 9512
rect 8944 9596 8996 9648
rect 10876 9639 10928 9648
rect 10876 9605 10885 9639
rect 10885 9605 10919 9639
rect 10919 9605 10928 9639
rect 10876 9596 10928 9605
rect 8576 9528 8628 9580
rect 7288 9460 7340 9512
rect 2228 9324 2280 9376
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 7012 9392 7064 9444
rect 6276 9367 6328 9376
rect 6276 9333 6285 9367
rect 6285 9333 6319 9367
rect 6319 9333 6328 9367
rect 6276 9324 6328 9333
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 7564 9392 7616 9444
rect 9312 9528 9364 9580
rect 9680 9528 9732 9580
rect 10048 9528 10100 9580
rect 10140 9503 10192 9512
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 10508 9460 10560 9512
rect 11888 9664 11940 9716
rect 11980 9596 12032 9648
rect 12348 9596 12400 9648
rect 11428 9571 11480 9580
rect 11428 9537 11437 9571
rect 11437 9537 11471 9571
rect 11471 9537 11480 9571
rect 11428 9528 11480 9537
rect 13452 9664 13504 9716
rect 16856 9707 16908 9716
rect 16856 9673 16865 9707
rect 16865 9673 16899 9707
rect 16899 9673 16908 9707
rect 16856 9664 16908 9673
rect 17592 9664 17644 9716
rect 19156 9664 19208 9716
rect 20536 9664 20588 9716
rect 20904 9707 20956 9716
rect 20904 9673 20913 9707
rect 20913 9673 20947 9707
rect 20947 9673 20956 9707
rect 20904 9664 20956 9673
rect 21272 9664 21324 9716
rect 21456 9664 21508 9716
rect 22284 9664 22336 9716
rect 23664 9664 23716 9716
rect 24216 9664 24268 9716
rect 14464 9596 14516 9648
rect 16764 9596 16816 9648
rect 17316 9596 17368 9648
rect 17776 9639 17828 9648
rect 17776 9605 17785 9639
rect 17785 9605 17819 9639
rect 17819 9605 17828 9639
rect 17776 9596 17828 9605
rect 20076 9596 20128 9648
rect 14280 9571 14332 9580
rect 12348 9460 12400 9512
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 13176 9460 13228 9512
rect 13820 9460 13872 9512
rect 20904 9528 20956 9580
rect 21180 9528 21232 9580
rect 22744 9596 22796 9648
rect 23940 9596 23992 9648
rect 10232 9392 10284 9444
rect 10692 9392 10744 9444
rect 15476 9503 15528 9512
rect 15476 9469 15485 9503
rect 15485 9469 15519 9503
rect 15519 9469 15528 9503
rect 15476 9460 15528 9469
rect 15568 9460 15620 9512
rect 6552 9324 6604 9333
rect 9404 9324 9456 9376
rect 9956 9324 10008 9376
rect 11612 9324 11664 9376
rect 13084 9324 13136 9376
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 13728 9324 13780 9376
rect 14556 9392 14608 9444
rect 15844 9392 15896 9444
rect 16120 9324 16172 9376
rect 18328 9324 18380 9376
rect 19524 9460 19576 9512
rect 20628 9460 20680 9512
rect 23296 9528 23348 9580
rect 23204 9460 23256 9512
rect 23572 9460 23624 9512
rect 20352 9392 20404 9444
rect 24308 9528 24360 9580
rect 24676 9528 24728 9580
rect 25964 9571 26016 9580
rect 25964 9537 25973 9571
rect 25973 9537 26007 9571
rect 26007 9537 26016 9571
rect 25964 9528 26016 9537
rect 25228 9503 25280 9512
rect 25228 9469 25237 9503
rect 25237 9469 25271 9503
rect 25271 9469 25280 9503
rect 25228 9460 25280 9469
rect 18972 9324 19024 9376
rect 21180 9324 21232 9376
rect 25504 9435 25556 9444
rect 23112 9324 23164 9376
rect 23572 9324 23624 9376
rect 25504 9401 25513 9435
rect 25513 9401 25547 9435
rect 25547 9401 25556 9435
rect 25504 9392 25556 9401
rect 26332 9367 26384 9376
rect 26332 9333 26341 9367
rect 26341 9333 26375 9367
rect 26375 9333 26384 9367
rect 26332 9324 26384 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2596 9120 2648 9172
rect 3884 9120 3936 9172
rect 4160 9120 4212 9172
rect 1584 9052 1636 9104
rect 2044 9052 2096 9104
rect 2044 8916 2096 8968
rect 2688 8916 2740 8968
rect 4436 9095 4488 9104
rect 4436 9061 4445 9095
rect 4445 9061 4479 9095
rect 4479 9061 4488 9095
rect 4436 9052 4488 9061
rect 4988 9120 5040 9172
rect 5540 9120 5592 9172
rect 6184 9120 6236 9172
rect 9312 9120 9364 9172
rect 6828 9052 6880 9104
rect 10876 9052 10928 9104
rect 11612 9120 11664 9172
rect 11796 9120 11848 9172
rect 13544 9120 13596 9172
rect 16580 9120 16632 9172
rect 17132 9120 17184 9172
rect 18420 9163 18472 9172
rect 18420 9129 18429 9163
rect 18429 9129 18463 9163
rect 18463 9129 18472 9163
rect 18420 9120 18472 9129
rect 18788 9120 18840 9172
rect 18972 9120 19024 9172
rect 19524 9163 19576 9172
rect 11336 9052 11388 9104
rect 5448 8984 5500 9036
rect 6460 8984 6512 9036
rect 7564 9027 7616 9036
rect 7564 8993 7573 9027
rect 7573 8993 7607 9027
rect 7607 8993 7616 9027
rect 7564 8984 7616 8993
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 12440 9052 12492 9104
rect 16304 9052 16356 9104
rect 16856 9052 16908 9104
rect 19524 9129 19533 9163
rect 19533 9129 19567 9163
rect 19567 9129 19576 9163
rect 19524 9120 19576 9129
rect 20352 9163 20404 9172
rect 20352 9129 20361 9163
rect 20361 9129 20395 9163
rect 20395 9129 20404 9163
rect 20352 9120 20404 9129
rect 21180 9120 21232 9172
rect 22008 9120 22060 9172
rect 22836 9120 22888 9172
rect 23480 9120 23532 9172
rect 25872 9120 25924 9172
rect 25964 9120 26016 9172
rect 26148 9120 26200 9172
rect 20720 9095 20772 9104
rect 20720 9061 20729 9095
rect 20729 9061 20763 9095
rect 20763 9061 20772 9095
rect 20720 9052 20772 9061
rect 21456 9095 21508 9104
rect 21456 9061 21465 9095
rect 21465 9061 21499 9095
rect 21499 9061 21508 9095
rect 21456 9052 21508 9061
rect 12072 8984 12124 9036
rect 15384 8984 15436 9036
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 18328 8984 18380 9036
rect 18788 8984 18840 9036
rect 21180 8984 21232 9036
rect 2136 8848 2188 8900
rect 2780 8848 2832 8900
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 8944 8916 8996 8968
rect 11060 8916 11112 8968
rect 17224 8916 17276 8968
rect 21640 9052 21692 9104
rect 22100 9052 22152 9104
rect 25688 9095 25740 9104
rect 22744 8984 22796 9036
rect 25688 9061 25697 9095
rect 25697 9061 25731 9095
rect 25731 9061 25740 9095
rect 25688 9052 25740 9061
rect 23296 8984 23348 9036
rect 25504 8984 25556 9036
rect 26148 8984 26200 9036
rect 24860 8916 24912 8968
rect 3148 8848 3200 8900
rect 4344 8848 4396 8900
rect 2228 8780 2280 8832
rect 3056 8780 3108 8832
rect 4712 8780 4764 8832
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 9312 8848 9364 8900
rect 9680 8848 9732 8900
rect 14556 8848 14608 8900
rect 20996 8891 21048 8900
rect 6368 8780 6420 8832
rect 7012 8823 7064 8832
rect 7012 8789 7021 8823
rect 7021 8789 7055 8823
rect 7055 8789 7064 8823
rect 7012 8780 7064 8789
rect 7932 8823 7984 8832
rect 7932 8789 7941 8823
rect 7941 8789 7975 8823
rect 7975 8789 7984 8823
rect 7932 8780 7984 8789
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 8760 8780 8812 8832
rect 11336 8780 11388 8832
rect 11796 8823 11848 8832
rect 11796 8789 11805 8823
rect 11805 8789 11839 8823
rect 11839 8789 11848 8823
rect 11796 8780 11848 8789
rect 12348 8780 12400 8832
rect 14280 8780 14332 8832
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 20996 8857 21005 8891
rect 21005 8857 21039 8891
rect 21039 8857 21048 8891
rect 20996 8848 21048 8857
rect 15936 8780 15988 8832
rect 17592 8780 17644 8832
rect 19248 8780 19300 8832
rect 21364 8780 21416 8832
rect 21824 8823 21876 8832
rect 21824 8789 21833 8823
rect 21833 8789 21867 8823
rect 21867 8789 21876 8823
rect 21824 8780 21876 8789
rect 22008 8823 22060 8832
rect 22008 8789 22017 8823
rect 22017 8789 22051 8823
rect 22051 8789 22060 8823
rect 22008 8780 22060 8789
rect 22560 8780 22612 8832
rect 23940 8780 23992 8832
rect 25596 8780 25648 8832
rect 25872 8780 25924 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 4252 8576 4304 8628
rect 4436 8576 4488 8628
rect 6736 8576 6788 8628
rect 6920 8619 6972 8628
rect 6920 8585 6929 8619
rect 6929 8585 6963 8619
rect 6963 8585 6972 8619
rect 6920 8576 6972 8585
rect 11060 8576 11112 8628
rect 3148 8508 3200 8560
rect 4068 8508 4120 8560
rect 4988 8551 5040 8560
rect 4988 8517 4997 8551
rect 4997 8517 5031 8551
rect 5031 8517 5040 8551
rect 4988 8508 5040 8517
rect 6368 8508 6420 8560
rect 8116 8508 8168 8560
rect 2596 8440 2648 8492
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 4620 8440 4672 8492
rect 8668 8440 8720 8492
rect 10048 8440 10100 8492
rect 4252 8415 4304 8424
rect 3056 8304 3108 8356
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4252 8372 4304 8381
rect 5448 8415 5500 8424
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 7380 8372 7432 8424
rect 10876 8372 10928 8424
rect 11980 8372 12032 8424
rect 3884 8304 3936 8356
rect 4344 8304 4396 8356
rect 4620 8304 4672 8356
rect 2596 8236 2648 8288
rect 3792 8236 3844 8288
rect 7564 8304 7616 8356
rect 8024 8304 8076 8356
rect 8484 8347 8536 8356
rect 8484 8313 8493 8347
rect 8493 8313 8527 8347
rect 8527 8313 8536 8347
rect 8484 8304 8536 8313
rect 9220 8304 9272 8356
rect 9404 8304 9456 8356
rect 9680 8304 9732 8356
rect 12440 8576 12492 8628
rect 14372 8619 14424 8628
rect 14372 8585 14381 8619
rect 14381 8585 14415 8619
rect 14415 8585 14424 8619
rect 14372 8576 14424 8585
rect 15568 8619 15620 8628
rect 15568 8585 15577 8619
rect 15577 8585 15611 8619
rect 15611 8585 15620 8619
rect 15568 8576 15620 8585
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 18972 8576 19024 8628
rect 19064 8576 19116 8628
rect 21272 8619 21324 8628
rect 21272 8585 21281 8619
rect 21281 8585 21315 8619
rect 21315 8585 21324 8619
rect 21272 8576 21324 8585
rect 21364 8576 21416 8628
rect 23112 8576 23164 8628
rect 24676 8619 24728 8628
rect 24676 8585 24685 8619
rect 24685 8585 24719 8619
rect 24719 8585 24728 8619
rect 24676 8576 24728 8585
rect 13820 8551 13872 8560
rect 13820 8517 13829 8551
rect 13829 8517 13863 8551
rect 13863 8517 13872 8551
rect 13820 8508 13872 8517
rect 14556 8508 14608 8560
rect 16672 8551 16724 8560
rect 16672 8517 16681 8551
rect 16681 8517 16715 8551
rect 16715 8517 16724 8551
rect 16672 8508 16724 8517
rect 17408 8551 17460 8560
rect 17408 8517 17417 8551
rect 17417 8517 17451 8551
rect 17451 8517 17460 8551
rect 17408 8508 17460 8517
rect 21456 8508 21508 8560
rect 23848 8508 23900 8560
rect 25044 8551 25096 8560
rect 25044 8517 25053 8551
rect 25053 8517 25087 8551
rect 25087 8517 25096 8551
rect 25044 8508 25096 8517
rect 25228 8508 25280 8560
rect 25596 8508 25648 8560
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 12992 8372 13044 8424
rect 18328 8372 18380 8424
rect 18972 8415 19024 8424
rect 18972 8381 19006 8415
rect 19006 8381 19024 8415
rect 18972 8372 19024 8381
rect 19248 8372 19300 8424
rect 23020 8372 23072 8424
rect 24676 8440 24728 8492
rect 10140 8236 10192 8288
rect 10876 8236 10928 8288
rect 12532 8304 12584 8356
rect 14188 8304 14240 8356
rect 16028 8347 16080 8356
rect 16028 8313 16037 8347
rect 16037 8313 16071 8347
rect 16071 8313 16080 8347
rect 16028 8304 16080 8313
rect 16212 8347 16264 8356
rect 16212 8313 16221 8347
rect 16221 8313 16255 8347
rect 16255 8313 16264 8347
rect 16212 8304 16264 8313
rect 16672 8304 16724 8356
rect 22008 8304 22060 8356
rect 23112 8347 23164 8356
rect 23112 8313 23121 8347
rect 23121 8313 23155 8347
rect 23155 8313 23164 8347
rect 25964 8576 26016 8628
rect 26148 8619 26200 8628
rect 26148 8585 26157 8619
rect 26157 8585 26191 8619
rect 26191 8585 26200 8619
rect 26148 8576 26200 8585
rect 23112 8304 23164 8313
rect 24400 8304 24452 8356
rect 13084 8236 13136 8288
rect 18328 8236 18380 8288
rect 21456 8236 21508 8288
rect 22284 8236 22336 8288
rect 22560 8236 22612 8288
rect 23388 8236 23440 8288
rect 23940 8236 23992 8288
rect 24124 8236 24176 8288
rect 25228 8236 25280 8288
rect 25412 8236 25464 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 3056 8032 3108 8084
rect 3424 8032 3476 8084
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 9220 8032 9272 8084
rect 9404 8032 9456 8084
rect 9864 8032 9916 8084
rect 10048 8032 10100 8084
rect 12072 8075 12124 8084
rect 12072 8041 12081 8075
rect 12081 8041 12115 8075
rect 12115 8041 12124 8075
rect 12072 8032 12124 8041
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 14464 8032 14516 8084
rect 14832 8032 14884 8084
rect 16304 8032 16356 8084
rect 18972 8075 19024 8084
rect 18972 8041 18981 8075
rect 18981 8041 19015 8075
rect 19015 8041 19024 8075
rect 18972 8032 19024 8041
rect 19340 8075 19392 8084
rect 19340 8041 19349 8075
rect 19349 8041 19383 8075
rect 19383 8041 19392 8075
rect 19340 8032 19392 8041
rect 19432 8032 19484 8084
rect 20812 8032 20864 8084
rect 21272 8032 21324 8084
rect 21824 8032 21876 8084
rect 24216 8075 24268 8084
rect 2964 8007 3016 8016
rect 2964 7973 2973 8007
rect 2973 7973 3007 8007
rect 3007 7973 3016 8007
rect 2964 7964 3016 7973
rect 4436 7964 4488 8016
rect 4896 7964 4948 8016
rect 7380 8007 7432 8016
rect 7380 7973 7414 8007
rect 7414 7973 7432 8007
rect 7380 7964 7432 7973
rect 10140 8007 10192 8016
rect 10140 7973 10174 8007
rect 10174 7973 10192 8007
rect 10140 7964 10192 7973
rect 2596 7896 2648 7948
rect 5264 7896 5316 7948
rect 6828 7896 6880 7948
rect 12992 7964 13044 8016
rect 16948 7964 17000 8016
rect 18604 7964 18656 8016
rect 21364 7964 21416 8016
rect 22008 7964 22060 8016
rect 22192 8007 22244 8016
rect 22192 7973 22226 8007
rect 22226 7973 22244 8007
rect 22192 7964 22244 7973
rect 24216 8041 24225 8075
rect 24225 8041 24259 8075
rect 24259 8041 24268 8075
rect 24216 8032 24268 8041
rect 24860 8032 24912 8084
rect 25688 8032 25740 8084
rect 26240 8075 26292 8084
rect 26240 8041 26249 8075
rect 26249 8041 26283 8075
rect 26283 8041 26292 8075
rect 26240 8032 26292 8041
rect 23756 7964 23808 8016
rect 24308 7964 24360 8016
rect 25412 8007 25464 8016
rect 25412 7973 25421 8007
rect 25421 7973 25455 8007
rect 25455 7973 25464 8007
rect 25412 7964 25464 7973
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 4620 7871 4672 7880
rect 2780 7760 2832 7812
rect 2412 7692 2464 7744
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 3976 7760 4028 7812
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 4344 7692 4396 7744
rect 6644 7828 6696 7880
rect 9864 7871 9916 7880
rect 6368 7760 6420 7812
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 12256 7828 12308 7880
rect 13728 7896 13780 7948
rect 17868 7896 17920 7948
rect 19432 7939 19484 7948
rect 19432 7905 19441 7939
rect 19441 7905 19475 7939
rect 19475 7905 19484 7939
rect 19432 7896 19484 7905
rect 21640 7896 21692 7948
rect 23572 7896 23624 7948
rect 24400 7896 24452 7948
rect 11244 7803 11296 7812
rect 11244 7769 11253 7803
rect 11253 7769 11287 7803
rect 11287 7769 11296 7803
rect 11244 7760 11296 7769
rect 12532 7760 12584 7812
rect 13820 7760 13872 7812
rect 14924 7760 14976 7812
rect 17592 7828 17644 7880
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 21824 7828 21876 7880
rect 24860 7871 24912 7880
rect 24860 7837 24869 7871
rect 24869 7837 24903 7871
rect 24903 7837 24912 7871
rect 24860 7828 24912 7837
rect 16856 7760 16908 7812
rect 21180 7760 21232 7812
rect 5540 7692 5592 7744
rect 6460 7692 6512 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 8300 7692 8352 7744
rect 8668 7692 8720 7744
rect 11152 7692 11204 7744
rect 11704 7692 11756 7744
rect 14096 7692 14148 7744
rect 16120 7735 16172 7744
rect 16120 7701 16129 7735
rect 16129 7701 16163 7735
rect 16163 7701 16172 7735
rect 16120 7692 16172 7701
rect 16580 7692 16632 7744
rect 17408 7735 17460 7744
rect 17408 7701 17417 7735
rect 17417 7701 17451 7735
rect 17451 7701 17460 7735
rect 17408 7692 17460 7701
rect 18512 7692 18564 7744
rect 21456 7735 21508 7744
rect 21456 7701 21465 7735
rect 21465 7701 21499 7735
rect 21499 7701 21508 7735
rect 21456 7692 21508 7701
rect 21640 7692 21692 7744
rect 23204 7760 23256 7812
rect 23296 7735 23348 7744
rect 23296 7701 23305 7735
rect 23305 7701 23339 7735
rect 23339 7701 23348 7735
rect 23296 7692 23348 7701
rect 24124 7760 24176 7812
rect 24676 7692 24728 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2964 7488 3016 7540
rect 4896 7531 4948 7540
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 6368 7488 6420 7540
rect 4344 7352 4396 7404
rect 8484 7488 8536 7540
rect 10140 7488 10192 7540
rect 10784 7488 10836 7540
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 11612 7488 11664 7540
rect 11888 7488 11940 7540
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 12900 7488 12952 7540
rect 13728 7488 13780 7540
rect 15936 7488 15988 7540
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 18236 7531 18288 7540
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 18696 7531 18748 7540
rect 18696 7497 18705 7531
rect 18705 7497 18739 7531
rect 18739 7497 18748 7531
rect 18696 7488 18748 7497
rect 21088 7531 21140 7540
rect 21088 7497 21097 7531
rect 21097 7497 21131 7531
rect 21131 7497 21140 7531
rect 21088 7488 21140 7497
rect 21732 7531 21784 7540
rect 21732 7497 21741 7531
rect 21741 7497 21775 7531
rect 21775 7497 21784 7531
rect 21732 7488 21784 7497
rect 22192 7488 22244 7540
rect 22560 7488 22612 7540
rect 22744 7531 22796 7540
rect 22744 7497 22753 7531
rect 22753 7497 22787 7531
rect 22787 7497 22796 7531
rect 23480 7531 23532 7540
rect 22744 7488 22796 7497
rect 9864 7420 9916 7472
rect 10876 7420 10928 7472
rect 12992 7463 13044 7472
rect 12992 7429 13001 7463
rect 13001 7429 13035 7463
rect 13035 7429 13044 7463
rect 12992 7420 13044 7429
rect 13544 7463 13596 7472
rect 13544 7429 13553 7463
rect 13553 7429 13587 7463
rect 13587 7429 13596 7463
rect 13544 7420 13596 7429
rect 18328 7420 18380 7472
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 22008 7420 22060 7472
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 24676 7531 24728 7540
rect 23480 7488 23532 7497
rect 12440 7352 12492 7361
rect 20352 7352 20404 7404
rect 23388 7420 23440 7472
rect 23572 7420 23624 7472
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 24952 7488 25004 7540
rect 25780 7488 25832 7540
rect 1860 7327 1912 7336
rect 1860 7293 1869 7327
rect 1869 7293 1903 7327
rect 1903 7293 1912 7327
rect 1860 7284 1912 7293
rect 3976 7284 4028 7336
rect 4620 7327 4672 7336
rect 4620 7293 4629 7327
rect 4629 7293 4663 7327
rect 4663 7293 4672 7327
rect 4620 7284 4672 7293
rect 5080 7284 5132 7336
rect 6920 7284 6972 7336
rect 8208 7284 8260 7336
rect 9772 7284 9824 7336
rect 10416 7284 10468 7336
rect 1676 7216 1728 7268
rect 2412 7216 2464 7268
rect 2688 7216 2740 7268
rect 4160 7216 4212 7268
rect 10048 7216 10100 7268
rect 14004 7284 14056 7336
rect 14372 7284 14424 7336
rect 18696 7284 18748 7336
rect 19248 7284 19300 7336
rect 21824 7284 21876 7336
rect 12256 7216 12308 7268
rect 3056 7148 3108 7200
rect 3424 7148 3476 7200
rect 4436 7148 4488 7200
rect 7380 7148 7432 7200
rect 9680 7148 9732 7200
rect 11704 7148 11756 7200
rect 13544 7148 13596 7200
rect 15200 7216 15252 7268
rect 17776 7216 17828 7268
rect 18328 7216 18380 7268
rect 19064 7216 19116 7268
rect 22192 7259 22244 7268
rect 22192 7225 22201 7259
rect 22201 7225 22235 7259
rect 22235 7225 22244 7259
rect 22192 7216 22244 7225
rect 15108 7148 15160 7200
rect 15384 7148 15436 7200
rect 16672 7148 16724 7200
rect 17592 7148 17644 7200
rect 17868 7191 17920 7200
rect 17868 7157 17877 7191
rect 17877 7157 17911 7191
rect 17911 7157 17920 7191
rect 17868 7148 17920 7157
rect 20260 7148 20312 7200
rect 24124 7216 24176 7268
rect 25504 7148 25556 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 3792 6944 3844 6996
rect 2596 6808 2648 6860
rect 4896 6876 4948 6928
rect 7380 6944 7432 6996
rect 8576 6944 8628 6996
rect 5448 6808 5500 6860
rect 6368 6808 6420 6860
rect 7472 6808 7524 6860
rect 8208 6808 8260 6860
rect 10048 6808 10100 6860
rect 2872 6783 2924 6792
rect 2872 6749 2881 6783
rect 2881 6749 2915 6783
rect 2915 6749 2924 6783
rect 2872 6740 2924 6749
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 5540 6740 5592 6792
rect 6460 6740 6512 6792
rect 2136 6672 2188 6724
rect 2504 6715 2556 6724
rect 2504 6681 2513 6715
rect 2513 6681 2547 6715
rect 2547 6681 2556 6715
rect 2504 6672 2556 6681
rect 1676 6604 1728 6656
rect 2596 6604 2648 6656
rect 4068 6604 4120 6656
rect 4344 6647 4396 6656
rect 4344 6613 4353 6647
rect 4353 6613 4387 6647
rect 4387 6613 4396 6647
rect 4344 6604 4396 6613
rect 4804 6647 4856 6656
rect 4804 6613 4813 6647
rect 4813 6613 4847 6647
rect 4847 6613 4856 6647
rect 4804 6604 4856 6613
rect 6644 6672 6696 6724
rect 6828 6740 6880 6792
rect 8484 6783 8536 6792
rect 7012 6672 7064 6724
rect 7380 6672 7432 6724
rect 7564 6672 7616 6724
rect 8208 6672 8260 6724
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 9496 6740 9548 6792
rect 9680 6740 9732 6792
rect 10876 6740 10928 6792
rect 11244 6876 11296 6928
rect 13544 6944 13596 6996
rect 12992 6876 13044 6928
rect 11244 6740 11296 6792
rect 12808 6851 12860 6860
rect 12808 6817 12842 6851
rect 12842 6817 12860 6851
rect 13820 6876 13872 6928
rect 14372 6944 14424 6996
rect 15200 6944 15252 6996
rect 14924 6876 14976 6928
rect 21640 6944 21692 6996
rect 22560 6944 22612 6996
rect 12808 6808 12860 6817
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 10692 6647 10744 6656
rect 10692 6613 10701 6647
rect 10701 6613 10735 6647
rect 10735 6613 10744 6647
rect 10692 6604 10744 6613
rect 11612 6647 11664 6656
rect 11612 6613 11621 6647
rect 11621 6613 11655 6647
rect 11655 6613 11664 6647
rect 11612 6604 11664 6613
rect 12348 6604 12400 6656
rect 12440 6647 12492 6656
rect 12440 6613 12449 6647
rect 12449 6613 12483 6647
rect 12483 6613 12492 6647
rect 14096 6672 14148 6724
rect 14280 6672 14332 6724
rect 14740 6672 14792 6724
rect 12440 6604 12492 6613
rect 13820 6604 13872 6656
rect 15384 6808 15436 6860
rect 15844 6808 15896 6860
rect 16212 6876 16264 6928
rect 16856 6876 16908 6928
rect 15200 6740 15252 6792
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 17592 6808 17644 6860
rect 19800 6876 19852 6928
rect 20352 6876 20404 6928
rect 22008 6876 22060 6928
rect 22652 6876 22704 6928
rect 23020 6919 23072 6928
rect 23020 6885 23029 6919
rect 23029 6885 23063 6919
rect 23063 6885 23072 6919
rect 23020 6876 23072 6885
rect 24584 6919 24636 6928
rect 17776 6808 17828 6860
rect 19064 6808 19116 6860
rect 19524 6808 19576 6860
rect 20444 6808 20496 6860
rect 20812 6808 20864 6860
rect 21732 6808 21784 6860
rect 23480 6851 23532 6860
rect 16488 6740 16540 6792
rect 19432 6740 19484 6792
rect 20536 6740 20588 6792
rect 20628 6740 20680 6792
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 23480 6817 23489 6851
rect 23489 6817 23523 6851
rect 23523 6817 23532 6851
rect 23480 6808 23532 6817
rect 24584 6885 24593 6919
rect 24593 6885 24627 6919
rect 24627 6885 24636 6919
rect 24584 6876 24636 6885
rect 25688 6876 25740 6928
rect 24216 6808 24268 6860
rect 25412 6851 25464 6860
rect 25412 6817 25421 6851
rect 25421 6817 25455 6851
rect 25455 6817 25464 6851
rect 25412 6808 25464 6817
rect 26424 6808 26476 6860
rect 20352 6672 20404 6724
rect 20996 6715 21048 6724
rect 20996 6681 21005 6715
rect 21005 6681 21039 6715
rect 21039 6681 21048 6715
rect 20996 6672 21048 6681
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 16948 6604 17000 6656
rect 17868 6604 17920 6656
rect 18696 6604 18748 6656
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 21916 6672 21968 6724
rect 21824 6604 21876 6656
rect 23204 6740 23256 6792
rect 24032 6672 24084 6724
rect 25044 6740 25096 6792
rect 25780 6783 25832 6792
rect 25780 6749 25789 6783
rect 25789 6749 25823 6783
rect 25823 6749 25832 6783
rect 25780 6740 25832 6749
rect 24860 6604 24912 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 5448 6400 5500 6452
rect 6092 6400 6144 6452
rect 6920 6443 6972 6452
rect 6920 6409 6929 6443
rect 6929 6409 6963 6443
rect 6963 6409 6972 6443
rect 6920 6400 6972 6409
rect 7932 6443 7984 6452
rect 7932 6409 7941 6443
rect 7941 6409 7975 6443
rect 7975 6409 7984 6443
rect 7932 6400 7984 6409
rect 8116 6400 8168 6452
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 4988 6332 5040 6384
rect 7012 6332 7064 6384
rect 7472 6264 7524 6316
rect 9404 6400 9456 6452
rect 10876 6400 10928 6452
rect 11244 6400 11296 6452
rect 12808 6400 12860 6452
rect 12992 6443 13044 6452
rect 12992 6409 13001 6443
rect 13001 6409 13035 6443
rect 13035 6409 13044 6443
rect 12992 6400 13044 6409
rect 14372 6400 14424 6452
rect 14740 6400 14792 6452
rect 15752 6400 15804 6452
rect 15844 6443 15896 6452
rect 15844 6409 15853 6443
rect 15853 6409 15887 6443
rect 15887 6409 15896 6443
rect 15844 6400 15896 6409
rect 16948 6400 17000 6452
rect 18512 6400 18564 6452
rect 19524 6443 19576 6452
rect 19524 6409 19533 6443
rect 19533 6409 19567 6443
rect 19567 6409 19576 6443
rect 19524 6400 19576 6409
rect 20444 6400 20496 6452
rect 21088 6400 21140 6452
rect 22560 6400 22612 6452
rect 25412 6443 25464 6452
rect 25412 6409 25421 6443
rect 25421 6409 25455 6443
rect 25455 6409 25464 6443
rect 25412 6400 25464 6409
rect 2504 6196 2556 6248
rect 3056 6196 3108 6248
rect 3240 6196 3292 6248
rect 3424 6196 3476 6248
rect 4620 6196 4672 6248
rect 10600 6264 10652 6316
rect 10876 6264 10928 6316
rect 11060 6264 11112 6316
rect 12256 6264 12308 6316
rect 5172 6128 5224 6180
rect 6828 6128 6880 6180
rect 7472 6171 7524 6180
rect 7472 6137 7481 6171
rect 7481 6137 7515 6171
rect 7515 6137 7524 6171
rect 7472 6128 7524 6137
rect 12992 6128 13044 6180
rect 13544 6128 13596 6180
rect 13820 6128 13872 6180
rect 17040 6332 17092 6384
rect 18144 6375 18196 6384
rect 18144 6341 18153 6375
rect 18153 6341 18187 6375
rect 18187 6341 18196 6375
rect 18144 6332 18196 6341
rect 19708 6375 19760 6384
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 19708 6341 19717 6375
rect 19717 6341 19751 6375
rect 19751 6341 19760 6375
rect 19708 6332 19760 6341
rect 21272 6375 21324 6384
rect 21272 6341 21281 6375
rect 21281 6341 21315 6375
rect 21315 6341 21324 6375
rect 21272 6332 21324 6341
rect 22008 6332 22060 6384
rect 23388 6332 23440 6384
rect 18696 6264 18748 6316
rect 16028 6196 16080 6248
rect 17592 6196 17644 6248
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 25964 6307 26016 6316
rect 25964 6273 25973 6307
rect 25973 6273 26007 6307
rect 26007 6273 26016 6307
rect 25964 6264 26016 6273
rect 18696 6171 18748 6180
rect 18696 6137 18705 6171
rect 18705 6137 18739 6171
rect 18739 6137 18748 6171
rect 18696 6128 18748 6137
rect 20812 6128 20864 6180
rect 22100 6196 22152 6248
rect 26608 6196 26660 6248
rect 21732 6171 21784 6180
rect 21732 6137 21741 6171
rect 21741 6137 21775 6171
rect 21775 6137 21784 6171
rect 21732 6128 21784 6137
rect 23020 6128 23072 6180
rect 24216 6128 24268 6180
rect 24492 6128 24544 6180
rect 25872 6128 25924 6180
rect 3240 6103 3292 6112
rect 3240 6069 3249 6103
rect 3249 6069 3283 6103
rect 3283 6069 3292 6103
rect 3240 6060 3292 6069
rect 5080 6060 5132 6112
rect 5540 6060 5592 6112
rect 5908 6060 5960 6112
rect 6368 6060 6420 6112
rect 7932 6060 7984 6112
rect 8300 6103 8352 6112
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 11520 6060 11572 6112
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 12808 6060 12860 6112
rect 15384 6103 15436 6112
rect 15384 6069 15393 6103
rect 15393 6069 15427 6103
rect 15427 6069 15436 6103
rect 15384 6060 15436 6069
rect 17776 6060 17828 6112
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 23204 6060 23256 6112
rect 25688 6060 25740 6112
rect 26332 6103 26384 6112
rect 26332 6069 26341 6103
rect 26341 6069 26375 6103
rect 26375 6069 26384 6103
rect 26332 6060 26384 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 2504 5899 2556 5908
rect 1768 5831 1820 5840
rect 1768 5797 1777 5831
rect 1777 5797 1811 5831
rect 1811 5797 1820 5831
rect 1768 5788 1820 5797
rect 2504 5865 2513 5899
rect 2513 5865 2547 5899
rect 2547 5865 2556 5899
rect 2504 5856 2556 5865
rect 3332 5856 3384 5908
rect 7104 5856 7156 5908
rect 8484 5856 8536 5908
rect 9496 5856 9548 5908
rect 12624 5856 12676 5908
rect 13820 5856 13872 5908
rect 14740 5899 14792 5908
rect 4620 5788 4672 5840
rect 2780 5720 2832 5772
rect 6920 5788 6972 5840
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 1952 5584 2004 5636
rect 2596 5584 2648 5636
rect 3240 5516 3292 5568
rect 4804 5516 4856 5568
rect 6276 5516 6328 5568
rect 6828 5720 6880 5772
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 8116 5788 8168 5840
rect 9772 5788 9824 5840
rect 10692 5788 10744 5840
rect 10784 5831 10836 5840
rect 10784 5797 10793 5831
rect 10793 5797 10827 5831
rect 10827 5797 10836 5831
rect 10784 5788 10836 5797
rect 11428 5788 11480 5840
rect 11796 5831 11848 5840
rect 11796 5797 11805 5831
rect 11805 5797 11839 5831
rect 11839 5797 11848 5831
rect 11796 5788 11848 5797
rect 7472 5720 7524 5772
rect 6920 5652 6972 5661
rect 9312 5652 9364 5704
rect 11244 5652 11296 5704
rect 13820 5720 13872 5772
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 16028 5856 16080 5908
rect 16304 5899 16356 5908
rect 16304 5865 16313 5899
rect 16313 5865 16347 5899
rect 16347 5865 16356 5899
rect 16304 5856 16356 5865
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 18696 5856 18748 5908
rect 20444 5856 20496 5908
rect 20812 5856 20864 5908
rect 21640 5856 21692 5908
rect 22652 5899 22704 5908
rect 22652 5865 22661 5899
rect 22661 5865 22695 5899
rect 22695 5865 22704 5899
rect 22652 5856 22704 5865
rect 14556 5788 14608 5840
rect 17040 5831 17092 5840
rect 17040 5797 17049 5831
rect 17049 5797 17083 5831
rect 17083 5797 17092 5831
rect 17040 5788 17092 5797
rect 17408 5788 17460 5840
rect 17868 5788 17920 5840
rect 18144 5788 18196 5840
rect 18972 5788 19024 5840
rect 22744 5788 22796 5840
rect 23388 5788 23440 5840
rect 25136 5856 25188 5908
rect 25872 5899 25924 5908
rect 25872 5865 25881 5899
rect 25881 5865 25915 5899
rect 25915 5865 25924 5899
rect 25872 5856 25924 5865
rect 14372 5720 14424 5772
rect 15660 5720 15712 5772
rect 16764 5720 16816 5772
rect 17960 5720 18012 5772
rect 9680 5584 9732 5636
rect 13176 5584 13228 5636
rect 8116 5516 8168 5568
rect 9312 5559 9364 5568
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 13084 5516 13136 5568
rect 13912 5652 13964 5704
rect 18604 5695 18656 5704
rect 16488 5584 16540 5636
rect 16028 5516 16080 5568
rect 17316 5516 17368 5568
rect 18604 5661 18613 5695
rect 18613 5661 18647 5695
rect 18647 5661 18656 5695
rect 18604 5652 18656 5661
rect 19340 5720 19392 5772
rect 19708 5763 19760 5772
rect 19708 5729 19717 5763
rect 19717 5729 19751 5763
rect 19751 5729 19760 5763
rect 19708 5720 19760 5729
rect 20076 5720 20128 5772
rect 21364 5720 21416 5772
rect 24216 5720 24268 5772
rect 24492 5720 24544 5772
rect 25228 5720 25280 5772
rect 25872 5720 25924 5772
rect 19248 5584 19300 5636
rect 20076 5584 20128 5636
rect 19524 5516 19576 5568
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 20628 5516 20680 5568
rect 24676 5652 24728 5704
rect 25136 5695 25188 5704
rect 25136 5661 25145 5695
rect 25145 5661 25179 5695
rect 25179 5661 25188 5695
rect 25136 5652 25188 5661
rect 25044 5584 25096 5636
rect 25964 5584 26016 5636
rect 22008 5516 22060 5568
rect 23940 5516 23992 5568
rect 25320 5516 25372 5568
rect 26240 5559 26292 5568
rect 26240 5525 26249 5559
rect 26249 5525 26283 5559
rect 26283 5525 26292 5559
rect 26240 5516 26292 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1492 5355 1544 5364
rect 1492 5321 1501 5355
rect 1501 5321 1535 5355
rect 1535 5321 1544 5355
rect 1492 5312 1544 5321
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 4620 5312 4672 5364
rect 8208 5312 8260 5364
rect 10048 5355 10100 5364
rect 10048 5321 10057 5355
rect 10057 5321 10091 5355
rect 10091 5321 10100 5355
rect 10048 5312 10100 5321
rect 11428 5312 11480 5364
rect 11612 5355 11664 5364
rect 11612 5321 11621 5355
rect 11621 5321 11655 5355
rect 11655 5321 11664 5355
rect 11612 5312 11664 5321
rect 13912 5312 13964 5364
rect 14372 5312 14424 5364
rect 5632 5244 5684 5296
rect 7288 5244 7340 5296
rect 12532 5287 12584 5296
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 2964 5219 3016 5228
rect 2964 5185 2973 5219
rect 2973 5185 3007 5219
rect 3007 5185 3016 5219
rect 2964 5176 3016 5185
rect 6736 5176 6788 5228
rect 9404 5176 9456 5228
rect 12532 5253 12541 5287
rect 12541 5253 12575 5287
rect 12575 5253 12584 5287
rect 12532 5244 12584 5253
rect 11612 5176 11664 5228
rect 12992 5219 13044 5228
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 13544 5176 13596 5228
rect 3240 5151 3292 5160
rect 2688 5040 2740 5092
rect 3240 5117 3274 5151
rect 3274 5117 3292 5151
rect 3240 5108 3292 5117
rect 5448 5151 5500 5160
rect 5448 5117 5457 5151
rect 5457 5117 5491 5151
rect 5491 5117 5500 5151
rect 5448 5108 5500 5117
rect 5540 5108 5592 5160
rect 5816 5108 5868 5160
rect 8116 5108 8168 5160
rect 10784 5108 10836 5160
rect 14464 5108 14516 5160
rect 17684 5312 17736 5364
rect 17868 5355 17920 5364
rect 17868 5321 17877 5355
rect 17877 5321 17911 5355
rect 17911 5321 17920 5355
rect 17868 5312 17920 5321
rect 18604 5312 18656 5364
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 18328 5244 18380 5296
rect 20628 5312 20680 5364
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 22008 5355 22060 5364
rect 22008 5321 22017 5355
rect 22017 5321 22051 5355
rect 22051 5321 22060 5355
rect 22008 5312 22060 5321
rect 23388 5312 23440 5364
rect 24860 5312 24912 5364
rect 25872 5312 25924 5364
rect 17776 5176 17828 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 18696 5219 18748 5228
rect 18696 5185 18705 5219
rect 18705 5185 18739 5219
rect 18739 5185 18748 5219
rect 18696 5176 18748 5185
rect 23020 5244 23072 5296
rect 26700 5244 26752 5296
rect 22284 5176 22336 5228
rect 25504 5219 25556 5228
rect 25504 5185 25513 5219
rect 25513 5185 25547 5219
rect 25547 5185 25556 5219
rect 25504 5176 25556 5185
rect 20260 5151 20312 5160
rect 20260 5117 20294 5151
rect 20294 5117 20312 5151
rect 20260 5108 20312 5117
rect 23480 5108 23532 5160
rect 2136 4972 2188 5024
rect 2964 4972 3016 5024
rect 3240 4972 3292 5024
rect 4804 4972 4856 5024
rect 6920 5040 6972 5092
rect 8760 5083 8812 5092
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 8760 5049 8769 5083
rect 8769 5049 8803 5083
rect 8803 5049 8812 5083
rect 8760 5040 8812 5049
rect 8944 5083 8996 5092
rect 8944 5049 8953 5083
rect 8953 5049 8987 5083
rect 8987 5049 8996 5083
rect 8944 5040 8996 5049
rect 13084 5083 13136 5092
rect 13084 5049 13093 5083
rect 13093 5049 13127 5083
rect 13127 5049 13136 5083
rect 13084 5040 13136 5049
rect 14740 5040 14792 5092
rect 6552 4972 6604 4981
rect 7656 4972 7708 5024
rect 10140 4972 10192 5024
rect 11060 4972 11112 5024
rect 12624 4972 12676 5024
rect 13912 4972 13964 5024
rect 16764 5040 16816 5092
rect 18604 5083 18656 5092
rect 18604 5049 18613 5083
rect 18613 5049 18647 5083
rect 18647 5049 18656 5083
rect 18604 5040 18656 5049
rect 22284 5083 22336 5092
rect 22284 5049 22293 5083
rect 22293 5049 22327 5083
rect 22327 5049 22336 5083
rect 22284 5040 22336 5049
rect 24676 5108 24728 5160
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 15384 4972 15436 5024
rect 17316 4972 17368 5024
rect 19984 4972 20036 5024
rect 22376 4972 22428 5024
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 23480 5015 23532 5024
rect 23480 4981 23489 5015
rect 23489 4981 23523 5015
rect 23523 4981 23532 5015
rect 25504 5040 25556 5092
rect 24216 5015 24268 5024
rect 23480 4972 23532 4981
rect 24216 4981 24225 5015
rect 24225 4981 24259 5015
rect 24259 4981 24268 5015
rect 24216 4972 24268 4981
rect 26332 5015 26384 5024
rect 26332 4981 26341 5015
rect 26341 4981 26375 5015
rect 26375 4981 26384 5015
rect 26332 4972 26384 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 2504 4768 2556 4820
rect 5080 4811 5132 4820
rect 5080 4777 5089 4811
rect 5089 4777 5123 4811
rect 5123 4777 5132 4811
rect 5080 4768 5132 4777
rect 5816 4768 5868 4820
rect 6000 4768 6052 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 6920 4811 6972 4820
rect 6920 4777 6929 4811
rect 6929 4777 6963 4811
rect 6963 4777 6972 4811
rect 6920 4768 6972 4777
rect 8300 4768 8352 4820
rect 8852 4768 8904 4820
rect 9404 4811 9456 4820
rect 9404 4777 9413 4811
rect 9413 4777 9447 4811
rect 9447 4777 9456 4811
rect 11244 4811 11296 4820
rect 9404 4768 9456 4777
rect 3516 4700 3568 4752
rect 6552 4700 6604 4752
rect 10048 4743 10100 4752
rect 4160 4632 4212 4684
rect 6000 4632 6052 4684
rect 8300 4632 8352 4684
rect 10048 4709 10057 4743
rect 10057 4709 10091 4743
rect 10091 4709 10100 4743
rect 10048 4700 10100 4709
rect 10232 4743 10284 4752
rect 10232 4709 10241 4743
rect 10241 4709 10275 4743
rect 10275 4709 10284 4743
rect 10232 4700 10284 4709
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 11612 4811 11664 4820
rect 11612 4777 11621 4811
rect 11621 4777 11655 4811
rect 11655 4777 11664 4811
rect 11612 4768 11664 4777
rect 12808 4768 12860 4820
rect 13636 4768 13688 4820
rect 14464 4768 14516 4820
rect 14740 4768 14792 4820
rect 15200 4768 15252 4820
rect 17408 4768 17460 4820
rect 20260 4768 20312 4820
rect 21364 4768 21416 4820
rect 24124 4768 24176 4820
rect 25136 4768 25188 4820
rect 25228 4768 25280 4820
rect 26240 4811 26292 4820
rect 26240 4777 26249 4811
rect 26249 4777 26283 4811
rect 26283 4777 26292 4811
rect 26240 4768 26292 4777
rect 10784 4743 10836 4752
rect 10784 4709 10793 4743
rect 10793 4709 10827 4743
rect 10827 4709 10836 4743
rect 10784 4700 10836 4709
rect 13820 4700 13872 4752
rect 10876 4632 10928 4684
rect 11244 4632 11296 4684
rect 12256 4632 12308 4684
rect 15384 4700 15436 4752
rect 15660 4743 15712 4752
rect 15660 4709 15669 4743
rect 15669 4709 15703 4743
rect 15703 4709 15712 4743
rect 15660 4700 15712 4709
rect 2504 4564 2556 4616
rect 3332 4564 3384 4616
rect 3976 4564 4028 4616
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 2320 4539 2372 4548
rect 2320 4505 2329 4539
rect 2329 4505 2363 4539
rect 2363 4505 2372 4539
rect 2320 4496 2372 4505
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 4344 4496 4396 4548
rect 6276 4564 6328 4616
rect 9680 4564 9732 4616
rect 10232 4564 10284 4616
rect 12624 4607 12676 4616
rect 12624 4573 12633 4607
rect 12633 4573 12667 4607
rect 12667 4573 12676 4607
rect 12624 4564 12676 4573
rect 14556 4632 14608 4684
rect 16672 4700 16724 4752
rect 18696 4700 18748 4752
rect 21180 4700 21232 4752
rect 22836 4743 22888 4752
rect 22836 4709 22845 4743
rect 22845 4709 22879 4743
rect 22879 4709 22888 4743
rect 22836 4700 22888 4709
rect 23020 4743 23072 4752
rect 23020 4709 23029 4743
rect 23029 4709 23063 4743
rect 23063 4709 23072 4743
rect 23020 4700 23072 4709
rect 16304 4632 16356 4684
rect 18144 4675 18196 4684
rect 18144 4641 18153 4675
rect 18153 4641 18187 4675
rect 18187 4641 18196 4675
rect 18328 4675 18380 4684
rect 18144 4632 18196 4641
rect 18328 4641 18337 4675
rect 18337 4641 18371 4675
rect 18371 4641 18380 4675
rect 18328 4632 18380 4641
rect 20904 4632 20956 4684
rect 21364 4632 21416 4684
rect 12992 4564 13044 4616
rect 5448 4496 5500 4548
rect 7656 4496 7708 4548
rect 8944 4496 8996 4548
rect 9772 4539 9824 4548
rect 9772 4505 9781 4539
rect 9781 4505 9815 4539
rect 9815 4505 9824 4539
rect 9772 4496 9824 4505
rect 12164 4539 12216 4548
rect 12164 4505 12173 4539
rect 12173 4505 12207 4539
rect 12207 4505 12216 4539
rect 12164 4496 12216 4505
rect 12440 4496 12492 4548
rect 13820 4496 13872 4548
rect 14464 4496 14516 4548
rect 1676 4428 1728 4437
rect 4068 4428 4120 4480
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 7288 4471 7340 4480
rect 4160 4428 4212 4437
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 14004 4428 14056 4480
rect 16488 4564 16540 4616
rect 17132 4607 17184 4616
rect 17132 4573 17141 4607
rect 17141 4573 17175 4607
rect 17175 4573 17184 4607
rect 17132 4564 17184 4573
rect 19432 4564 19484 4616
rect 22008 4632 22060 4684
rect 22192 4632 22244 4684
rect 24492 4700 24544 4752
rect 24124 4632 24176 4684
rect 15844 4496 15896 4548
rect 20996 4539 21048 4548
rect 20996 4505 21005 4539
rect 21005 4505 21039 4539
rect 21039 4505 21048 4539
rect 20996 4496 21048 4505
rect 21548 4607 21600 4616
rect 21548 4573 21557 4607
rect 21557 4573 21591 4607
rect 21591 4573 21600 4607
rect 21548 4564 21600 4573
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 22468 4496 22520 4548
rect 24216 4496 24268 4548
rect 17868 4428 17920 4480
rect 20628 4471 20680 4480
rect 20628 4437 20637 4471
rect 20637 4437 20671 4471
rect 20671 4437 20680 4471
rect 20628 4428 20680 4437
rect 22560 4471 22612 4480
rect 22560 4437 22569 4471
rect 22569 4437 22603 4471
rect 22603 4437 22612 4471
rect 25412 4471 25464 4480
rect 22560 4428 22612 4437
rect 25412 4437 25421 4471
rect 25421 4437 25455 4471
rect 25455 4437 25464 4471
rect 25412 4428 25464 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2136 4267 2188 4276
rect 2136 4233 2145 4267
rect 2145 4233 2179 4267
rect 2179 4233 2188 4267
rect 2136 4224 2188 4233
rect 3240 4267 3292 4276
rect 3240 4233 3249 4267
rect 3249 4233 3283 4267
rect 3283 4233 3292 4267
rect 3240 4224 3292 4233
rect 5448 4267 5500 4276
rect 5448 4233 5457 4267
rect 5457 4233 5491 4267
rect 5491 4233 5500 4267
rect 5448 4224 5500 4233
rect 6368 4267 6420 4276
rect 6368 4233 6377 4267
rect 6377 4233 6411 4267
rect 6411 4233 6420 4267
rect 6368 4224 6420 4233
rect 7012 4224 7064 4276
rect 8852 4224 8904 4276
rect 10140 4224 10192 4276
rect 12164 4267 12216 4276
rect 12164 4233 12173 4267
rect 12173 4233 12207 4267
rect 12207 4233 12216 4267
rect 12164 4224 12216 4233
rect 12624 4224 12676 4276
rect 12808 4224 12860 4276
rect 14188 4224 14240 4276
rect 14556 4224 14608 4276
rect 14740 4267 14792 4276
rect 14740 4233 14749 4267
rect 14749 4233 14783 4267
rect 14783 4233 14792 4267
rect 14740 4224 14792 4233
rect 17408 4267 17460 4276
rect 17408 4233 17417 4267
rect 17417 4233 17451 4267
rect 17451 4233 17460 4267
rect 17408 4224 17460 4233
rect 21640 4267 21692 4276
rect 21640 4233 21649 4267
rect 21649 4233 21683 4267
rect 21683 4233 21692 4267
rect 21640 4224 21692 4233
rect 22192 4224 22244 4276
rect 23020 4224 23072 4276
rect 23756 4267 23808 4276
rect 23756 4233 23765 4267
rect 23765 4233 23799 4267
rect 23799 4233 23808 4267
rect 23756 4224 23808 4233
rect 3516 4156 3568 4208
rect 8760 4199 8812 4208
rect 8760 4165 8769 4199
rect 8769 4165 8803 4199
rect 8803 4165 8812 4199
rect 8760 4156 8812 4165
rect 10232 4156 10284 4208
rect 10784 4156 10836 4208
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 3608 4088 3660 4140
rect 3884 4088 3936 4140
rect 7380 4088 7432 4140
rect 8300 4088 8352 4140
rect 9404 4088 9456 4140
rect 9864 4088 9916 4140
rect 10968 4131 11020 4140
rect 2228 4020 2280 4072
rect 2412 4063 2464 4072
rect 2412 4029 2421 4063
rect 2421 4029 2455 4063
rect 2455 4029 2464 4063
rect 2412 4020 2464 4029
rect 2320 3952 2372 4004
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 2044 3884 2096 3936
rect 2780 3884 2832 3936
rect 3976 3952 4028 4004
rect 4160 4020 4212 4072
rect 6000 4063 6052 4072
rect 6000 4029 6009 4063
rect 6009 4029 6043 4063
rect 6043 4029 6052 4063
rect 6000 4020 6052 4029
rect 6920 4020 6972 4072
rect 7288 4020 7340 4072
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 12256 4088 12308 4140
rect 14464 4156 14516 4208
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 14004 4131 14056 4140
rect 14004 4097 14013 4131
rect 14013 4097 14047 4131
rect 14047 4097 14056 4131
rect 22836 4156 22888 4208
rect 24124 4156 24176 4208
rect 14004 4088 14056 4097
rect 7748 3952 7800 4004
rect 8484 3952 8536 4004
rect 9496 3995 9548 4004
rect 9496 3961 9505 3995
rect 9505 3961 9539 3995
rect 9539 3961 9548 3995
rect 9496 3952 9548 3961
rect 10048 3952 10100 4004
rect 11888 3952 11940 4004
rect 14096 3952 14148 4004
rect 14740 4020 14792 4072
rect 16304 4020 16356 4072
rect 18144 3952 18196 4004
rect 22284 4131 22336 4140
rect 22284 4097 22293 4131
rect 22293 4097 22327 4131
rect 22327 4097 22336 4131
rect 22284 4088 22336 4097
rect 21548 4020 21600 4072
rect 22376 4020 22428 4072
rect 23388 4020 23440 4072
rect 23756 4020 23808 4072
rect 24584 4020 24636 4072
rect 25136 4063 25188 4072
rect 25136 4029 25145 4063
rect 25145 4029 25179 4063
rect 25179 4029 25188 4063
rect 25136 4020 25188 4029
rect 25412 4020 25464 4072
rect 20168 3952 20220 4004
rect 20904 3995 20956 4004
rect 20904 3961 20913 3995
rect 20913 3961 20947 3995
rect 20947 3961 20956 3995
rect 20904 3952 20956 3961
rect 22744 3952 22796 4004
rect 24216 3995 24268 4004
rect 24216 3961 24225 3995
rect 24225 3961 24259 3995
rect 24259 3961 24268 3995
rect 24216 3952 24268 3961
rect 24308 3995 24360 4004
rect 24308 3961 24317 3995
rect 24317 3961 24351 3995
rect 24351 3961 24360 3995
rect 24308 3952 24360 3961
rect 25504 3952 25556 4004
rect 3240 3884 3292 3936
rect 4068 3884 4120 3936
rect 6644 3884 6696 3936
rect 7932 3884 7984 3936
rect 11336 3884 11388 3936
rect 15292 3884 15344 3936
rect 15936 3884 15988 3936
rect 17868 3884 17920 3936
rect 18236 3884 18288 3936
rect 18696 3884 18748 3936
rect 19984 3927 20036 3936
rect 19984 3893 19993 3927
rect 19993 3893 20027 3927
rect 20027 3893 20036 3927
rect 19984 3884 20036 3893
rect 22008 3884 22060 3936
rect 22560 3884 22612 3936
rect 23388 3884 23440 3936
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 25136 3884 25188 3936
rect 26424 3884 26476 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 4160 3680 4212 3732
rect 5448 3680 5500 3732
rect 6276 3723 6328 3732
rect 6276 3689 6285 3723
rect 6285 3689 6319 3723
rect 6319 3689 6328 3723
rect 6276 3680 6328 3689
rect 10968 3680 11020 3732
rect 12992 3680 13044 3732
rect 15384 3680 15436 3732
rect 15844 3723 15896 3732
rect 15844 3689 15853 3723
rect 15853 3689 15887 3723
rect 15887 3689 15896 3723
rect 15844 3680 15896 3689
rect 17132 3723 17184 3732
rect 17132 3689 17141 3723
rect 17141 3689 17175 3723
rect 17175 3689 17184 3723
rect 17132 3680 17184 3689
rect 17408 3680 17460 3732
rect 18696 3723 18748 3732
rect 1676 3655 1728 3664
rect 1676 3621 1685 3655
rect 1685 3621 1719 3655
rect 1719 3621 1728 3655
rect 1676 3612 1728 3621
rect 2872 3612 2924 3664
rect 4528 3655 4580 3664
rect 4528 3621 4562 3655
rect 4562 3621 4580 3655
rect 4528 3612 4580 3621
rect 15660 3655 15712 3664
rect 3884 3544 3936 3596
rect 4068 3544 4120 3596
rect 2504 3451 2556 3460
rect 2504 3417 2513 3451
rect 2513 3417 2547 3451
rect 2547 3417 2556 3451
rect 2504 3408 2556 3417
rect 2044 3340 2096 3392
rect 3332 3476 3384 3528
rect 4896 3544 4948 3596
rect 7104 3544 7156 3596
rect 7288 3587 7340 3596
rect 7288 3553 7322 3587
rect 7322 3553 7340 3587
rect 7288 3544 7340 3553
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 11612 3544 11664 3596
rect 15660 3621 15669 3655
rect 15669 3621 15703 3655
rect 15703 3621 15712 3655
rect 15660 3612 15712 3621
rect 15936 3655 15988 3664
rect 15936 3621 15945 3655
rect 15945 3621 15979 3655
rect 15979 3621 15988 3655
rect 15936 3612 15988 3621
rect 17224 3612 17276 3664
rect 18236 3655 18288 3664
rect 18236 3621 18245 3655
rect 18245 3621 18279 3655
rect 18279 3621 18288 3655
rect 18236 3612 18288 3621
rect 18696 3689 18705 3723
rect 18705 3689 18739 3723
rect 18739 3689 18748 3723
rect 18696 3680 18748 3689
rect 19432 3680 19484 3732
rect 20812 3680 20864 3732
rect 21088 3680 21140 3732
rect 21640 3680 21692 3732
rect 22376 3723 22428 3732
rect 22376 3689 22385 3723
rect 22385 3689 22419 3723
rect 22419 3689 22428 3723
rect 22376 3680 22428 3689
rect 22652 3680 22704 3732
rect 24308 3680 24360 3732
rect 21548 3655 21600 3664
rect 21548 3621 21557 3655
rect 21557 3621 21591 3655
rect 21591 3621 21600 3655
rect 21548 3612 21600 3621
rect 23388 3612 23440 3664
rect 26240 3723 26292 3732
rect 26240 3689 26249 3723
rect 26249 3689 26283 3723
rect 26283 3689 26292 3723
rect 26240 3680 26292 3689
rect 26332 3612 26384 3664
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 14648 3544 14700 3553
rect 16856 3587 16908 3596
rect 16856 3553 16865 3587
rect 16865 3553 16899 3587
rect 16899 3553 16908 3587
rect 16856 3544 16908 3553
rect 20628 3544 20680 3596
rect 22468 3544 22520 3596
rect 24216 3544 24268 3596
rect 10968 3476 11020 3528
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 14372 3476 14424 3528
rect 19892 3519 19944 3528
rect 19892 3485 19901 3519
rect 19901 3485 19935 3519
rect 19935 3485 19944 3519
rect 19892 3476 19944 3485
rect 21548 3476 21600 3528
rect 23020 3519 23072 3528
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 25044 3519 25096 3528
rect 9496 3408 9548 3460
rect 13636 3451 13688 3460
rect 13636 3417 13645 3451
rect 13645 3417 13679 3451
rect 13679 3417 13688 3451
rect 13636 3408 13688 3417
rect 16580 3408 16632 3460
rect 17776 3451 17828 3460
rect 17776 3417 17785 3451
rect 17785 3417 17819 3451
rect 17819 3417 17828 3451
rect 17776 3408 17828 3417
rect 19340 3451 19392 3460
rect 19340 3417 19349 3451
rect 19349 3417 19383 3451
rect 19383 3417 19392 3451
rect 19340 3408 19392 3417
rect 21180 3408 21232 3460
rect 22376 3408 22428 3460
rect 22928 3408 22980 3460
rect 24032 3408 24084 3460
rect 24308 3408 24360 3460
rect 25044 3485 25053 3519
rect 25053 3485 25087 3519
rect 25087 3485 25096 3519
rect 25044 3476 25096 3485
rect 3516 3383 3568 3392
rect 3516 3349 3525 3383
rect 3525 3349 3559 3383
rect 3559 3349 3568 3383
rect 3516 3340 3568 3349
rect 6920 3383 6972 3392
rect 6920 3349 6929 3383
rect 6929 3349 6963 3383
rect 6963 3349 6972 3383
rect 6920 3340 6972 3349
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 12440 3383 12492 3392
rect 12440 3349 12449 3383
rect 12449 3349 12483 3383
rect 12483 3349 12492 3383
rect 12440 3340 12492 3349
rect 15292 3340 15344 3392
rect 16488 3383 16540 3392
rect 16488 3349 16497 3383
rect 16497 3349 16531 3383
rect 16531 3349 16540 3383
rect 16488 3340 16540 3349
rect 19064 3383 19116 3392
rect 19064 3349 19073 3383
rect 19073 3349 19107 3383
rect 19107 3349 19116 3383
rect 19064 3340 19116 3349
rect 22560 3383 22612 3392
rect 22560 3349 22569 3383
rect 22569 3349 22603 3383
rect 22603 3349 22612 3383
rect 22560 3340 22612 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1768 3136 1820 3188
rect 3332 3136 3384 3188
rect 3884 3136 3936 3188
rect 4068 3179 4120 3188
rect 4068 3145 4077 3179
rect 4077 3145 4111 3179
rect 4111 3145 4120 3179
rect 4068 3136 4120 3145
rect 4528 3136 4580 3188
rect 6368 3136 6420 3188
rect 7012 3136 7064 3188
rect 7104 3136 7156 3188
rect 3056 3068 3108 3120
rect 3424 3068 3476 3120
rect 1768 3000 1820 3052
rect 2504 3000 2556 3052
rect 3240 3043 3292 3052
rect 3240 3009 3249 3043
rect 3249 3009 3283 3043
rect 3283 3009 3292 3043
rect 3240 3000 3292 3009
rect 8484 3136 8536 3188
rect 9588 3136 9640 3188
rect 11428 3136 11480 3188
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 14740 3179 14792 3188
rect 14740 3145 14749 3179
rect 14749 3145 14783 3179
rect 14783 3145 14792 3179
rect 14740 3136 14792 3145
rect 15936 3136 15988 3188
rect 17224 3136 17276 3188
rect 17684 3179 17736 3188
rect 17684 3145 17693 3179
rect 17693 3145 17727 3179
rect 17727 3145 17736 3179
rect 17684 3136 17736 3145
rect 18144 3179 18196 3188
rect 18144 3145 18153 3179
rect 18153 3145 18187 3179
rect 18187 3145 18196 3179
rect 18144 3136 18196 3145
rect 22652 3136 22704 3188
rect 23020 3136 23072 3188
rect 23204 3179 23256 3188
rect 23204 3145 23213 3179
rect 23213 3145 23247 3179
rect 23247 3145 23256 3179
rect 23204 3136 23256 3145
rect 24216 3136 24268 3188
rect 26332 3179 26384 3188
rect 26332 3145 26341 3179
rect 26341 3145 26375 3179
rect 26375 3145 26384 3179
rect 26332 3136 26384 3145
rect 2964 2975 3016 2984
rect 2964 2941 2973 2975
rect 2973 2941 3007 2975
rect 3007 2941 3016 2975
rect 2964 2932 3016 2941
rect 7012 3000 7064 3052
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 14372 3000 14424 3052
rect 14556 3000 14608 3052
rect 16304 3111 16356 3120
rect 16304 3077 16313 3111
rect 16313 3077 16347 3111
rect 16347 3077 16356 3111
rect 16304 3068 16356 3077
rect 19340 3068 19392 3120
rect 20076 3068 20128 3120
rect 21548 3068 21600 3120
rect 23756 3111 23808 3120
rect 17960 3000 18012 3052
rect 18696 3000 18748 3052
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 21640 3043 21692 3052
rect 21640 3009 21649 3043
rect 21649 3009 21683 3043
rect 21683 3009 21692 3043
rect 21640 3000 21692 3009
rect 23756 3077 23765 3111
rect 23765 3077 23799 3111
rect 23799 3077 23808 3111
rect 23756 3068 23808 3077
rect 24860 3068 24912 3120
rect 24952 3000 25004 3052
rect 25412 3043 25464 3052
rect 25412 3009 25421 3043
rect 25421 3009 25455 3043
rect 25455 3009 25464 3043
rect 25412 3000 25464 3009
rect 5080 2932 5132 2984
rect 7288 2932 7340 2984
rect 8208 2932 8260 2984
rect 9312 2932 9364 2984
rect 9496 2975 9548 2984
rect 9496 2941 9519 2975
rect 9519 2941 9548 2975
rect 9496 2932 9548 2941
rect 2044 2907 2096 2916
rect 2044 2873 2053 2907
rect 2053 2873 2087 2907
rect 2087 2873 2096 2907
rect 2044 2864 2096 2873
rect 3516 2864 3568 2916
rect 5356 2864 5408 2916
rect 7748 2864 7800 2916
rect 9680 2864 9732 2916
rect 11428 2864 11480 2916
rect 13452 2932 13504 2984
rect 19064 2932 19116 2984
rect 19984 2932 20036 2984
rect 25228 2975 25280 2984
rect 25228 2941 25237 2975
rect 25237 2941 25271 2975
rect 25271 2941 25280 2975
rect 25228 2932 25280 2941
rect 15384 2864 15436 2916
rect 18604 2907 18656 2916
rect 18604 2873 18613 2907
rect 18613 2873 18647 2907
rect 18647 2873 18656 2907
rect 18604 2864 18656 2873
rect 18696 2907 18748 2916
rect 18696 2873 18705 2907
rect 18705 2873 18739 2907
rect 18739 2873 18748 2907
rect 18696 2864 18748 2873
rect 19892 2864 19944 2916
rect 20076 2864 20128 2916
rect 20628 2864 20680 2916
rect 21732 2907 21784 2916
rect 21732 2873 21741 2907
rect 21741 2873 21775 2907
rect 21775 2873 21784 2907
rect 21732 2864 21784 2873
rect 26148 2864 26200 2916
rect 1216 2796 1268 2848
rect 1676 2796 1728 2848
rect 2504 2839 2556 2848
rect 2504 2805 2513 2839
rect 2513 2805 2547 2839
rect 2547 2805 2556 2839
rect 2504 2796 2556 2805
rect 5172 2796 5224 2848
rect 7564 2796 7616 2848
rect 10692 2796 10744 2848
rect 10876 2796 10928 2848
rect 11060 2796 11112 2848
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 14556 2796 14608 2848
rect 19984 2796 20036 2848
rect 25596 2796 25648 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 204 2592 256 2644
rect 1584 2592 1636 2644
rect 3424 2592 3476 2644
rect 5448 2635 5500 2644
rect 2044 2567 2096 2576
rect 2044 2533 2053 2567
rect 2053 2533 2087 2567
rect 2087 2533 2096 2567
rect 2044 2524 2096 2533
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 9220 2592 9272 2644
rect 5080 2567 5132 2576
rect 664 2456 716 2508
rect 3424 2456 3476 2508
rect 3792 2456 3844 2508
rect 5080 2533 5089 2567
rect 5089 2533 5123 2567
rect 5123 2533 5132 2567
rect 5080 2524 5132 2533
rect 6368 2456 6420 2508
rect 7472 2499 7524 2508
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 7472 2465 7506 2499
rect 7506 2465 7524 2499
rect 7472 2456 7524 2465
rect 10876 2592 10928 2644
rect 11428 2635 11480 2644
rect 11428 2601 11437 2635
rect 11437 2601 11471 2635
rect 11471 2601 11480 2635
rect 11428 2592 11480 2601
rect 14280 2592 14332 2644
rect 13268 2524 13320 2576
rect 19524 2592 19576 2644
rect 22468 2635 22520 2644
rect 14740 2524 14792 2576
rect 10324 2499 10376 2508
rect 10324 2465 10358 2499
rect 10358 2465 10376 2499
rect 10324 2456 10376 2465
rect 11060 2456 11112 2508
rect 1860 2320 1912 2372
rect 4252 2320 4304 2372
rect 5908 2363 5960 2372
rect 5908 2329 5917 2363
rect 5917 2329 5951 2363
rect 5951 2329 5960 2363
rect 5908 2320 5960 2329
rect 16764 2524 16816 2576
rect 18880 2567 18932 2576
rect 18880 2533 18889 2567
rect 18889 2533 18923 2567
rect 18923 2533 18932 2567
rect 18880 2524 18932 2533
rect 15752 2499 15804 2508
rect 15752 2465 15786 2499
rect 15786 2465 15804 2499
rect 15752 2456 15804 2465
rect 16672 2456 16724 2508
rect 22468 2601 22477 2635
rect 22477 2601 22511 2635
rect 22511 2601 22520 2635
rect 22468 2592 22520 2601
rect 23664 2592 23716 2644
rect 25136 2635 25188 2644
rect 20904 2524 20956 2576
rect 25136 2601 25145 2635
rect 25145 2601 25179 2635
rect 25179 2601 25188 2635
rect 25136 2592 25188 2601
rect 8208 2252 8260 2304
rect 8944 2252 8996 2304
rect 12900 2295 12952 2304
rect 12900 2261 12909 2295
rect 12909 2261 12943 2295
rect 12943 2261 12952 2295
rect 12900 2252 12952 2261
rect 13268 2295 13320 2304
rect 13268 2261 13277 2295
rect 13277 2261 13311 2295
rect 13311 2261 13320 2295
rect 13268 2252 13320 2261
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 14740 2252 14792 2304
rect 17408 2252 17460 2304
rect 19064 2388 19116 2440
rect 21548 2456 21600 2508
rect 21916 2456 21968 2508
rect 23756 2456 23808 2508
rect 21732 2431 21784 2440
rect 20076 2320 20128 2372
rect 21732 2397 21741 2431
rect 21741 2397 21775 2431
rect 21775 2397 21784 2431
rect 21732 2388 21784 2397
rect 23480 2388 23532 2440
rect 25412 2431 25464 2440
rect 21364 2320 21416 2372
rect 24032 2320 24084 2372
rect 24768 2320 24820 2372
rect 25412 2397 25421 2431
rect 25421 2397 25455 2431
rect 25455 2397 25464 2431
rect 25412 2388 25464 2397
rect 25596 2431 25648 2440
rect 25596 2397 25605 2431
rect 25605 2397 25639 2431
rect 25639 2397 25648 2431
rect 25596 2388 25648 2397
rect 18420 2295 18472 2304
rect 18420 2261 18429 2295
rect 18429 2261 18463 2295
rect 18463 2261 18472 2295
rect 18420 2252 18472 2261
rect 20168 2295 20220 2304
rect 20168 2261 20177 2295
rect 20177 2261 20211 2295
rect 20211 2261 20220 2295
rect 20168 2252 20220 2261
rect 20904 2295 20956 2304
rect 20904 2261 20913 2295
rect 20913 2261 20947 2295
rect 20947 2261 20956 2295
rect 20904 2252 20956 2261
rect 23664 2252 23716 2304
rect 25228 2252 25280 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 14648 2048 14700 2100
rect 15660 2048 15712 2100
rect 24124 2048 24176 2100
rect 25780 2048 25832 2100
rect 11520 1980 11572 2032
rect 18604 1980 18656 2032
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3054 27520 3110 28000
rect 3606 27520 3662 28000
rect 4158 27520 4214 28000
rect 4710 27520 4766 28000
rect 5262 27520 5318 28000
rect 5814 27520 5870 28000
rect 6366 27520 6422 28000
rect 6918 27520 6974 28000
rect 7562 27520 7618 28000
rect 8114 27520 8170 28000
rect 8666 27520 8722 28000
rect 9218 27520 9274 28000
rect 9770 27520 9826 28000
rect 10322 27520 10378 28000
rect 10874 27520 10930 28000
rect 11426 27520 11482 28000
rect 11978 27520 12034 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 15934 27520 15990 28000
rect 16486 27520 16542 28000
rect 17038 27520 17094 28000
rect 17590 27520 17646 28000
rect 18142 27520 18198 28000
rect 18694 27520 18750 28000
rect 19246 27520 19302 28000
rect 19798 27520 19854 28000
rect 20350 27520 20406 28000
rect 20902 27520 20958 28000
rect 21178 27704 21234 27713
rect 21178 27639 21234 27648
rect 308 25945 336 27520
rect 294 25936 350 25945
rect 294 25871 350 25880
rect 860 25702 888 27520
rect 1122 27024 1178 27033
rect 1122 26959 1178 26968
rect 848 25696 900 25702
rect 848 25638 900 25644
rect 1136 20398 1164 26959
rect 1412 26466 1440 27520
rect 1412 26438 1716 26466
rect 1398 26344 1454 26353
rect 1398 26279 1454 26288
rect 1308 26240 1360 26246
rect 1308 26182 1360 26188
rect 1214 25800 1270 25809
rect 1214 25735 1270 25744
rect 1228 21622 1256 25735
rect 1320 22114 1348 26182
rect 1412 23866 1440 26279
rect 1582 25664 1638 25673
rect 1582 25599 1638 25608
rect 1490 24984 1546 24993
rect 1490 24919 1546 24928
rect 1400 23860 1452 23866
rect 1400 23802 1452 23808
rect 1504 23322 1532 24919
rect 1596 24410 1624 25599
rect 1688 24886 1716 26438
rect 1964 25906 1992 27520
rect 2134 26208 2190 26217
rect 2134 26143 2190 26152
rect 1952 25900 2004 25906
rect 1952 25842 2004 25848
rect 1766 24984 1822 24993
rect 1766 24919 1822 24928
rect 1676 24880 1728 24886
rect 1676 24822 1728 24828
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1582 24304 1638 24313
rect 1582 24239 1638 24248
rect 1492 23316 1544 23322
rect 1492 23258 1544 23264
rect 1596 22710 1624 24239
rect 1780 24018 1808 24919
rect 1688 23990 1808 24018
rect 1584 22704 1636 22710
rect 1584 22646 1636 22652
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 1412 22234 1440 22510
rect 1400 22228 1452 22234
rect 1400 22170 1452 22176
rect 1320 22086 1440 22114
rect 1308 21684 1360 21690
rect 1308 21626 1360 21632
rect 1216 21616 1268 21622
rect 1216 21558 1268 21564
rect 1124 20392 1176 20398
rect 1124 20334 1176 20340
rect 1320 20262 1348 21626
rect 1308 20256 1360 20262
rect 1308 20198 1360 20204
rect 1412 18970 1440 22086
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1492 21616 1544 21622
rect 1492 21558 1544 21564
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1398 18864 1454 18873
rect 1398 18799 1454 18808
rect 1412 18222 1440 18799
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 16833 1440 17614
rect 1398 16824 1454 16833
rect 1398 16759 1454 16768
rect 1400 16040 1452 16046
rect 1398 16008 1400 16017
rect 1452 16008 1454 16017
rect 1398 15943 1454 15952
rect 1398 15600 1454 15609
rect 1398 15535 1400 15544
rect 1452 15535 1454 15544
rect 1400 15506 1452 15512
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12889 1440 13262
rect 1398 12880 1454 12889
rect 1398 12815 1454 12824
rect 1398 12744 1454 12753
rect 1398 12679 1454 12688
rect 1412 12442 1440 12679
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1504 12345 1532 21558
rect 1596 20369 1624 21830
rect 1688 21690 1716 23990
rect 1768 23112 1820 23118
rect 1768 23054 1820 23060
rect 1780 22438 1808 23054
rect 1952 22976 2004 22982
rect 1952 22918 2004 22924
rect 1768 22432 1820 22438
rect 1768 22374 1820 22380
rect 1676 21684 1728 21690
rect 1676 21626 1728 21632
rect 1674 21584 1730 21593
rect 1674 21519 1730 21528
rect 1582 20360 1638 20369
rect 1582 20295 1638 20304
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 18290 1624 20198
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1584 18148 1636 18154
rect 1584 18090 1636 18096
rect 1596 16046 1624 18090
rect 1688 16250 1716 21519
rect 1780 21146 1808 22374
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1872 21350 1900 21966
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1768 20800 1820 20806
rect 1768 20742 1820 20748
rect 1780 20534 1808 20742
rect 1768 20528 1820 20534
rect 1872 20505 1900 21286
rect 1964 21010 1992 22918
rect 2044 22228 2096 22234
rect 2044 22170 2096 22176
rect 2056 21554 2084 22170
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 1952 21004 2004 21010
rect 1952 20946 2004 20952
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1768 20470 1820 20476
rect 1858 20496 1914 20505
rect 1964 20466 1992 20742
rect 1858 20431 1914 20440
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 1766 20360 1822 20369
rect 1766 20295 1822 20304
rect 1860 20324 1912 20330
rect 1780 17134 1808 20295
rect 1860 20266 1912 20272
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1780 15162 1808 16594
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1676 14544 1728 14550
rect 1676 14486 1728 14492
rect 1688 13938 1716 14486
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1688 13530 1716 13874
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1872 13274 1900 20266
rect 1964 20058 1992 20402
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 2056 19281 2084 21082
rect 2148 20262 2176 26143
rect 2516 24449 2544 27520
rect 2686 26072 2742 26081
rect 3068 26042 3096 27520
rect 2686 26007 2742 26016
rect 3056 26036 3108 26042
rect 2700 24993 2728 26007
rect 3056 25978 3108 25984
rect 2686 24984 2742 24993
rect 2686 24919 2742 24928
rect 3068 24857 3096 25978
rect 3620 24857 3648 27520
rect 3054 24848 3110 24857
rect 3054 24783 3110 24792
rect 3606 24848 3662 24857
rect 3606 24783 3662 24792
rect 2502 24440 2558 24449
rect 2502 24375 2558 24384
rect 2228 24268 2280 24274
rect 2228 24210 2280 24216
rect 2240 23526 2268 24210
rect 3698 24168 3754 24177
rect 3698 24103 3754 24112
rect 2594 23624 2650 23633
rect 2594 23559 2650 23568
rect 2228 23520 2280 23526
rect 2228 23462 2280 23468
rect 2412 23520 2464 23526
rect 2412 23462 2464 23468
rect 2240 21554 2268 23462
rect 2424 23225 2452 23462
rect 2410 23216 2466 23225
rect 2410 23151 2466 23160
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2228 21004 2280 21010
rect 2228 20946 2280 20952
rect 2136 20256 2188 20262
rect 2136 20198 2188 20204
rect 2148 20058 2176 20198
rect 2136 20052 2188 20058
rect 2136 19994 2188 20000
rect 2042 19272 2098 19281
rect 2240 19258 2268 20946
rect 2042 19207 2098 19216
rect 2148 19230 2268 19258
rect 1950 19136 2006 19145
rect 1950 19071 2006 19080
rect 1964 16538 1992 19071
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2056 17241 2084 18702
rect 2148 17626 2176 19230
rect 2228 19168 2280 19174
rect 2228 19110 2280 19116
rect 2240 18057 2268 19110
rect 2226 18048 2282 18057
rect 2226 17983 2282 17992
rect 2148 17598 2268 17626
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 2042 17232 2098 17241
rect 2042 17167 2098 17176
rect 2148 16697 2176 17478
rect 2134 16688 2190 16697
rect 2134 16623 2190 16632
rect 1964 16510 2084 16538
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 15978 1992 16390
rect 1952 15972 2004 15978
rect 1952 15914 2004 15920
rect 1964 15706 1992 15914
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1964 15026 1992 15642
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 2056 13802 2084 16510
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 1952 13796 2004 13802
rect 1952 13738 2004 13744
rect 2044 13796 2096 13802
rect 2044 13738 2096 13744
rect 1964 13394 1992 13738
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1872 13246 2084 13274
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1398 11384 1454 11393
rect 1398 11319 1400 11328
rect 1452 11319 1454 11328
rect 1400 11290 1452 11296
rect 1596 11121 1624 11630
rect 1676 11620 1728 11626
rect 1676 11562 1728 11568
rect 1582 11112 1638 11121
rect 1582 11047 1638 11056
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9217 1440 9998
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1216 2848 1268 2854
rect 1216 2790 1268 2796
rect 204 2644 256 2650
rect 204 2586 256 2592
rect 216 480 244 2586
rect 664 2508 716 2514
rect 664 2450 716 2456
rect 676 480 704 2450
rect 1228 480 1256 2790
rect 1412 785 1440 7822
rect 1490 5808 1546 5817
rect 1490 5743 1546 5752
rect 1504 5370 1532 5743
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1596 4049 1624 9046
rect 1688 8537 1716 11562
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1964 10266 1992 10474
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1950 9752 2006 9761
rect 1950 9687 2006 9696
rect 1674 8528 1730 8537
rect 1674 8463 1730 8472
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1688 6662 1716 7210
rect 1766 6760 1822 6769
rect 1766 6695 1822 6704
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 4486 1716 6598
rect 1780 5846 1808 6695
rect 1872 6322 1900 7278
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1964 5914 1992 9687
rect 2056 9110 2084 13246
rect 2148 12866 2176 16458
rect 2240 14890 2268 17598
rect 2332 14958 2360 22918
rect 2424 22273 2452 22918
rect 2410 22264 2466 22273
rect 2410 22199 2466 22208
rect 2504 22092 2556 22098
rect 2504 22034 2556 22040
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2424 21486 2452 21830
rect 2516 21570 2544 22034
rect 2608 21962 2636 23559
rect 3240 23520 3292 23526
rect 3240 23462 3292 23468
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2686 22944 2742 22953
rect 2686 22879 2742 22888
rect 2700 22778 2728 22879
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2792 22438 2820 23122
rect 2964 23044 3016 23050
rect 2964 22986 3016 22992
rect 2872 22500 2924 22506
rect 2872 22442 2924 22448
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2596 21956 2648 21962
rect 2596 21898 2648 21904
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 2516 21542 2636 21570
rect 2412 21480 2464 21486
rect 2412 21422 2464 21428
rect 2424 20369 2452 21422
rect 2608 21350 2636 21542
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 2608 21185 2636 21286
rect 2594 21176 2650 21185
rect 2594 21111 2650 21120
rect 2700 20890 2728 21626
rect 2792 21078 2820 22374
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 2516 20862 2728 20890
rect 2410 20360 2466 20369
rect 2410 20295 2466 20304
rect 2516 20244 2544 20862
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2596 20528 2648 20534
rect 2596 20470 2648 20476
rect 2700 20482 2728 20742
rect 2792 20602 2820 21014
rect 2884 20641 2912 22442
rect 2870 20632 2926 20641
rect 2780 20596 2832 20602
rect 2870 20567 2926 20576
rect 2780 20538 2832 20544
rect 2424 20216 2544 20244
rect 2424 19310 2452 20216
rect 2502 20088 2558 20097
rect 2502 20023 2558 20032
rect 2516 19786 2544 20023
rect 2504 19780 2556 19786
rect 2504 19722 2556 19728
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2608 19242 2636 20470
rect 2700 20454 2820 20482
rect 2792 19922 2820 20454
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19394 2820 19858
rect 2700 19366 2820 19394
rect 2596 19236 2648 19242
rect 2596 19178 2648 19184
rect 2504 19168 2556 19174
rect 2504 19110 2556 19116
rect 2516 17898 2544 19110
rect 2594 17912 2650 17921
rect 2516 17870 2594 17898
rect 2700 17882 2728 19366
rect 2884 18902 2912 19994
rect 2976 19145 3004 22986
rect 3056 22976 3108 22982
rect 3056 22918 3108 22924
rect 3148 22976 3200 22982
rect 3148 22918 3200 22924
rect 3068 22545 3096 22918
rect 3054 22536 3110 22545
rect 3054 22471 3110 22480
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 3068 20806 3096 21830
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 3054 20632 3110 20641
rect 3054 20567 3056 20576
rect 3108 20567 3110 20576
rect 3056 20538 3108 20544
rect 3068 19446 3096 20538
rect 3056 19440 3108 19446
rect 3056 19382 3108 19388
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2962 19136 3018 19145
rect 2962 19071 3018 19080
rect 3068 18986 3096 19246
rect 2976 18958 3096 18986
rect 2872 18896 2924 18902
rect 2872 18838 2924 18844
rect 2872 18760 2924 18766
rect 2870 18728 2872 18737
rect 2924 18728 2926 18737
rect 2870 18663 2926 18672
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2792 18057 2820 18294
rect 2778 18048 2834 18057
rect 2778 17983 2834 17992
rect 2594 17847 2650 17856
rect 2688 17876 2740 17882
rect 2608 17814 2636 17847
rect 2688 17818 2740 17824
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2596 17808 2648 17814
rect 2502 17776 2558 17785
rect 2596 17750 2648 17756
rect 2502 17711 2558 17720
rect 2688 17740 2740 17746
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2424 16794 2452 17274
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2516 16590 2544 17711
rect 2688 17682 2740 17688
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2516 16250 2544 16526
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2608 16182 2636 16662
rect 2700 16522 2728 17682
rect 2792 17066 2820 17818
rect 2872 17808 2924 17814
rect 2872 17750 2924 17756
rect 2884 17134 2912 17750
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2870 16552 2926 16561
rect 2688 16516 2740 16522
rect 2870 16487 2926 16496
rect 2688 16458 2740 16464
rect 2884 16454 2912 16487
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2596 16176 2648 16182
rect 2596 16118 2648 16124
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2502 15736 2558 15745
rect 2502 15671 2558 15680
rect 2516 15434 2544 15671
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 2240 12986 2268 14826
rect 2332 13258 2360 14894
rect 2608 14550 2636 15982
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2700 15162 2728 15438
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2884 14618 2912 14962
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2412 13796 2464 13802
rect 2412 13738 2464 13744
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2148 12838 2268 12866
rect 2134 11248 2190 11257
rect 2134 11183 2190 11192
rect 2148 9654 2176 11183
rect 2240 10538 2268 12838
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2332 12714 2360 12786
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 2332 12442 2360 12650
rect 2424 12646 2452 13738
rect 2778 13560 2834 13569
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2688 13524 2740 13530
rect 2778 13495 2834 13504
rect 2688 13466 2740 13472
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2332 10674 2360 11290
rect 2424 11082 2452 12582
rect 2504 12368 2556 12374
rect 2502 12336 2504 12345
rect 2556 12336 2558 12345
rect 2502 12271 2558 12280
rect 2608 11830 2636 13466
rect 2700 12170 2728 13466
rect 2792 12782 2820 13495
rect 2870 13016 2926 13025
rect 2870 12951 2926 12960
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2792 11898 2820 12718
rect 2884 12617 2912 12951
rect 2870 12608 2926 12617
rect 2870 12543 2926 12552
rect 2976 12458 3004 18958
rect 3056 18896 3108 18902
rect 3056 18838 3108 18844
rect 3068 18426 3096 18838
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3056 18148 3108 18154
rect 3056 18090 3108 18096
rect 3068 17921 3096 18090
rect 3054 17912 3110 17921
rect 3054 17847 3110 17856
rect 3160 17105 3188 22918
rect 3252 20398 3280 23462
rect 3606 23080 3662 23089
rect 3606 23015 3662 23024
rect 3516 22432 3568 22438
rect 3436 22392 3516 22420
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 3344 21078 3372 22034
rect 3332 21072 3384 21078
rect 3332 21014 3384 21020
rect 3332 20936 3384 20942
rect 3330 20904 3332 20913
rect 3384 20904 3386 20913
rect 3330 20839 3386 20848
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3252 19961 3280 20198
rect 3238 19952 3294 19961
rect 3238 19887 3294 19896
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 3252 19174 3280 19790
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3252 18193 3280 18226
rect 3238 18184 3294 18193
rect 3238 18119 3294 18128
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 3146 17096 3202 17105
rect 3056 17060 3108 17066
rect 3146 17031 3202 17040
rect 3056 17002 3108 17008
rect 3068 16794 3096 17002
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3068 15162 3096 15506
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3160 14822 3188 15574
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3068 14278 3096 14418
rect 3160 14414 3188 14758
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3068 14074 3096 14214
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3068 13462 3096 14010
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 3146 13424 3202 13433
rect 3068 12850 3096 13398
rect 3146 13359 3202 13368
rect 3160 13326 3188 13359
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3252 13025 3280 17206
rect 3344 13530 3372 20742
rect 3436 19009 3464 22392
rect 3516 22374 3568 22380
rect 3516 21956 3568 21962
rect 3516 21898 3568 21904
rect 3528 20058 3556 21898
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3422 19000 3478 19009
rect 3422 18935 3478 18944
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3436 16794 3464 18702
rect 3620 18086 3648 23015
rect 3712 21962 3740 24103
rect 3976 23588 4028 23594
rect 3976 23530 4028 23536
rect 3792 23520 3844 23526
rect 3792 23462 3844 23468
rect 3700 21956 3752 21962
rect 3700 21898 3752 21904
rect 3700 21616 3752 21622
rect 3700 21558 3752 21564
rect 3712 20777 3740 21558
rect 3698 20768 3754 20777
rect 3698 20703 3754 20712
rect 3698 20632 3754 20641
rect 3698 20567 3754 20576
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 3514 17912 3570 17921
rect 3620 17882 3648 18022
rect 3514 17847 3516 17856
rect 3568 17847 3570 17856
rect 3608 17876 3660 17882
rect 3516 17818 3568 17824
rect 3608 17818 3660 17824
rect 3712 17762 3740 20567
rect 3804 20058 3832 23462
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 3896 20602 3924 21966
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 3988 20262 4016 23530
rect 4172 23497 4200 27520
rect 4344 26308 4396 26314
rect 4344 26250 4396 26256
rect 4158 23488 4214 23497
rect 4158 23423 4214 23432
rect 4068 22704 4120 22710
rect 4068 22646 4120 22652
rect 4080 21690 4108 22646
rect 4160 22500 4212 22506
rect 4160 22442 4212 22448
rect 4172 22166 4200 22442
rect 4160 22160 4212 22166
rect 4160 22102 4212 22108
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4172 21570 4200 21898
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4080 21542 4200 21570
rect 4080 21418 4108 21542
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 4080 21321 4108 21354
rect 4160 21344 4212 21350
rect 4066 21312 4122 21321
rect 4264 21332 4292 21830
rect 4212 21304 4292 21332
rect 4160 21286 4212 21292
rect 4066 21247 4122 21256
rect 4172 21185 4200 21286
rect 4158 21176 4214 21185
rect 4158 21111 4214 21120
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 4068 20936 4120 20942
rect 4120 20896 4200 20924
rect 4068 20878 4120 20884
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 4080 20534 4108 20742
rect 4172 20602 4200 20896
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 4264 20466 4292 20946
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 3976 20256 4028 20262
rect 4252 20256 4304 20262
rect 4028 20216 4108 20244
rect 3976 20198 4028 20204
rect 3974 20088 4030 20097
rect 3792 20052 3844 20058
rect 3974 20023 4030 20032
rect 3792 19994 3844 20000
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 3804 19009 3832 19382
rect 3790 19000 3846 19009
rect 3896 18970 3924 19654
rect 3790 18935 3846 18944
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 3790 18728 3846 18737
rect 3790 18663 3846 18672
rect 3804 18426 3832 18663
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 3712 17734 3832 17762
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3620 17338 3648 17614
rect 3700 17604 3752 17610
rect 3700 17546 3752 17552
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3422 15464 3478 15473
rect 3422 15399 3478 15408
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3238 13016 3294 13025
rect 3238 12951 3294 12960
rect 3148 12912 3200 12918
rect 3148 12854 3200 12860
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3160 12730 3188 12854
rect 2884 12430 3004 12458
rect 3068 12702 3188 12730
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2792 10826 2820 11698
rect 2700 10810 2820 10826
rect 2688 10804 2820 10810
rect 2740 10798 2820 10804
rect 2688 10746 2740 10752
rect 2884 10724 2912 12430
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2976 12209 3004 12310
rect 2962 12200 3018 12209
rect 2962 12135 3018 12144
rect 2964 11280 3016 11286
rect 2962 11248 2964 11257
rect 3016 11248 3018 11257
rect 2962 11183 3018 11192
rect 3068 11150 3096 12702
rect 3344 12617 3372 13330
rect 3330 12608 3386 12617
rect 3330 12543 3386 12552
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3146 11928 3202 11937
rect 3146 11863 3202 11872
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3054 10976 3110 10985
rect 3054 10911 3110 10920
rect 2792 10696 2912 10724
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2332 10266 2360 10610
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2410 10024 2466 10033
rect 2410 9959 2466 9968
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1952 5908 2004 5914
rect 1872 5868 1952 5896
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1582 4040 1638 4049
rect 1582 3975 1638 3984
rect 1596 2650 1624 3975
rect 1688 3942 1716 4422
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1688 2854 1716 3606
rect 1780 3194 1808 5782
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1398 776 1454 785
rect 1398 711 1454 720
rect 1780 480 1808 2994
rect 1872 2378 1900 5868
rect 1952 5850 2004 5856
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 1964 5234 1992 5578
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 2056 4729 2084 8910
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 2148 7585 2176 8842
rect 2240 8838 2268 9318
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2134 7576 2190 7585
rect 2134 7511 2190 7520
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 2148 5030 2176 6666
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2042 4720 2098 4729
rect 2042 4655 2098 4664
rect 2134 4312 2190 4321
rect 2134 4247 2136 4256
rect 2188 4247 2190 4256
rect 2136 4218 2188 4224
rect 2240 4162 2268 8774
rect 2424 8634 2452 9959
rect 2516 9518 2544 10202
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2700 9722 2728 9998
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2608 9178 2636 9522
rect 2792 9353 2820 10696
rect 3068 10305 3096 10911
rect 3054 10296 3110 10305
rect 3054 10231 3110 10240
rect 2964 10192 3016 10198
rect 2870 10160 2926 10169
rect 3016 10152 3096 10180
rect 2964 10134 3016 10140
rect 2870 10095 2926 10104
rect 2778 9344 2834 9353
rect 2778 9279 2834 9288
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2686 9072 2742 9081
rect 2686 9007 2742 9016
rect 2700 8974 2728 9007
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2412 8628 2464 8634
rect 2700 8616 2728 8910
rect 2792 8906 2820 9279
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2464 8588 2544 8616
rect 2412 8570 2464 8576
rect 2318 7984 2374 7993
rect 2318 7919 2374 7928
rect 2332 4554 2360 7919
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7274 2452 7686
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2516 7154 2544 8588
rect 2608 8588 2728 8616
rect 2608 8498 2636 8588
rect 2884 8498 2912 10095
rect 3068 9926 3096 10152
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2962 9480 3018 9489
rect 2962 9415 3018 9424
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2608 8294 2636 8434
rect 2596 8288 2648 8294
rect 2884 8242 2912 8434
rect 2596 8230 2648 8236
rect 2792 8214 2912 8242
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2424 7126 2544 7154
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2148 4134 2268 4162
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2056 3398 2084 3878
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2056 2922 2084 3334
rect 2044 2916 2096 2922
rect 2044 2858 2096 2864
rect 2056 2582 2084 2858
rect 2044 2576 2096 2582
rect 2044 2518 2096 2524
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 2148 1329 2176 4134
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2134 1320 2190 1329
rect 2134 1255 2190 1264
rect 2240 480 2268 4014
rect 2332 4010 2360 4490
rect 2424 4078 2452 7126
rect 2502 6896 2558 6905
rect 2608 6866 2636 7890
rect 2792 7818 2820 8214
rect 2870 8120 2926 8129
rect 2870 8055 2926 8064
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2502 6831 2558 6840
rect 2596 6860 2648 6866
rect 2516 6730 2544 6831
rect 2596 6802 2648 6808
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2516 5914 2544 6190
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2516 5370 2544 5850
rect 2608 5642 2636 6598
rect 2700 6338 2728 7210
rect 2884 6798 2912 8055
rect 2976 8022 3004 9415
rect 3068 9382 3096 9862
rect 3160 9654 3188 11863
rect 3252 11354 3280 12378
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3344 11694 3372 12174
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3344 11354 3372 11630
rect 3436 11626 3464 15399
rect 3528 12186 3556 17070
rect 3620 17066 3648 17274
rect 3608 17060 3660 17066
rect 3608 17002 3660 17008
rect 3712 16998 3740 17546
rect 3700 16992 3752 16998
rect 3606 16960 3662 16969
rect 3700 16934 3752 16940
rect 3606 16895 3662 16904
rect 3620 15065 3648 16895
rect 3606 15056 3662 15065
rect 3606 14991 3662 15000
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3620 12442 3648 12786
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3528 12158 3648 12186
rect 3514 11792 3570 11801
rect 3514 11727 3570 11736
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 10810 3280 11154
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3238 10704 3294 10713
rect 3238 10639 3294 10648
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 8838 3096 9318
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3160 8566 3188 8842
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 3160 8401 3188 8502
rect 3146 8392 3202 8401
rect 3056 8356 3108 8362
rect 3146 8327 3202 8336
rect 3056 8298 3108 8304
rect 3068 8090 3096 8298
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2976 7546 3004 7958
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 3160 7426 3188 8327
rect 2976 7398 3188 7426
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2700 6310 2912 6338
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2792 5681 2820 5714
rect 2778 5672 2834 5681
rect 2596 5636 2648 5642
rect 2778 5607 2834 5616
rect 2596 5578 2648 5584
rect 2884 5386 2912 6310
rect 2976 6100 3004 7398
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3068 6798 3096 7142
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3068 6254 3096 6734
rect 3146 6352 3202 6361
rect 3146 6287 3202 6296
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2976 6072 3096 6100
rect 2964 5704 3016 5710
rect 2962 5672 2964 5681
rect 3016 5672 3018 5681
rect 2962 5607 3018 5616
rect 2504 5364 2556 5370
rect 2884 5358 3004 5386
rect 2504 5306 2556 5312
rect 2516 4826 2544 5306
rect 2976 5234 3004 5358
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2688 5092 2740 5098
rect 2688 5034 2740 5040
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 2516 3466 2544 4558
rect 2700 4146 2728 5034
rect 2976 5030 3004 5170
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2962 4856 3018 4865
rect 2962 4791 3018 4800
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2870 3904 2926 3913
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2516 2854 2544 2994
rect 2504 2848 2556 2854
rect 2502 2816 2504 2825
rect 2556 2816 2558 2825
rect 2502 2751 2558 2760
rect 2792 480 2820 3878
rect 2870 3839 2926 3848
rect 2884 3670 2912 3839
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2976 2990 3004 4791
rect 3068 3126 3096 6072
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2964 2440 3016 2446
rect 2962 2408 2964 2417
rect 3016 2408 3018 2417
rect 2962 2343 3018 2352
rect 3160 2009 3188 6287
rect 3252 6254 3280 10639
rect 3344 9081 3372 11086
rect 3436 9994 3464 11562
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3528 9489 3556 11727
rect 3514 9480 3570 9489
rect 3514 9415 3570 9424
rect 3330 9072 3386 9081
rect 3330 9007 3386 9016
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3436 7206 3464 8026
rect 3516 7744 3568 7750
rect 3514 7712 3516 7721
rect 3568 7712 3570 7721
rect 3514 7647 3570 7656
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 5574 3280 6054
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 5166 3280 5510
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3252 4282 3280 4966
rect 3344 4622 3372 5850
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3252 3942 3280 4218
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3238 3768 3294 3777
rect 3238 3703 3294 3712
rect 3252 3058 3280 3703
rect 3332 3528 3384 3534
rect 3436 3505 3464 6190
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3528 4214 3556 4694
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3620 4146 3648 12158
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3332 3470 3384 3476
rect 3422 3496 3478 3505
rect 3344 3194 3372 3470
rect 3422 3431 3478 3440
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3146 2000 3202 2009
rect 3146 1935 3202 1944
rect 3344 480 3372 3130
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3436 2650 3464 3062
rect 3528 2922 3556 3334
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3422 2544 3478 2553
rect 3422 2479 3424 2488
rect 3476 2479 3478 2488
rect 3424 2450 3476 2456
rect 3712 2394 3740 16934
rect 3804 15026 3832 17734
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 3896 16794 3924 17138
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3988 16726 4016 20023
rect 4080 19514 4108 20216
rect 4252 20198 4304 20204
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4160 19304 4212 19310
rect 4158 19272 4160 19281
rect 4212 19272 4214 19281
rect 4158 19207 4214 19216
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4080 18902 4108 19110
rect 4068 18896 4120 18902
rect 4068 18838 4120 18844
rect 4066 18320 4122 18329
rect 4066 18255 4122 18264
rect 3976 16720 4028 16726
rect 4080 16697 4108 18255
rect 4264 16998 4292 20198
rect 4356 17338 4384 26250
rect 4724 26178 4752 27520
rect 4712 26172 4764 26178
rect 4712 26114 4764 26120
rect 5276 24698 5304 27520
rect 5828 25265 5856 27520
rect 6276 25424 6328 25430
rect 6276 25366 6328 25372
rect 5814 25256 5870 25265
rect 5814 25191 5870 25200
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6092 24948 6144 24954
rect 6092 24890 6144 24896
rect 5276 24670 5488 24698
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 4620 23656 4672 23662
rect 4620 23598 4672 23604
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4448 20913 4476 21830
rect 4540 21593 4568 22918
rect 4526 21584 4582 21593
rect 4526 21519 4582 21528
rect 4528 21412 4580 21418
rect 4528 21354 4580 21360
rect 4434 20904 4490 20913
rect 4434 20839 4490 20848
rect 4436 20800 4488 20806
rect 4436 20742 4488 20748
rect 4448 18834 4476 20742
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4448 18086 4476 18566
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4356 16776 4384 17274
rect 4264 16748 4384 16776
rect 3976 16662 4028 16668
rect 4066 16688 4122 16697
rect 4066 16623 4122 16632
rect 4264 16572 4292 16748
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4080 16544 4292 16572
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15706 3924 15846
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3804 13977 3832 14826
rect 3790 13968 3846 13977
rect 3790 13903 3846 13912
rect 3896 13852 3924 14826
rect 3988 14074 4016 15506
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3804 13824 3924 13852
rect 3804 12646 3832 13824
rect 3988 13802 4016 14010
rect 3976 13796 4028 13802
rect 3896 13756 3976 13784
rect 3896 12850 3924 13756
rect 3976 13738 4028 13744
rect 4080 13394 4108 16544
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4264 16250 4292 16390
rect 4252 16244 4304 16250
rect 4172 16204 4252 16232
rect 4172 16046 4200 16204
rect 4252 16186 4304 16192
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4250 16008 4306 16017
rect 4172 15638 4200 15982
rect 4356 15978 4384 16594
rect 4250 15943 4306 15952
rect 4344 15972 4396 15978
rect 4264 15706 4292 15943
rect 4344 15914 4396 15920
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 4344 15632 4396 15638
rect 4344 15574 4396 15580
rect 4356 15162 4384 15574
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4342 14648 4398 14657
rect 4342 14583 4398 14592
rect 4356 14550 4384 14583
rect 4344 14544 4396 14550
rect 4344 14486 4396 14492
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 4172 13841 4200 14282
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4158 13832 4214 13841
rect 4158 13767 4214 13776
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 4066 13152 4122 13161
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3882 12608 3938 12617
rect 3882 12543 3938 12552
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 9761 3832 12038
rect 3790 9752 3846 9761
rect 3790 9687 3846 9696
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3804 9489 3832 9522
rect 3896 9518 3924 12543
rect 3884 9512 3936 9518
rect 3790 9480 3846 9489
rect 3884 9454 3936 9460
rect 3790 9415 3846 9424
rect 3896 9178 3924 9454
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3884 8356 3936 8362
rect 3988 8344 4016 13126
rect 4066 13087 4122 13096
rect 4080 12714 4108 13087
rect 4172 12986 4200 13767
rect 4264 13705 4292 14214
rect 4250 13696 4306 13705
rect 4250 13631 4306 13640
rect 4344 13320 4396 13326
rect 4342 13288 4344 13297
rect 4396 13288 4398 13297
rect 4342 13223 4398 13232
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4448 12832 4476 17614
rect 4172 12804 4476 12832
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 4066 12336 4122 12345
rect 4066 12271 4122 12280
rect 4080 11762 4108 12271
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4080 9738 4108 10202
rect 4172 9926 4200 12804
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4080 9710 4200 9738
rect 4172 9586 4200 9710
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4172 9178 4200 9318
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4264 8634 4292 12650
rect 4434 12608 4490 12617
rect 4434 12543 4490 12552
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4356 11880 4384 12378
rect 4448 12170 4476 12543
rect 4436 12164 4488 12170
rect 4436 12106 4488 12112
rect 4436 11892 4488 11898
rect 4356 11852 4436 11880
rect 4436 11834 4488 11840
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4356 11354 4384 11630
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4356 10266 4384 11290
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4356 10062 4384 10202
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4356 8906 4384 9522
rect 4434 9208 4490 9217
rect 4434 9143 4490 9152
rect 4448 9110 4476 9143
rect 4436 9104 4488 9110
rect 4436 9046 4488 9052
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4448 8634 4476 9046
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 3936 8316 4016 8344
rect 3884 8298 3936 8304
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3804 7002 3832 8230
rect 3988 7818 4016 8316
rect 4080 8129 4108 8502
rect 4264 8430 4292 8570
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 4356 7750 4384 8298
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4356 7410 4384 7686
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3804 2514 3832 6938
rect 3882 5264 3938 5273
rect 3882 5199 3938 5208
rect 3896 4457 3924 5199
rect 3988 5001 4016 7278
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4068 6656 4120 6662
rect 4172 6644 4200 7210
rect 4356 6662 4384 7346
rect 4448 7206 4476 7958
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4344 6656 4396 6662
rect 4120 6616 4292 6644
rect 4068 6598 4120 6604
rect 4158 5944 4214 5953
rect 4158 5879 4214 5888
rect 3974 4992 4030 5001
rect 3974 4927 4030 4936
rect 4172 4690 4200 5879
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3882 4448 3938 4457
rect 3882 4383 3938 4392
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3896 3602 3924 4082
rect 3988 4010 4016 4558
rect 4172 4486 4200 4626
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4080 4162 4108 4422
rect 4080 4134 4200 4162
rect 4172 4078 4200 4134
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3602 4108 3878
rect 4172 3738 4200 4014
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3896 3194 3924 3538
rect 4080 3194 4108 3538
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3712 2366 3832 2394
rect 3698 2272 3754 2281
rect 3698 2207 3754 2216
rect 3712 1057 3740 2207
rect 3804 1601 3832 2366
rect 3790 1592 3846 1601
rect 3790 1527 3846 1536
rect 3698 1048 3754 1057
rect 3698 983 3754 992
rect 3896 626 3924 3130
rect 4264 2378 4292 6616
rect 4344 6598 4396 6604
rect 4356 4554 4384 6598
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4342 4176 4398 4185
rect 4342 4111 4398 4120
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 3896 598 4016 626
rect 3896 480 3924 598
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2226 0 2282 480
rect 2778 0 2834 480
rect 3330 0 3386 480
rect 3882 0 3938 480
rect 3988 105 4016 598
rect 4356 480 4384 4111
rect 4448 3641 4476 7142
rect 4540 3670 4568 21354
rect 4632 16046 4660 23598
rect 4724 22030 4752 24550
rect 5172 24200 5224 24206
rect 5172 24142 5224 24148
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4710 21856 4766 21865
rect 4710 21791 4766 21800
rect 4724 17678 4752 21791
rect 4816 18698 4844 23530
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4724 17134 4752 17478
rect 4816 17202 4844 18634
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4802 17096 4858 17105
rect 4802 17031 4804 17040
rect 4856 17031 4858 17040
rect 4804 17002 4856 17008
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4632 15434 4660 15982
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4724 15314 4752 16934
rect 4816 16250 4844 17002
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4632 15286 4752 15314
rect 4632 13802 4660 15286
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4724 14618 4752 15030
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4724 14278 4752 14418
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4618 13560 4674 13569
rect 4618 13495 4674 13504
rect 4632 12374 4660 13495
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4632 11665 4660 12106
rect 4618 11656 4674 11665
rect 4618 11591 4674 11600
rect 4724 11529 4752 14214
rect 4816 13433 4844 16050
rect 4908 15706 4936 23462
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 5000 22642 5028 23122
rect 5080 23112 5132 23118
rect 5080 23054 5132 23060
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 4986 21992 5042 22001
rect 4986 21927 4988 21936
rect 5040 21927 5042 21936
rect 4988 21898 5040 21904
rect 4988 21140 5040 21146
rect 4988 21082 5040 21088
rect 5000 20262 5028 21082
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 5000 19378 5028 19790
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 5000 18970 5028 19314
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 5000 16114 5028 18770
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 4908 14346 4936 15642
rect 5000 14414 5028 15846
rect 5092 14958 5120 23054
rect 5184 21418 5212 24142
rect 5172 21412 5224 21418
rect 5172 21354 5224 21360
rect 5276 21332 5304 24550
rect 5356 24132 5408 24138
rect 5356 24074 5408 24080
rect 5368 21434 5396 24074
rect 5460 23497 5488 24670
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5446 23488 5502 23497
rect 5446 23423 5502 23432
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5460 22642 5488 22918
rect 5448 22636 5500 22642
rect 5448 22578 5500 22584
rect 5552 22488 5580 24550
rect 6104 24410 6132 24890
rect 6092 24404 6144 24410
rect 6092 24346 6144 24352
rect 6184 24200 6236 24206
rect 6184 24142 6236 24148
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5630 23352 5686 23361
rect 5630 23287 5632 23296
rect 5684 23287 5686 23296
rect 5632 23258 5684 23264
rect 6092 22976 6144 22982
rect 6092 22918 6144 22924
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5632 22568 5684 22574
rect 5632 22510 5684 22516
rect 5460 22460 5580 22488
rect 5460 22234 5488 22460
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5460 21690 5488 22170
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5552 21622 5580 21966
rect 5644 21962 5672 22510
rect 5724 22432 5776 22438
rect 5722 22400 5724 22409
rect 5776 22400 5778 22409
rect 5722 22335 5778 22344
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21672 6040 21830
rect 5828 21644 6040 21672
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5368 21406 5488 21434
rect 5356 21344 5408 21350
rect 5276 21304 5356 21332
rect 5356 21286 5408 21292
rect 5264 21072 5316 21078
rect 5264 21014 5316 21020
rect 5276 20398 5304 21014
rect 5368 20534 5396 21286
rect 5460 21078 5488 21406
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 5448 21072 5500 21078
rect 5448 21014 5500 21020
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5460 20602 5488 20878
rect 5448 20596 5500 20602
rect 5448 20538 5500 20544
rect 5356 20528 5408 20534
rect 5552 20482 5580 21354
rect 5644 20913 5672 21490
rect 5828 21418 5856 21644
rect 5998 21448 6054 21457
rect 5816 21412 5868 21418
rect 5998 21383 6000 21392
rect 5816 21354 5868 21360
rect 6052 21383 6054 21392
rect 6000 21354 6052 21360
rect 5828 21010 5856 21354
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 6000 20936 6052 20942
rect 5630 20904 5686 20913
rect 6000 20878 6052 20884
rect 5630 20839 5686 20848
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5356 20470 5408 20476
rect 5460 20454 5580 20482
rect 5630 20496 5686 20505
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 5184 19242 5212 19926
rect 5276 19514 5304 19994
rect 5368 19514 5396 20266
rect 5460 19786 5488 20454
rect 6012 20466 6040 20878
rect 5630 20431 5686 20440
rect 6000 20460 6052 20466
rect 5540 19916 5592 19922
rect 5644 19904 5672 20431
rect 6000 20402 6052 20408
rect 6104 20346 6132 22918
rect 6196 21894 6224 24142
rect 6288 23866 6316 25366
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6276 23588 6328 23594
rect 6276 23530 6328 23536
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 5908 20324 5960 20330
rect 5908 20266 5960 20272
rect 6012 20318 6132 20346
rect 5920 19922 5948 20266
rect 5592 19876 5672 19904
rect 5908 19916 5960 19922
rect 5540 19858 5592 19864
rect 5908 19858 5960 19864
rect 5448 19780 5500 19786
rect 5448 19722 5500 19728
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5552 19310 5580 19858
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5540 19304 5592 19310
rect 5262 19272 5318 19281
rect 5172 19236 5224 19242
rect 5262 19207 5318 19216
rect 5368 19264 5540 19292
rect 5172 19178 5224 19184
rect 5276 18902 5304 19207
rect 5264 18896 5316 18902
rect 5264 18838 5316 18844
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5184 17814 5212 18362
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 5184 17338 5212 17750
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5184 16454 5212 17274
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5276 15960 5304 18226
rect 5184 15932 5304 15960
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5184 14906 5212 15932
rect 5368 15858 5396 19264
rect 5540 19246 5592 19252
rect 6012 19224 6040 20318
rect 6196 20262 6224 21830
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6092 19984 6144 19990
rect 6092 19926 6144 19932
rect 6104 19378 6132 19926
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6012 19196 6132 19224
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5998 19136 6054 19145
rect 5448 18896 5500 18902
rect 5448 18838 5500 18844
rect 5460 18358 5488 18838
rect 5920 18834 5948 19110
rect 5998 19071 6054 19080
rect 6012 18970 6040 19071
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6012 18873 6040 18906
rect 5998 18864 6054 18873
rect 5908 18828 5960 18834
rect 5998 18799 6054 18808
rect 5908 18770 5960 18776
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5460 17202 5488 18090
rect 5552 18086 5580 18702
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17746 5580 18022
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5460 16794 5488 17138
rect 5552 16998 5580 17682
rect 6000 17604 6052 17610
rect 6000 17546 6052 17552
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 5644 17105 5672 17206
rect 5630 17096 5686 17105
rect 5630 17031 5686 17040
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5276 15830 5396 15858
rect 5276 15502 5304 15830
rect 5460 15706 5488 16730
rect 5552 16114 5580 16934
rect 6012 16726 6040 17546
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5448 15700 5500 15706
rect 5368 15660 5448 15688
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5276 15094 5304 15438
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 5368 15026 5396 15660
rect 5448 15642 5500 15648
rect 5448 15156 5500 15162
rect 5552 15144 5580 15914
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5500 15116 5580 15144
rect 5448 15098 5500 15104
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 4896 14340 4948 14346
rect 4896 14282 4948 14288
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4802 13424 4858 13433
rect 4802 13359 4858 13368
rect 4816 12617 4844 13359
rect 4802 12608 4858 12617
rect 4802 12543 4858 12552
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4816 11937 4844 12310
rect 4802 11928 4858 11937
rect 4802 11863 4858 11872
rect 4710 11520 4766 11529
rect 4710 11455 4766 11464
rect 4908 11370 4936 14010
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 4724 11342 4936 11370
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4632 10130 4660 10474
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4632 9722 4660 10066
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4724 9654 4752 11342
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4816 10470 4844 11154
rect 5000 10849 5028 13738
rect 5092 13326 5120 14894
rect 5184 14878 5304 14906
rect 5172 14816 5224 14822
rect 5170 14784 5172 14793
rect 5224 14784 5226 14793
rect 5170 14719 5226 14728
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5092 12918 5120 13126
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4986 10840 5042 10849
rect 4986 10775 5042 10784
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4894 10432 4950 10441
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4618 9208 4674 9217
rect 4618 9143 4674 9152
rect 4632 8498 4660 9143
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 8362 4660 8434
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4632 7342 4660 7822
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4632 5846 4660 6190
rect 4620 5840 4672 5846
rect 4620 5782 4672 5788
rect 4632 5370 4660 5782
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4618 5128 4674 5137
rect 4618 5063 4674 5072
rect 4632 4622 4660 5063
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4724 4162 4752 8774
rect 4816 7449 4844 10406
rect 4894 10367 4950 10376
rect 4908 9994 4936 10367
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4908 8022 4936 9590
rect 5000 9178 5028 10775
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5000 8566 5028 9114
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5092 8090 5120 12582
rect 5184 11665 5212 14554
rect 5276 14074 5304 14878
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5460 13530 5488 14486
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5460 13433 5488 13466
rect 5446 13424 5502 13433
rect 5552 13394 5580 13670
rect 5920 13462 5948 13942
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 5446 13359 5502 13368
rect 5540 13388 5592 13394
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5262 12880 5318 12889
rect 5262 12815 5318 12824
rect 5276 12714 5304 12815
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5276 12442 5304 12650
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5170 11656 5226 11665
rect 5170 11591 5226 11600
rect 5172 11008 5224 11014
rect 5276 10985 5304 11698
rect 5172 10950 5224 10956
rect 5262 10976 5318 10985
rect 5184 10713 5212 10950
rect 5262 10911 5318 10920
rect 5170 10704 5226 10713
rect 5170 10639 5226 10648
rect 5184 10198 5212 10639
rect 5262 10568 5318 10577
rect 5262 10503 5318 10512
rect 5276 10266 5304 10503
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 9518 5212 9998
rect 5264 9648 5316 9654
rect 5262 9616 5264 9625
rect 5316 9616 5318 9625
rect 5262 9551 5318 9560
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5262 9072 5318 9081
rect 5262 9007 5318 9016
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4894 7848 4950 7857
rect 4894 7783 4950 7792
rect 4908 7546 4936 7783
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4802 7440 4858 7449
rect 4802 7375 4858 7384
rect 4908 6934 4936 7482
rect 5092 7342 5120 8026
rect 5276 7954 5304 9007
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4986 7168 5042 7177
rect 4986 7103 5042 7112
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4816 6225 4844 6598
rect 5000 6390 5028 7103
rect 5170 7032 5226 7041
rect 5170 6967 5226 6976
rect 5078 6896 5134 6905
rect 5078 6831 5134 6840
rect 4988 6384 5040 6390
rect 5092 6361 5120 6831
rect 4988 6326 5040 6332
rect 5078 6352 5134 6361
rect 4802 6216 4858 6225
rect 4802 6151 4858 6160
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 5030 4844 5510
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 5000 4321 5028 6326
rect 5078 6287 5134 6296
rect 5184 6186 5212 6967
rect 5264 6792 5316 6798
rect 5368 6780 5396 13194
rect 5460 12306 5488 13359
rect 5540 13330 5592 13336
rect 5552 12374 5580 13330
rect 5920 13258 5948 13398
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 13025 6040 16390
rect 6104 15978 6132 19196
rect 6196 17814 6224 19314
rect 6288 18902 6316 23530
rect 6380 22273 6408 27520
rect 6932 25974 6960 27520
rect 7576 26722 7604 27520
rect 7564 26716 7616 26722
rect 7564 26658 7616 26664
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 6920 25968 6972 25974
rect 6920 25910 6972 25916
rect 6460 25288 6512 25294
rect 6460 25230 6512 25236
rect 6472 24410 6500 25230
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 6552 24064 6604 24070
rect 6552 24006 6604 24012
rect 6564 23633 6592 24006
rect 6550 23624 6606 23633
rect 6550 23559 6606 23568
rect 6552 23248 6604 23254
rect 6552 23190 6604 23196
rect 6458 23080 6514 23089
rect 6458 23015 6514 23024
rect 6472 22982 6500 23015
rect 6460 22976 6512 22982
rect 6460 22918 6512 22924
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 6366 22264 6422 22273
rect 6472 22250 6500 22578
rect 6564 22438 6592 23190
rect 6552 22432 6604 22438
rect 6550 22400 6552 22409
rect 6604 22400 6606 22409
rect 6550 22335 6606 22344
rect 6472 22222 6592 22250
rect 6366 22199 6422 22208
rect 6458 22128 6514 22137
rect 6458 22063 6514 22072
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 6380 20806 6408 21898
rect 6472 21146 6500 22063
rect 6460 21140 6512 21146
rect 6460 21082 6512 21088
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6472 20262 6500 20402
rect 6460 20256 6512 20262
rect 6460 20198 6512 20204
rect 6472 19922 6500 20198
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6276 18896 6328 18902
rect 6276 18838 6328 18844
rect 6276 18692 6328 18698
rect 6276 18634 6328 18640
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6196 16726 6224 17478
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6196 16250 6224 16662
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6288 15858 6316 18634
rect 6380 18222 6408 19178
rect 6472 18902 6500 19450
rect 6460 18896 6512 18902
rect 6460 18838 6512 18844
rect 6472 18426 6500 18838
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6564 17320 6592 22222
rect 6656 22001 6684 25094
rect 6932 24818 6960 25910
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7194 25120 7250 25129
rect 7194 25055 7250 25064
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6736 24744 6788 24750
rect 6736 24686 6788 24692
rect 7010 24712 7066 24721
rect 6748 23769 6776 24686
rect 7010 24647 7066 24656
rect 7104 24676 7156 24682
rect 7024 24614 7052 24647
rect 7104 24618 7156 24624
rect 7012 24608 7064 24614
rect 7012 24550 7064 24556
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6734 23760 6790 23769
rect 6734 23695 6790 23704
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6642 21992 6698 22001
rect 6642 21927 6698 21936
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6656 20942 6684 21286
rect 6644 20936 6696 20942
rect 6644 20878 6696 20884
rect 6656 20330 6684 20878
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6656 19242 6684 19858
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6644 18624 6696 18630
rect 6644 18566 6696 18572
rect 6656 18193 6684 18566
rect 6642 18184 6698 18193
rect 6642 18119 6698 18128
rect 6642 17776 6698 17785
rect 6642 17711 6698 17720
rect 6656 17377 6684 17711
rect 6196 15830 6316 15858
rect 6380 17292 6592 17320
rect 6642 17368 6698 17377
rect 6642 17303 6698 17312
rect 6196 15570 6224 15830
rect 6380 15722 6408 17292
rect 6748 17218 6776 23462
rect 6840 23225 6868 24006
rect 6932 23594 6960 24210
rect 7010 24032 7066 24041
rect 7010 23967 7066 23976
rect 6920 23588 6972 23594
rect 6920 23530 6972 23536
rect 6826 23216 6882 23225
rect 7024 23202 7052 23967
rect 6932 23186 7052 23202
rect 6826 23151 6882 23160
rect 6920 23180 7052 23186
rect 6972 23174 7052 23180
rect 6920 23122 6972 23128
rect 6828 23044 6880 23050
rect 6828 22986 6880 22992
rect 6840 19281 6868 22986
rect 6932 22778 6960 23122
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6932 22574 6960 22714
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 7024 22522 7052 23054
rect 7116 22642 7144 24618
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7024 22494 7144 22522
rect 7116 22438 7144 22494
rect 7104 22432 7156 22438
rect 7102 22400 7104 22409
rect 7156 22400 7158 22409
rect 7102 22335 7158 22344
rect 7208 22166 7236 25055
rect 7300 24410 7328 25842
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7288 24404 7340 24410
rect 7288 24346 7340 24352
rect 7484 24177 7512 24550
rect 7470 24168 7526 24177
rect 7470 24103 7526 24112
rect 7576 24018 7604 26522
rect 7748 26104 7800 26110
rect 7748 26046 7800 26052
rect 7760 25498 7788 26046
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 7748 25356 7800 25362
rect 7748 25298 7800 25304
rect 7654 25256 7710 25265
rect 7654 25191 7710 25200
rect 7484 23990 7604 24018
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7288 23044 7340 23050
rect 7288 22986 7340 22992
rect 7196 22160 7248 22166
rect 7116 22120 7196 22148
rect 7012 22024 7064 22030
rect 6918 21992 6974 22001
rect 7012 21966 7064 21972
rect 6918 21927 6974 21936
rect 6932 21486 6960 21927
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 7024 21418 7052 21966
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 7024 21321 7052 21354
rect 7010 21312 7066 21321
rect 7010 21247 7066 21256
rect 7116 21146 7144 22120
rect 7196 22102 7248 22108
rect 7300 22098 7328 22986
rect 7288 22092 7340 22098
rect 7288 22034 7340 22040
rect 7196 21412 7248 21418
rect 7196 21354 7248 21360
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7208 21049 7236 21354
rect 7010 21040 7066 21049
rect 7010 20975 7066 20984
rect 7194 21040 7250 21049
rect 7194 20975 7250 20984
rect 7288 21004 7340 21010
rect 7024 19514 7052 20975
rect 7288 20946 7340 20952
rect 7102 20904 7158 20913
rect 7102 20839 7158 20848
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6932 19292 6960 19382
rect 6932 19281 7052 19292
rect 6826 19272 6882 19281
rect 6932 19272 7066 19281
rect 6932 19264 7010 19272
rect 6826 19207 6882 19216
rect 7010 19207 7066 19216
rect 6840 18306 6868 19207
rect 7024 18873 7052 19207
rect 7010 18864 7066 18873
rect 7010 18799 7066 18808
rect 7116 18442 7144 20839
rect 7194 20088 7250 20097
rect 7300 20058 7328 20946
rect 7392 20097 7420 23530
rect 7378 20088 7434 20097
rect 7194 20023 7250 20032
rect 7288 20052 7340 20058
rect 7208 19553 7236 20023
rect 7378 20023 7434 20032
rect 7288 19994 7340 20000
rect 7194 19544 7250 19553
rect 7194 19479 7250 19488
rect 7194 19000 7250 19009
rect 7194 18935 7250 18944
rect 7208 18834 7236 18935
rect 7288 18896 7340 18902
rect 7288 18838 7340 18844
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7024 18414 7144 18442
rect 6840 18278 6960 18306
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 6840 17882 6868 18090
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6840 17785 6868 17818
rect 6826 17776 6882 17785
rect 6826 17711 6882 17720
rect 6932 17338 6960 18278
rect 7024 17746 7052 18414
rect 7208 18306 7236 18770
rect 7116 18278 7236 18306
rect 7116 17882 7144 18278
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 6288 15694 6408 15722
rect 6564 17190 6776 17218
rect 6460 15700 6512 15706
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6092 15360 6144 15366
rect 6090 15328 6092 15337
rect 6144 15328 6146 15337
rect 6090 15263 6146 15272
rect 6196 14793 6224 15506
rect 6182 14784 6238 14793
rect 6182 14719 6238 14728
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6104 13734 6132 14418
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6104 13569 6132 13670
rect 6090 13560 6146 13569
rect 6090 13495 6146 13504
rect 6196 13326 6224 14350
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 5998 13016 6054 13025
rect 5998 12951 6054 12960
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6012 12442 6040 12650
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 11830 5488 12038
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5460 11082 5488 11562
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5460 9042 5488 11018
rect 5552 10810 5580 12310
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5906 11384 5962 11393
rect 5906 11319 5908 11328
rect 5960 11319 5962 11328
rect 5908 11290 5960 11296
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5538 10296 5594 10305
rect 5644 10266 5672 10542
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5538 10231 5594 10240
rect 5632 10260 5684 10266
rect 5552 9178 5580 10231
rect 5632 10202 5684 10208
rect 5920 10062 5948 10406
rect 5724 10056 5776 10062
rect 5722 10024 5724 10033
rect 5908 10056 5960 10062
rect 5776 10024 5778 10033
rect 5908 9998 5960 10004
rect 5722 9959 5778 9968
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5644 8974 5672 9454
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5446 8528 5502 8537
rect 5446 8463 5502 8472
rect 5460 8430 5488 8463
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5552 7993 5580 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5538 7984 5594 7993
rect 5538 7919 5594 7928
rect 5540 7744 5592 7750
rect 5446 7712 5502 7721
rect 5502 7692 5540 7698
rect 5502 7686 5592 7692
rect 5502 7670 5580 7686
rect 5446 7647 5502 7656
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5316 6752 5396 6780
rect 5460 6769 5488 6802
rect 5552 6798 5580 7670
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5540 6792 5592 6798
rect 5446 6760 5502 6769
rect 5264 6734 5316 6740
rect 5540 6734 5592 6740
rect 5446 6695 5502 6704
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 4978 5120 6054
rect 5184 5817 5212 6122
rect 5170 5808 5226 5817
rect 5170 5743 5226 5752
rect 5460 5166 5488 6394
rect 5552 6118 5580 6734
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5552 5166 5580 6054
rect 5920 5817 5948 6054
rect 5906 5808 5962 5817
rect 5906 5743 5962 5752
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5092 4950 5212 4978
rect 5078 4856 5134 4865
rect 5078 4791 5080 4800
rect 5132 4791 5134 4800
rect 5080 4762 5132 4768
rect 4986 4312 5042 4321
rect 4986 4247 5042 4256
rect 4724 4134 4844 4162
rect 4528 3664 4580 3670
rect 4434 3632 4490 3641
rect 4528 3606 4580 3612
rect 4434 3567 4490 3576
rect 4540 3194 4568 3606
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4816 2666 4844 4134
rect 4894 3632 4950 3641
rect 4894 3567 4896 3576
rect 4948 3567 4950 3576
rect 4896 3538 4948 3544
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4816 2638 4936 2666
rect 4434 1592 4490 1601
rect 4434 1527 4490 1536
rect 3974 96 4030 105
rect 3974 31 4030 40
rect 4342 0 4398 480
rect 4448 377 4476 1527
rect 4908 480 4936 2638
rect 5092 2582 5120 2926
rect 5184 2854 5212 4950
rect 5262 4856 5318 4865
rect 5262 4791 5318 4800
rect 5276 3913 5304 4791
rect 5644 4570 5672 5238
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5828 4826 5856 5102
rect 6012 4826 6040 12242
rect 6104 10452 6132 13194
rect 6196 12986 6224 13262
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11354 6224 12242
rect 6288 11778 6316 15694
rect 6460 15642 6512 15648
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6380 15162 6408 15574
rect 6472 15162 6500 15642
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6366 14648 6422 14657
rect 6366 14583 6422 14592
rect 6380 13462 6408 14583
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 6472 13394 6500 14894
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 11898 6408 13126
rect 6472 12986 6500 13330
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6472 12374 6500 12786
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 6564 12306 6592 17190
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6932 16833 6960 17002
rect 6918 16824 6974 16833
rect 6918 16759 6920 16768
rect 6972 16759 6974 16768
rect 6920 16730 6972 16736
rect 6918 16688 6974 16697
rect 6828 16652 6880 16658
rect 6918 16623 6974 16632
rect 6828 16594 6880 16600
rect 6642 16416 6698 16425
rect 6642 16351 6698 16360
rect 6656 15638 6684 16351
rect 6734 15736 6790 15745
rect 6734 15671 6736 15680
rect 6788 15671 6790 15680
rect 6736 15642 6788 15648
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6642 15192 6698 15201
rect 6642 15127 6698 15136
rect 6656 14618 6684 15127
rect 6748 14890 6776 15438
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6748 14793 6776 14826
rect 6734 14784 6790 14793
rect 6734 14719 6790 14728
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6656 14113 6684 14418
rect 6734 14376 6790 14385
rect 6734 14311 6790 14320
rect 6642 14104 6698 14113
rect 6642 14039 6644 14048
rect 6696 14039 6698 14048
rect 6644 14010 6696 14016
rect 6644 13864 6696 13870
rect 6642 13832 6644 13841
rect 6696 13832 6698 13841
rect 6642 13767 6698 13776
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6288 11750 6408 11778
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6288 10962 6316 11494
rect 6196 10934 6316 10962
rect 6196 10520 6224 10934
rect 6274 10840 6330 10849
rect 6380 10826 6408 11750
rect 6472 11694 6500 12174
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6472 11014 6500 11630
rect 6564 11150 6592 12038
rect 6656 11801 6684 12922
rect 6642 11792 6698 11801
rect 6642 11727 6698 11736
rect 6642 11384 6698 11393
rect 6642 11319 6698 11328
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6656 11082 6684 11319
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6642 10976 6698 10985
rect 6642 10911 6698 10920
rect 6380 10798 6592 10826
rect 6274 10775 6330 10784
rect 6288 10690 6316 10775
rect 6288 10662 6408 10690
rect 6196 10492 6316 10520
rect 6104 10424 6224 10452
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6104 6458 6132 9998
rect 6196 9586 6224 10424
rect 6288 9722 6316 10492
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6380 9489 6408 10662
rect 6366 9480 6422 9489
rect 6564 9466 6592 10798
rect 6366 9415 6422 9424
rect 6472 9438 6592 9466
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5552 4542 5672 4570
rect 5460 4282 5488 4490
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5262 3904 5318 3913
rect 5262 3839 5318 3848
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5354 3088 5410 3097
rect 5354 3023 5410 3032
rect 5368 2922 5396 3023
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5460 2650 5488 3674
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5080 2576 5132 2582
rect 5552 2530 5580 4542
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4078 6040 4626
rect 6000 4072 6052 4078
rect 5998 4040 6000 4049
rect 6052 4040 6054 4049
rect 5998 3975 6054 3984
rect 6196 3924 6224 9114
rect 6288 5658 6316 9318
rect 6472 9194 6500 9438
rect 6552 9376 6604 9382
rect 6550 9344 6552 9353
rect 6604 9344 6606 9353
rect 6550 9279 6606 9288
rect 6472 9166 6592 9194
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6380 8566 6408 8774
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6380 7818 6408 8502
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6380 7546 6408 7754
rect 6472 7750 6500 8978
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6380 6118 6408 6802
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6288 5630 6408 5658
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 5030 6316 5510
rect 6380 5273 6408 5630
rect 6366 5264 6422 5273
rect 6366 5199 6422 5208
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4622 6316 4966
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6012 3896 6224 3924
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 2802 6040 3896
rect 6288 3738 6316 4558
rect 6380 4282 6408 4762
rect 6472 4593 6500 6734
rect 6564 5030 6592 9166
rect 6656 8129 6684 10911
rect 6748 8634 6776 14311
rect 6840 13818 6868 16594
rect 6932 15162 6960 16623
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6918 15056 6974 15065
rect 6918 14991 6974 15000
rect 6932 14618 6960 14991
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6840 13790 6960 13818
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13258 6868 13670
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6932 12986 6960 13790
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 11558 6868 12718
rect 6932 11558 6960 12922
rect 7024 11914 7052 17274
rect 7196 17264 7248 17270
rect 7196 17206 7248 17212
rect 7208 16658 7236 17206
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7208 15910 7236 16594
rect 7196 15904 7248 15910
rect 7102 15872 7158 15881
rect 7196 15846 7248 15852
rect 7102 15807 7158 15816
rect 7116 13734 7144 15807
rect 7208 14822 7236 15846
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 14278 7236 14309
rect 7196 14272 7248 14278
rect 7194 14240 7196 14249
rect 7248 14240 7250 14249
rect 7194 14175 7250 14184
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7116 12714 7144 13330
rect 7208 12850 7236 14175
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7300 12782 7328 18838
rect 7484 18766 7512 23990
rect 7562 23896 7618 23905
rect 7562 23831 7564 23840
rect 7616 23831 7618 23840
rect 7564 23802 7616 23808
rect 7564 23520 7616 23526
rect 7564 23462 7616 23468
rect 7576 22982 7604 23462
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7472 18624 7524 18630
rect 7378 18592 7434 18601
rect 7472 18566 7524 18572
rect 7378 18527 7434 18536
rect 7392 18154 7420 18527
rect 7484 18290 7512 18566
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7392 17066 7420 17818
rect 7484 17202 7512 18226
rect 7576 17746 7604 22918
rect 7668 20602 7696 25191
rect 7760 24274 7788 25298
rect 7840 25152 7892 25158
rect 7840 25094 7892 25100
rect 8024 25152 8076 25158
rect 8024 25094 8076 25100
rect 7748 24268 7800 24274
rect 7748 24210 7800 24216
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7760 23594 7788 24006
rect 7748 23588 7800 23594
rect 7748 23530 7800 23536
rect 7760 23050 7788 23530
rect 7748 23044 7800 23050
rect 7748 22986 7800 22992
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7760 21690 7788 22510
rect 7852 22438 7880 25094
rect 8036 24750 8064 25094
rect 8024 24744 8076 24750
rect 8024 24686 8076 24692
rect 8128 24426 8156 27520
rect 8208 25220 8260 25226
rect 8208 25162 8260 25168
rect 7944 24398 8156 24426
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7852 22234 7880 22374
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 7838 22128 7894 22137
rect 7838 22063 7894 22072
rect 7852 22030 7880 22063
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7852 21418 7880 21966
rect 7840 21412 7892 21418
rect 7840 21354 7892 21360
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7654 19272 7710 19281
rect 7654 19207 7710 19216
rect 7668 19174 7696 19207
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7760 18952 7788 21082
rect 7852 19718 7880 21354
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7668 18924 7788 18952
rect 7668 18358 7696 18924
rect 7746 18864 7802 18873
rect 7746 18799 7802 18808
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7760 17864 7788 18799
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7852 18057 7880 18566
rect 7838 18048 7894 18057
rect 7838 17983 7894 17992
rect 7760 17836 7880 17864
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7668 16130 7696 17478
rect 7484 16102 7696 16130
rect 7378 15872 7434 15881
rect 7378 15807 7434 15816
rect 7392 15473 7420 15807
rect 7378 15464 7434 15473
rect 7378 15399 7434 15408
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7288 12776 7340 12782
rect 7208 12724 7288 12730
rect 7208 12718 7340 12724
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7208 12702 7328 12718
rect 7208 12102 7236 12702
rect 7392 12594 7420 15302
rect 7484 13530 7512 16102
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7668 15366 7696 15914
rect 7656 15360 7708 15366
rect 7562 15328 7618 15337
rect 7656 15302 7708 15308
rect 7562 15263 7618 15272
rect 7576 13802 7604 15263
rect 7668 14482 7696 15302
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7668 13938 7696 14418
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7300 12566 7420 12594
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7024 11898 7236 11914
rect 7024 11892 7248 11898
rect 7024 11886 7196 11892
rect 7196 11834 7248 11840
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6840 9110 6868 11494
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10198 6960 10950
rect 7024 10577 7052 11766
rect 7116 11286 7144 11766
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7010 10568 7066 10577
rect 7010 10503 7066 10512
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 7024 9568 7052 10406
rect 7116 10305 7144 11222
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 10538 7236 11086
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7102 10296 7158 10305
rect 7208 10266 7236 10474
rect 7102 10231 7158 10240
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7024 9540 7144 9568
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6840 8809 6868 9046
rect 7024 8838 7052 9386
rect 7012 8832 7064 8838
rect 6826 8800 6882 8809
rect 7012 8774 7064 8780
rect 6826 8735 6882 8744
rect 6918 8664 6974 8673
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6840 8608 6918 8616
rect 6840 8588 6920 8608
rect 6734 8256 6790 8265
rect 6734 8191 6790 8200
rect 6642 8120 6698 8129
rect 6642 8055 6698 8064
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6656 7721 6684 7822
rect 6642 7712 6698 7721
rect 6642 7647 6698 7656
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6564 4758 6592 4966
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6458 4584 6514 4593
rect 6458 4519 6514 4528
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6366 4176 6422 4185
rect 6366 4111 6422 4120
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6380 3194 6408 4111
rect 6656 3942 6684 6666
rect 6748 5234 6776 8191
rect 6840 7954 6868 8588
rect 6972 8599 6974 8608
rect 6920 8570 6972 8576
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6920 7744 6972 7750
rect 7024 7732 7052 8774
rect 6972 7704 7052 7732
rect 6920 7686 6972 7692
rect 6826 7576 6882 7585
rect 6826 7511 6882 7520
rect 6840 6882 6868 7511
rect 6932 7342 6960 7686
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6840 6854 7052 6882
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6186 6868 6734
rect 7024 6730 7052 6854
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6918 6488 6974 6497
rect 6918 6423 6920 6432
rect 6972 6423 6974 6432
rect 6920 6394 6972 6400
rect 7024 6390 7052 6666
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 6840 5778 6868 6122
rect 7116 5914 7144 9540
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 6920 5840 6972 5846
rect 6918 5808 6920 5817
rect 6972 5808 6974 5817
rect 6828 5772 6880 5778
rect 6918 5743 6974 5752
rect 6828 5714 6880 5720
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6932 5098 6960 5646
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6932 4826 6960 5034
rect 6920 4820 6972 4826
rect 6972 4780 7144 4808
rect 6920 4762 6972 4768
rect 7010 4312 7066 4321
rect 7010 4247 7012 4256
rect 7064 4247 7066 4256
rect 7012 4218 7064 4224
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 7010 4040 7066 4049
rect 6644 3936 6696 3942
rect 6550 3904 6606 3913
rect 6644 3878 6696 3884
rect 6550 3839 6606 3848
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 5920 2774 6040 2802
rect 5920 2666 5948 2774
rect 5920 2638 6040 2666
rect 5080 2518 5132 2524
rect 5460 2502 5580 2530
rect 5460 480 5488 2502
rect 5906 2408 5962 2417
rect 5906 2343 5908 2352
rect 5960 2343 5962 2352
rect 5908 2314 5960 2320
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6012 480 6040 2638
rect 6380 2514 6408 3130
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6564 1034 6592 3839
rect 6932 3398 6960 4014
rect 7010 3975 7066 3984
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6932 3097 6960 3334
rect 7024 3194 7052 3975
rect 7116 3602 7144 4780
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7116 3194 7144 3538
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 6918 3088 6974 3097
rect 7012 3052 7064 3058
rect 6974 3032 7012 3040
rect 6918 3023 7012 3032
rect 6932 3012 7012 3023
rect 7012 2994 7064 3000
rect 7208 2938 7236 9862
rect 7300 9518 7328 12566
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7392 9897 7420 12242
rect 7378 9888 7434 9897
rect 7378 9823 7434 9832
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7392 8514 7420 9823
rect 7300 8486 7420 8514
rect 7300 5302 7328 8486
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 8022 7420 8366
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7392 7206 7420 7958
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7392 7002 7420 7142
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7484 6866 7512 13262
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7576 12850 7604 13126
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7576 11354 7604 12786
rect 7668 12714 7696 13738
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7668 12442 7696 12650
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7576 10674 7604 11290
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7576 10130 7604 10406
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9722 7604 10066
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7668 9489 7696 12038
rect 7760 9926 7788 17682
rect 7852 15502 7880 17836
rect 7944 17338 7972 24398
rect 8022 24304 8078 24313
rect 8022 24239 8024 24248
rect 8076 24239 8078 24248
rect 8024 24210 8076 24216
rect 8220 24138 8248 25162
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8208 24132 8260 24138
rect 8208 24074 8260 24080
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8024 23724 8076 23730
rect 8024 23666 8076 23672
rect 8036 23089 8064 23666
rect 8114 23352 8170 23361
rect 8114 23287 8170 23296
rect 8022 23080 8078 23089
rect 8128 23050 8156 23287
rect 8022 23015 8078 23024
rect 8116 23044 8168 23050
rect 8116 22986 8168 22992
rect 8114 22944 8170 22953
rect 8114 22879 8170 22888
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 8036 22001 8064 22578
rect 8022 21992 8078 22001
rect 8022 21927 8078 21936
rect 8024 21616 8076 21622
rect 8024 21558 8076 21564
rect 8036 21146 8064 21558
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8036 15688 8064 20198
rect 8128 18986 8156 22879
rect 8220 22681 8248 23802
rect 8312 23526 8340 24210
rect 8300 23520 8352 23526
rect 8300 23462 8352 23468
rect 8206 22672 8262 22681
rect 8206 22607 8262 22616
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8220 22098 8248 22510
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 8312 21729 8340 23462
rect 8404 23254 8432 25094
rect 8484 24676 8536 24682
rect 8484 24618 8536 24624
rect 8392 23248 8444 23254
rect 8392 23190 8444 23196
rect 8404 22778 8432 23190
rect 8496 22817 8524 24618
rect 8576 23248 8628 23254
rect 8574 23216 8576 23225
rect 8628 23216 8630 23225
rect 8574 23151 8630 23160
rect 8482 22808 8538 22817
rect 8392 22772 8444 22778
rect 8588 22778 8616 23151
rect 8482 22743 8538 22752
rect 8576 22772 8628 22778
rect 8392 22714 8444 22720
rect 8576 22714 8628 22720
rect 8680 22556 8708 27520
rect 8760 26036 8812 26042
rect 8760 25978 8812 25984
rect 8772 25498 8800 25978
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 9036 25356 9088 25362
rect 9036 25298 9088 25304
rect 8944 24880 8996 24886
rect 8944 24822 8996 24828
rect 8760 24676 8812 24682
rect 8760 24618 8812 24624
rect 8772 24177 8800 24618
rect 8852 24336 8904 24342
rect 8852 24278 8904 24284
rect 8758 24168 8814 24177
rect 8758 24103 8814 24112
rect 8864 23526 8892 24278
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 8760 23248 8812 23254
rect 8864 23225 8892 23462
rect 8760 23190 8812 23196
rect 8850 23216 8906 23225
rect 8772 22710 8800 23190
rect 8850 23151 8906 23160
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8864 22556 8892 23151
rect 8496 22528 8708 22556
rect 8772 22528 8892 22556
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8298 21720 8354 21729
rect 8298 21655 8354 21664
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 8220 20913 8248 21422
rect 8206 20904 8262 20913
rect 8206 20839 8262 20848
rect 8404 20466 8432 21830
rect 8392 20460 8444 20466
rect 8312 20420 8392 20448
rect 8312 20058 8340 20420
rect 8392 20402 8444 20408
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8312 19700 8340 19994
rect 8404 19825 8432 20198
rect 8390 19816 8446 19825
rect 8390 19751 8446 19760
rect 8312 19672 8432 19700
rect 8298 19408 8354 19417
rect 8298 19343 8354 19352
rect 8128 18958 8248 18986
rect 8116 18896 8168 18902
rect 8116 18838 8168 18844
rect 8128 18426 8156 18838
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 8220 17762 8248 18958
rect 8312 18426 8340 19343
rect 8404 19242 8432 19672
rect 8392 19236 8444 19242
rect 8392 19178 8444 19184
rect 8496 18952 8524 22528
rect 8666 22400 8722 22409
rect 8666 22335 8722 22344
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8588 21078 8616 21966
rect 8576 21072 8628 21078
rect 8576 21014 8628 21020
rect 8404 18924 8524 18952
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8220 17734 8340 17762
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8128 17066 8156 17614
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 8114 16960 8170 16969
rect 8114 16895 8170 16904
rect 7944 15660 8064 15688
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7852 15201 7880 15302
rect 7838 15192 7894 15201
rect 7944 15162 7972 15660
rect 7838 15127 7894 15136
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7852 13190 7880 14214
rect 7944 13870 7972 14758
rect 8024 14000 8076 14006
rect 8128 13988 8156 16895
rect 8220 16658 8248 17546
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 14074 8248 16594
rect 8312 16561 8340 17734
rect 8298 16552 8354 16561
rect 8298 16487 8354 16496
rect 8404 15586 8432 18924
rect 8588 18902 8616 21014
rect 8576 18896 8628 18902
rect 8482 18864 8538 18873
rect 8576 18838 8628 18844
rect 8482 18799 8538 18808
rect 8496 18766 8524 18799
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8496 17882 8524 18702
rect 8574 18048 8630 18057
rect 8574 17983 8630 17992
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8588 16046 8616 17983
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8404 15558 8616 15586
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8390 14920 8446 14929
rect 8496 14890 8524 15438
rect 8390 14855 8446 14864
rect 8484 14884 8536 14890
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8076 13960 8156 13988
rect 8024 13942 8076 13948
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7930 13424 7986 13433
rect 7930 13359 7986 13368
rect 7840 13184 7892 13190
rect 7944 13161 7972 13359
rect 8036 13326 8064 13942
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 8128 13530 8156 13670
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7840 13126 7892 13132
rect 7930 13152 7986 13161
rect 7852 12918 7880 13126
rect 7930 13087 7986 13096
rect 8128 12986 8156 13466
rect 8208 13252 8260 13258
rect 8312 13240 8340 14486
rect 8404 14414 8432 14855
rect 8484 14826 8536 14832
rect 8496 14414 8524 14826
rect 8588 14521 8616 15558
rect 8574 14512 8630 14521
rect 8574 14447 8630 14456
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8404 14006 8432 14350
rect 8496 14278 8524 14350
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 14074 8524 14214
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8260 13212 8340 13240
rect 8208 13194 8260 13200
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7852 11830 7880 12038
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7838 11656 7894 11665
rect 7838 11591 7894 11600
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7654 9480 7710 9489
rect 7564 9444 7616 9450
rect 7654 9415 7710 9424
rect 7564 9386 7616 9392
rect 7576 9042 7604 9386
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7654 8936 7710 8945
rect 7654 8871 7710 8880
rect 7562 8800 7618 8809
rect 7562 8735 7618 8744
rect 7576 8362 7604 8735
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7378 6760 7434 6769
rect 7378 6695 7380 6704
rect 7432 6695 7434 6704
rect 7380 6666 7432 6672
rect 7484 6322 7512 6802
rect 7576 6730 7604 8298
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7484 5778 7512 6122
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7668 5030 7696 8871
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4554 7696 4966
rect 7746 4584 7802 4593
rect 7656 4548 7708 4554
rect 7746 4519 7802 4528
rect 7656 4490 7708 4496
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 4078 7328 4422
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7300 2990 7328 3538
rect 6472 1006 6592 1034
rect 7024 2910 7236 2938
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 6472 480 6500 1006
rect 7024 480 7052 2910
rect 7392 2553 7420 4082
rect 7760 4010 7788 4519
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7654 3632 7710 3641
rect 7654 3567 7710 3576
rect 7668 2961 7696 3567
rect 7746 3360 7802 3369
rect 7746 3295 7802 3304
rect 7654 2952 7710 2961
rect 7760 2922 7788 3295
rect 7654 2887 7710 2896
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7378 2544 7434 2553
rect 7378 2479 7434 2488
rect 7472 2508 7524 2514
rect 7392 921 7420 2479
rect 7472 2450 7524 2456
rect 7484 2281 7512 2450
rect 7470 2272 7526 2281
rect 7470 2207 7526 2216
rect 7576 2145 7604 2790
rect 7562 2136 7618 2145
rect 7562 2071 7618 2080
rect 7852 1306 7880 11591
rect 7944 9081 7972 12582
rect 8128 12481 8156 12922
rect 8114 12472 8170 12481
rect 8114 12407 8170 12416
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8036 11121 8064 12242
rect 8220 12209 8248 12310
rect 8300 12232 8352 12238
rect 8206 12200 8262 12209
rect 8300 12174 8352 12180
rect 8206 12135 8262 12144
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8114 11792 8170 11801
rect 8114 11727 8170 11736
rect 8128 11218 8156 11727
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8022 11112 8078 11121
rect 8220 11098 8248 11834
rect 8312 11694 8340 12174
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8298 11520 8354 11529
rect 8298 11455 8354 11464
rect 8312 11150 8340 11455
rect 8022 11047 8078 11056
rect 8128 11070 8248 11098
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8128 9874 8156 11070
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8312 10248 8340 10950
rect 8220 10220 8340 10248
rect 8220 10010 8248 10220
rect 8298 10160 8354 10169
rect 8298 10095 8300 10104
rect 8352 10095 8354 10104
rect 8300 10066 8352 10072
rect 8220 9982 8340 10010
rect 8128 9846 8248 9874
rect 7930 9072 7986 9081
rect 7930 9007 7986 9016
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7944 7041 7972 8774
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7930 7032 7986 7041
rect 7930 6967 7986 6976
rect 7930 6624 7986 6633
rect 7930 6559 7986 6568
rect 7944 6458 7972 6559
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7944 6118 7972 6394
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7944 1737 7972 3878
rect 8036 3369 8064 8298
rect 8128 6458 8156 8502
rect 8220 8401 8248 9846
rect 8312 9217 8340 9982
rect 8298 9208 8354 9217
rect 8298 9143 8354 9152
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8206 8392 8262 8401
rect 8206 8327 8262 8336
rect 8312 7857 8340 8774
rect 8298 7848 8354 7857
rect 8298 7783 8354 7792
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8220 6866 8248 7278
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8128 5846 8156 6394
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8128 5166 8156 5510
rect 8220 5370 8248 6666
rect 8312 6118 8340 7686
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8312 4826 8340 6054
rect 8404 4842 8432 13942
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8588 12986 8616 13262
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8482 11928 8538 11937
rect 8482 11863 8484 11872
rect 8536 11863 8538 11872
rect 8484 11834 8536 11840
rect 8496 11286 8524 11834
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8496 9160 8524 11086
rect 8588 9586 8616 12786
rect 8680 12782 8708 22335
rect 8772 16810 8800 22528
rect 8956 22488 8984 24822
rect 9048 24614 9076 25298
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 9048 23866 9076 24550
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 9140 23662 9168 24006
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9048 23118 9076 23598
rect 9140 23254 9168 23598
rect 9128 23248 9180 23254
rect 9128 23190 9180 23196
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9128 22976 9180 22982
rect 9128 22918 9180 22924
rect 8864 22460 8984 22488
rect 8864 22098 8892 22460
rect 9048 22386 9076 22918
rect 8956 22358 9076 22386
rect 8956 22098 8984 22358
rect 9140 22250 9168 22918
rect 9232 22273 9260 27520
rect 9588 26716 9640 26722
rect 9588 26658 9640 26664
rect 9402 25392 9458 25401
rect 9402 25327 9458 25336
rect 9310 24440 9366 24449
rect 9310 24375 9366 24384
rect 9324 22982 9352 24375
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9310 22536 9366 22545
rect 9310 22471 9366 22480
rect 9048 22222 9168 22250
rect 9218 22264 9274 22273
rect 8852 22092 8904 22098
rect 8852 22034 8904 22040
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8850 21720 8906 21729
rect 8850 21655 8906 21664
rect 8864 19417 8892 21655
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8850 19408 8906 19417
rect 8850 19343 8906 19352
rect 8864 16969 8892 19343
rect 8956 18329 8984 20742
rect 8942 18320 8998 18329
rect 8942 18255 8998 18264
rect 8956 18057 8984 18255
rect 8942 18048 8998 18057
rect 8942 17983 8998 17992
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8956 17338 8984 17614
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8850 16960 8906 16969
rect 8850 16895 8906 16904
rect 8772 16782 8984 16810
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8772 15706 8800 16118
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8864 14793 8892 16662
rect 8850 14784 8906 14793
rect 8850 14719 8906 14728
rect 8864 14618 8892 14719
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8864 13870 8892 14554
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8864 13682 8892 13806
rect 8772 13654 8892 13682
rect 8772 13462 8800 13654
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8680 12442 8708 12718
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8772 12209 8800 12854
rect 8864 12646 8892 13466
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8864 12442 8892 12582
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8758 12200 8814 12209
rect 8668 12164 8720 12170
rect 8758 12135 8814 12144
rect 8668 12106 8720 12112
rect 8680 9625 8708 12106
rect 8956 11778 8984 16782
rect 9048 13530 9076 22222
rect 9218 22199 9274 22208
rect 9128 22160 9180 22166
rect 9128 22102 9180 22108
rect 9140 17218 9168 22102
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 9232 20641 9260 21830
rect 9218 20632 9274 20641
rect 9324 20602 9352 22471
rect 9416 22166 9444 25327
rect 9600 24993 9628 26658
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 9586 24984 9642 24993
rect 9508 24942 9586 24970
rect 9508 24585 9536 24942
rect 9586 24919 9642 24928
rect 9692 24698 9720 25094
rect 9784 24857 9812 27520
rect 10138 26480 10194 26489
rect 10138 26415 10194 26424
rect 9954 26344 10010 26353
rect 9954 26279 10010 26288
rect 9864 26172 9916 26178
rect 9864 26114 9916 26120
rect 9876 25140 9904 26114
rect 9968 25702 9996 26279
rect 10048 26172 10100 26178
rect 10048 26114 10100 26120
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 10060 25498 10088 26114
rect 10152 25537 10180 26415
rect 10336 25786 10364 27520
rect 10784 26852 10836 26858
rect 10784 26794 10836 26800
rect 10336 25758 10732 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10138 25528 10194 25537
rect 10048 25492 10100 25498
rect 10289 25520 10585 25540
rect 10138 25463 10194 25472
rect 10048 25434 10100 25440
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9876 25112 9996 25140
rect 9770 24848 9826 24857
rect 9770 24783 9826 24792
rect 9692 24670 9812 24698
rect 9588 24608 9640 24614
rect 9494 24576 9550 24585
rect 9588 24550 9640 24556
rect 9494 24511 9550 24520
rect 9600 24313 9628 24550
rect 9586 24304 9642 24313
rect 9586 24239 9642 24248
rect 9496 24064 9548 24070
rect 9496 24006 9548 24012
rect 9404 22160 9456 22166
rect 9404 22102 9456 22108
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9416 21593 9444 21966
rect 9508 21865 9536 24006
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9494 21856 9550 21865
rect 9494 21791 9550 21800
rect 9402 21584 9458 21593
rect 9402 21519 9458 21528
rect 9600 21434 9628 22918
rect 9416 21406 9628 21434
rect 9416 20777 9444 21406
rect 9496 21344 9548 21350
rect 9496 21286 9548 21292
rect 9402 20768 9458 20777
rect 9402 20703 9458 20712
rect 9218 20567 9274 20576
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9508 20505 9536 21286
rect 9692 21078 9720 23462
rect 9784 22506 9812 24670
rect 9864 24676 9916 24682
rect 9864 24618 9916 24624
rect 9876 24070 9904 24618
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9876 23361 9904 24006
rect 9862 23352 9918 23361
rect 9862 23287 9918 23296
rect 9968 22658 9996 25112
rect 10060 24614 10088 25230
rect 10140 24676 10192 24682
rect 10140 24618 10192 24624
rect 10048 24608 10100 24614
rect 10048 24550 10100 24556
rect 10060 22778 10088 24550
rect 10152 23662 10180 24618
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10612 23662 10640 24142
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 9968 22630 10180 22658
rect 9772 22500 9824 22506
rect 9772 22442 9824 22448
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9784 21146 9812 22034
rect 9862 21992 9918 22001
rect 9862 21927 9864 21936
rect 9916 21927 9918 21936
rect 9864 21898 9916 21904
rect 10046 21856 10102 21865
rect 10046 21791 10102 21800
rect 10060 21434 10088 21791
rect 9864 21412 9916 21418
rect 9864 21354 9916 21360
rect 9968 21406 10088 21434
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9680 21072 9732 21078
rect 9600 21020 9680 21026
rect 9600 21014 9732 21020
rect 9600 20998 9720 21014
rect 9494 20496 9550 20505
rect 9494 20431 9550 20440
rect 9600 20058 9628 20998
rect 9680 20936 9732 20942
rect 9678 20904 9680 20913
rect 9732 20904 9734 20913
rect 9678 20839 9734 20848
rect 9692 20534 9720 20839
rect 9770 20768 9826 20777
rect 9770 20703 9826 20712
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9784 20330 9812 20703
rect 9772 20324 9824 20330
rect 9772 20266 9824 20272
rect 9680 20256 9732 20262
rect 9678 20224 9680 20233
rect 9732 20224 9734 20233
rect 9678 20159 9734 20168
rect 9770 20088 9826 20097
rect 9588 20052 9640 20058
rect 9770 20023 9826 20032
rect 9588 19994 9640 20000
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9508 19009 9536 19382
rect 9494 19000 9550 19009
rect 9692 18986 9720 19926
rect 9784 19825 9812 20023
rect 9876 19854 9904 21354
rect 9968 20466 9996 21406
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9954 20088 10010 20097
rect 9954 20023 10010 20032
rect 9864 19848 9916 19854
rect 9770 19816 9826 19825
rect 9864 19790 9916 19796
rect 9770 19751 9826 19760
rect 9772 19712 9824 19718
rect 9968 19700 9996 20023
rect 9772 19654 9824 19660
rect 9876 19672 9996 19700
rect 9784 19145 9812 19654
rect 9770 19136 9826 19145
rect 9770 19071 9826 19080
rect 9600 18970 9720 18986
rect 9494 18935 9550 18944
rect 9588 18964 9720 18970
rect 9640 18958 9720 18964
rect 9588 18906 9640 18912
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9508 18086 9536 18702
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9140 17190 9260 17218
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9140 16250 9168 17002
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9034 13016 9090 13025
rect 9034 12951 9090 12960
rect 9048 12918 9076 12951
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 9140 12850 9168 15982
rect 9232 12986 9260 17190
rect 9324 16425 9352 18022
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9310 16416 9366 16425
rect 9310 16351 9366 16360
rect 9416 15745 9444 17682
rect 9402 15736 9458 15745
rect 9402 15671 9458 15680
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14482 9352 14758
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9128 12708 9180 12714
rect 9048 12668 9128 12696
rect 9048 12345 9076 12668
rect 9128 12650 9180 12656
rect 9232 12356 9260 12922
rect 9324 12782 9352 13126
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9034 12336 9090 12345
rect 9034 12271 9036 12280
rect 9088 12271 9090 12280
rect 9140 12328 9260 12356
rect 9036 12242 9088 12248
rect 9048 12211 9076 12242
rect 9140 12050 9168 12328
rect 8772 11750 8984 11778
rect 9048 12022 9168 12050
rect 8772 11218 8800 11750
rect 8942 11656 8998 11665
rect 8942 11591 8944 11600
rect 8996 11591 8998 11600
rect 8944 11562 8996 11568
rect 8850 11520 8906 11529
rect 8850 11455 8906 11464
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8666 9616 8722 9625
rect 8576 9580 8628 9586
rect 8666 9551 8722 9560
rect 8576 9522 8628 9528
rect 8496 9132 8616 9160
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8362 8524 8978
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8496 8265 8524 8298
rect 8482 8256 8538 8265
rect 8482 8191 8538 8200
rect 8482 8120 8538 8129
rect 8482 8055 8538 8064
rect 8496 7546 8524 8055
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8588 7002 8616 9132
rect 8680 8498 8708 9551
rect 8772 8945 8800 11018
rect 8758 8936 8814 8945
rect 8758 8871 8814 8880
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8680 7177 8708 7686
rect 8666 7168 8722 7177
rect 8666 7103 8722 7112
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8496 5914 8524 6734
rect 8588 6225 8616 6938
rect 8772 6905 8800 8774
rect 8758 6896 8814 6905
rect 8758 6831 8814 6840
rect 8666 6760 8722 6769
rect 8666 6695 8722 6704
rect 8574 6216 8630 6225
rect 8574 6151 8630 6160
rect 8680 5953 8708 6695
rect 8666 5944 8722 5953
rect 8484 5908 8536 5914
rect 8666 5879 8722 5888
rect 8484 5850 8536 5856
rect 8758 5128 8814 5137
rect 8758 5063 8760 5072
rect 8812 5063 8814 5072
rect 8760 5034 8812 5040
rect 8300 4820 8352 4826
rect 8404 4814 8616 4842
rect 8864 4826 8892 11455
rect 8956 9654 8984 11562
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 6769 8984 8910
rect 8942 6760 8998 6769
rect 8942 6695 8998 6704
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 5098 8984 6598
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 8300 4762 8352 4768
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 4146 8340 4626
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 8484 4004 8536 4010
rect 8022 3360 8078 3369
rect 8022 3295 8078 3304
rect 7930 1728 7986 1737
rect 7930 1663 7986 1672
rect 7576 1278 7880 1306
rect 7378 912 7434 921
rect 7378 847 7434 856
rect 7576 480 7604 1278
rect 8128 480 8156 3975
rect 8484 3946 8536 3952
rect 8496 3194 8524 3946
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8220 2310 8248 2926
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8588 480 8616 4814
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8758 4720 8814 4729
rect 8758 4655 8814 4664
rect 8772 4214 8800 4655
rect 8864 4282 8892 4762
rect 8956 4554 8984 5034
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 9048 4049 9076 12022
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9034 4040 9090 4049
rect 9034 3975 9090 3984
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8956 1873 8984 2246
rect 8942 1864 8998 1873
rect 8942 1799 8998 1808
rect 9140 480 9168 11834
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9232 10810 9260 11630
rect 9324 11014 9352 12718
rect 9416 12696 9444 15671
rect 9508 15065 9536 18022
rect 9600 17678 9628 18022
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9692 17610 9720 18958
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9588 17536 9640 17542
rect 9640 17484 9720 17490
rect 9588 17478 9720 17484
rect 9600 17462 9720 17478
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9600 15745 9628 15846
rect 9586 15736 9642 15745
rect 9586 15671 9642 15680
rect 9494 15056 9550 15065
rect 9494 14991 9550 15000
rect 9600 14958 9628 15671
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9692 14278 9720 17462
rect 9784 16114 9812 18702
rect 9876 17746 9904 19672
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9968 18630 9996 19246
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 18154 9996 18566
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9862 17640 9918 17649
rect 9862 17575 9918 17584
rect 9876 16794 9904 17575
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9876 16153 9904 16526
rect 9862 16144 9918 16153
rect 9772 16108 9824 16114
rect 9862 16079 9918 16088
rect 9772 16050 9824 16056
rect 9770 16008 9826 16017
rect 9770 15943 9826 15952
rect 9784 15706 9812 15943
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9770 15192 9826 15201
rect 9770 15127 9826 15136
rect 9784 14618 9812 15127
rect 9876 14958 9904 16079
rect 9968 15609 9996 17070
rect 9954 15600 10010 15609
rect 9954 15535 10010 15544
rect 9954 15464 10010 15473
rect 9954 15399 10010 15408
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9862 14376 9918 14385
rect 9862 14311 9918 14320
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9494 14104 9550 14113
rect 9494 14039 9550 14048
rect 9508 12866 9536 14039
rect 9678 13968 9734 13977
rect 9678 13903 9734 13912
rect 9692 13818 9720 13903
rect 9600 13790 9720 13818
rect 9770 13832 9826 13841
rect 9600 13734 9628 13790
rect 9770 13767 9826 13776
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9678 13696 9734 13705
rect 9678 13631 9734 13640
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9600 12986 9628 13398
rect 9692 13394 9720 13631
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9678 13016 9734 13025
rect 9588 12980 9640 12986
rect 9678 12951 9734 12960
rect 9588 12922 9640 12928
rect 9692 12866 9720 12951
rect 9508 12838 9720 12866
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9416 12668 9536 12696
rect 9508 12306 9536 12668
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9324 10266 9352 10950
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9232 9897 9260 9930
rect 9218 9888 9274 9897
rect 9218 9823 9274 9832
rect 9324 9586 9352 10202
rect 9402 10024 9458 10033
rect 9402 9959 9458 9968
rect 9508 9976 9536 12038
rect 9600 11898 9628 12718
rect 9692 12481 9720 12838
rect 9678 12472 9734 12481
rect 9678 12407 9734 12416
rect 9680 12368 9732 12374
rect 9678 12336 9680 12345
rect 9732 12336 9734 12345
rect 9678 12271 9734 12280
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9600 11608 9628 11698
rect 9784 11608 9812 13767
rect 9876 12714 9904 14311
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9968 12594 9996 15399
rect 10060 14770 10088 21286
rect 10152 18766 10180 22630
rect 10244 22574 10272 23122
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10336 22506 10364 22918
rect 10324 22500 10376 22506
rect 10324 22442 10376 22448
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10232 22160 10284 22166
rect 10232 22102 10284 22108
rect 10244 21486 10272 22102
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10232 21480 10284 21486
rect 10232 21422 10284 21428
rect 10520 21418 10548 21966
rect 10704 21593 10732 25758
rect 10796 25430 10824 26794
rect 10784 25424 10836 25430
rect 10784 25366 10836 25372
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 10796 23905 10824 25230
rect 10782 23896 10838 23905
rect 10782 23831 10838 23840
rect 10796 22642 10824 23831
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10888 22386 10916 27520
rect 11440 26602 11468 27520
rect 11440 26574 11928 26602
rect 11704 26512 11756 26518
rect 11704 26454 11756 26460
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11150 25800 11206 25809
rect 11150 25735 11206 25744
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 10980 24614 11008 25298
rect 11072 24886 11100 25434
rect 11164 25265 11192 25735
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 11336 25356 11388 25362
rect 11336 25298 11388 25304
rect 11150 25256 11206 25265
rect 11150 25191 11206 25200
rect 11060 24880 11112 24886
rect 11060 24822 11112 24828
rect 11348 24818 11376 25298
rect 11440 24954 11468 25638
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10796 22358 10916 22386
rect 10796 21978 10824 22358
rect 10980 22250 11008 24550
rect 11244 24404 11296 24410
rect 11244 24346 11296 24352
rect 11058 24168 11114 24177
rect 11058 24103 11114 24112
rect 10888 22222 11008 22250
rect 11072 22234 11100 24103
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 11164 23186 11192 23462
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 11256 22642 11284 24346
rect 11428 24268 11480 24274
rect 11428 24210 11480 24216
rect 11440 23798 11468 24210
rect 11428 23792 11480 23798
rect 11428 23734 11480 23740
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11336 22976 11388 22982
rect 11336 22918 11388 22924
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11242 22264 11298 22273
rect 11060 22228 11112 22234
rect 10888 22098 10916 22222
rect 11242 22199 11298 22208
rect 11060 22170 11112 22176
rect 10966 22128 11022 22137
rect 10876 22092 10928 22098
rect 10966 22063 11022 22072
rect 10876 22034 10928 22040
rect 10796 21950 10916 21978
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10690 21584 10746 21593
rect 10690 21519 10746 21528
rect 10508 21412 10560 21418
rect 10508 21354 10560 21360
rect 10796 21350 10824 21830
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10796 20466 10824 21286
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10888 20346 10916 21950
rect 10980 21690 11008 22063
rect 11150 21992 11206 22001
rect 11150 21927 11206 21936
rect 11060 21888 11112 21894
rect 11058 21856 11060 21865
rect 11112 21856 11114 21865
rect 11058 21791 11114 21800
rect 11058 21720 11114 21729
rect 10968 21684 11020 21690
rect 11058 21655 11114 21664
rect 10968 21626 11020 21632
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10980 20602 11008 21490
rect 11072 21146 11100 21655
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 10704 20318 10916 20346
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10612 19514 10640 19858
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10152 17746 10180 18566
rect 10244 18426 10272 18702
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10704 18306 10732 20318
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10796 19174 10824 19790
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10888 19553 10916 19722
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10874 19544 10930 19553
rect 10874 19479 10930 19488
rect 10980 19292 11008 19654
rect 11072 19446 11100 20742
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 10980 19264 11100 19292
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10612 18278 10732 18306
rect 10612 18222 10640 18278
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10324 17808 10376 17814
rect 10322 17776 10324 17785
rect 10376 17776 10378 17785
rect 10140 17740 10192 17746
rect 10322 17711 10378 17720
rect 10140 17682 10192 17688
rect 10152 15162 10180 17682
rect 10704 17678 10732 18090
rect 10796 18086 10824 19110
rect 10888 18902 10916 19178
rect 11072 19174 11100 19264
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10888 18358 10916 18838
rect 11072 18426 11100 19110
rect 11164 18465 11192 21927
rect 11256 20806 11284 22199
rect 11348 21962 11376 22918
rect 11440 22642 11468 23190
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 11440 22166 11468 22578
rect 11428 22160 11480 22166
rect 11428 22102 11480 22108
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11348 21418 11376 21898
rect 11428 21616 11480 21622
rect 11428 21558 11480 21564
rect 11336 21412 11388 21418
rect 11336 21354 11388 21360
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11242 20632 11298 20641
rect 11242 20567 11298 20576
rect 11256 20330 11284 20567
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 11256 19281 11284 20266
rect 11348 20233 11376 20402
rect 11334 20224 11390 20233
rect 11334 20159 11390 20168
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 11242 19272 11298 19281
rect 11242 19207 11298 19216
rect 11348 19174 11376 19926
rect 11244 19168 11296 19174
rect 11336 19168 11388 19174
rect 11244 19110 11296 19116
rect 11334 19136 11336 19145
rect 11388 19136 11390 19145
rect 11150 18456 11206 18465
rect 11060 18420 11112 18426
rect 11150 18391 11206 18400
rect 11060 18362 11112 18368
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16794 10732 17614
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10322 16688 10378 16697
rect 10232 16652 10284 16658
rect 10322 16623 10378 16632
rect 10232 16594 10284 16600
rect 10244 15978 10272 16594
rect 10336 16046 10364 16623
rect 10796 16590 10824 17478
rect 10888 16697 10916 18158
rect 11072 17610 11100 18226
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 10968 17536 11020 17542
rect 11020 17484 11100 17490
rect 10968 17478 11100 17484
rect 10980 17462 11100 17478
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10980 16726 11008 17206
rect 11072 16998 11100 17462
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16794 11100 16934
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10968 16720 11020 16726
rect 10874 16688 10930 16697
rect 10968 16662 11020 16668
rect 10874 16623 10930 16632
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 16114 10916 16390
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15706 10732 15982
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10888 15745 10916 15846
rect 10874 15736 10930 15745
rect 10692 15700 10744 15706
rect 10744 15660 10824 15688
rect 10980 15706 11008 16662
rect 10874 15671 10930 15680
rect 10968 15700 11020 15706
rect 10692 15642 10744 15648
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10060 14742 10180 14770
rect 10046 14648 10102 14657
rect 10046 14583 10102 14592
rect 10060 14550 10088 14583
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 10046 14104 10102 14113
rect 10046 14039 10048 14048
rect 10100 14039 10102 14048
rect 10048 14010 10100 14016
rect 10046 13560 10102 13569
rect 10046 13495 10048 13504
rect 10100 13495 10102 13504
rect 10048 13466 10100 13472
rect 9968 12566 10088 12594
rect 9862 12472 9918 12481
rect 9862 12407 9918 12416
rect 9600 11580 9812 11608
rect 9692 9994 9720 11580
rect 9770 11384 9826 11393
rect 9770 11319 9826 11328
rect 9784 10554 9812 11319
rect 9876 10810 9904 12407
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9784 10526 9904 10554
rect 9770 10432 9826 10441
rect 9770 10367 9826 10376
rect 9680 9988 9732 9994
rect 9416 9926 9444 9959
rect 9508 9948 9628 9976
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9494 9888 9550 9897
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9324 9178 9352 9522
rect 9416 9382 9444 9862
rect 9494 9823 9550 9832
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9232 8090 9260 8298
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9218 7440 9274 7449
rect 9218 7375 9220 7384
rect 9272 7375 9274 7384
rect 9220 7346 9272 7352
rect 9324 5710 9352 8842
rect 9416 8362 9444 9318
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9416 6458 9444 8026
rect 9508 6798 9536 9823
rect 9600 7585 9628 9948
rect 9680 9930 9732 9936
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 8906 9720 9522
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9586 7576 9642 7585
rect 9586 7511 9642 7520
rect 9692 7426 9720 8298
rect 9784 7449 9812 10367
rect 9876 9081 9904 10526
rect 9968 9466 9996 12242
rect 10060 9586 10088 12566
rect 10152 11898 10180 14742
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 14074 10548 14350
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 10336 12782 10364 13398
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10520 12714 10548 13126
rect 10612 12782 10640 13330
rect 10704 13297 10732 15506
rect 10796 15162 10824 15660
rect 10968 15642 11020 15648
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10796 15008 10824 15098
rect 11072 15026 11100 16730
rect 11164 15570 11192 18022
rect 11256 17082 11284 19110
rect 11334 19071 11390 19080
rect 11348 18193 11376 19071
rect 11440 18290 11468 21558
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11334 18184 11390 18193
rect 11334 18119 11390 18128
rect 11334 17368 11390 17377
rect 11334 17303 11390 17312
rect 11348 17202 11376 17303
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11256 17054 11376 17082
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11060 15020 11112 15026
rect 10796 14980 10916 15008
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10690 13288 10746 13297
rect 10690 13223 10746 13232
rect 10796 13172 10824 14826
rect 10704 13144 10824 13172
rect 10600 12776 10652 12782
rect 10598 12744 10600 12753
rect 10652 12744 10654 12753
rect 10508 12708 10560 12714
rect 10598 12679 10654 12688
rect 10508 12650 10560 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12424 10732 13144
rect 10888 13002 10916 14980
rect 11060 14962 11112 14968
rect 11058 14784 11114 14793
rect 11058 14719 11114 14728
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10980 13138 11008 14214
rect 11072 13977 11100 14719
rect 11164 14618 11192 15506
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11058 13968 11114 13977
rect 11058 13903 11114 13912
rect 11164 13734 11192 14418
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11058 13560 11114 13569
rect 11058 13495 11114 13504
rect 11072 13462 11100 13495
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 10980 13110 11100 13138
rect 10888 12974 11008 13002
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10612 12396 10732 12424
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11898 10548 12174
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10152 11286 10180 11698
rect 10612 11676 10640 12396
rect 10784 12300 10836 12306
rect 10888 12288 10916 12854
rect 10836 12260 10916 12288
rect 10784 12242 10836 12248
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11830 10732 12038
rect 10692 11824 10744 11830
rect 10690 11792 10692 11801
rect 10744 11792 10746 11801
rect 10690 11727 10746 11736
rect 10888 11694 10916 12260
rect 10876 11688 10928 11694
rect 10612 11648 10732 11676
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10322 11112 10378 11121
rect 10322 11047 10378 11056
rect 10336 10742 10364 11047
rect 10704 10826 10732 11648
rect 10876 11630 10928 11636
rect 10876 11552 10928 11558
rect 10782 11520 10838 11529
rect 10876 11494 10928 11500
rect 10782 11455 10838 11464
rect 10796 10962 10824 11455
rect 10888 11064 10916 11494
rect 10980 11286 11008 12974
rect 11072 11626 11100 13110
rect 11164 12458 11192 13670
rect 11256 13462 11284 16934
rect 11348 14278 11376 17054
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11440 15910 11468 16390
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11440 15366 11468 15846
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11440 14822 11468 15302
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11440 13530 11468 14554
rect 11532 13802 11560 26318
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 11624 19854 11652 24550
rect 11716 22273 11744 26454
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 11808 24886 11836 25298
rect 11796 24880 11848 24886
rect 11796 24822 11848 24828
rect 11794 24168 11850 24177
rect 11794 24103 11850 24112
rect 11808 23633 11836 24103
rect 11900 24041 11928 26574
rect 11992 24274 12020 27520
rect 12440 26648 12492 26654
rect 12440 26590 12492 26596
rect 12254 24712 12310 24721
rect 12254 24647 12310 24656
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 11980 24064 12032 24070
rect 11886 24032 11942 24041
rect 11980 24006 12032 24012
rect 11886 23967 11942 23976
rect 11794 23624 11850 23633
rect 11900 23610 11928 23967
rect 11992 23730 12020 24006
rect 11980 23724 12032 23730
rect 11980 23666 12032 23672
rect 11978 23624 12034 23633
rect 11900 23582 11978 23610
rect 11794 23559 11850 23568
rect 11978 23559 12034 23568
rect 11808 22778 11836 23559
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11702 22264 11758 22273
rect 11702 22199 11758 22208
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 11716 20942 11744 22034
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 11704 20936 11756 20942
rect 11702 20904 11704 20913
rect 11756 20904 11758 20913
rect 11702 20839 11758 20848
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11624 19174 11652 19790
rect 11704 19780 11756 19786
rect 11808 19768 11836 21966
rect 11900 20233 11928 22374
rect 11992 21554 12020 22918
rect 12176 22574 12204 23122
rect 12268 23050 12296 24647
rect 12452 24206 12480 26590
rect 12544 25362 12572 27520
rect 13096 25498 13124 27520
rect 13176 26444 13228 26450
rect 13176 26386 13228 26392
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12532 25152 12584 25158
rect 12716 25152 12768 25158
rect 12584 25112 12664 25140
rect 12532 25094 12584 25100
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12544 24410 12572 24550
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12530 24168 12586 24177
rect 12530 24103 12586 24112
rect 12544 23866 12572 24103
rect 12348 23860 12400 23866
rect 12532 23860 12584 23866
rect 12400 23820 12480 23848
rect 12348 23802 12400 23808
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 12360 23338 12388 23530
rect 12452 23508 12480 23820
rect 12532 23802 12584 23808
rect 12636 23662 12664 25112
rect 12716 25094 12768 25100
rect 12728 24410 12756 25094
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12728 23594 12756 24346
rect 12820 24138 12848 25230
rect 12992 25220 13044 25226
rect 12992 25162 13044 25168
rect 13004 24682 13032 25162
rect 13082 24848 13138 24857
rect 13082 24783 13084 24792
rect 13136 24783 13138 24792
rect 13084 24754 13136 24760
rect 12992 24676 13044 24682
rect 12992 24618 13044 24624
rect 13084 24676 13136 24682
rect 13084 24618 13136 24624
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12820 23798 12848 24074
rect 12808 23792 12860 23798
rect 12808 23734 12860 23740
rect 12716 23588 12768 23594
rect 12716 23530 12768 23536
rect 12452 23480 12572 23508
rect 12360 23322 12480 23338
rect 12360 23316 12492 23322
rect 12360 23310 12440 23316
rect 12256 23044 12308 23050
rect 12256 22986 12308 22992
rect 12164 22568 12216 22574
rect 12162 22536 12164 22545
rect 12216 22536 12218 22545
rect 12162 22471 12218 22480
rect 12072 22160 12124 22166
rect 12360 22137 12388 23310
rect 12440 23258 12492 23264
rect 12544 22545 12572 23480
rect 12806 23488 12862 23497
rect 12806 23423 12862 23432
rect 12530 22536 12586 22545
rect 12530 22471 12586 22480
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12072 22102 12124 22108
rect 12346 22128 12402 22137
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11980 21344 12032 21350
rect 12084 21332 12112 22102
rect 12346 22063 12402 22072
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12032 21304 12112 21332
rect 11980 21286 12032 21292
rect 11886 20224 11942 20233
rect 11886 20159 11942 20168
rect 11808 19740 11928 19768
rect 11704 19722 11756 19728
rect 11716 19666 11744 19722
rect 11716 19638 11836 19666
rect 11808 19446 11836 19638
rect 11704 19440 11756 19446
rect 11704 19382 11756 19388
rect 11796 19440 11848 19446
rect 11796 19382 11848 19388
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 11624 18329 11652 19110
rect 11610 18320 11666 18329
rect 11610 18255 11666 18264
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11624 13682 11652 18255
rect 11716 17354 11744 19382
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11808 18970 11836 19246
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11808 18086 11836 18770
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11808 17746 11836 18022
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11716 17326 11836 17354
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 14618 11744 15846
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11702 13968 11758 13977
rect 11702 13903 11758 13912
rect 11532 13654 11652 13682
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11256 12850 11284 13194
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11440 12782 11468 13126
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11244 12640 11296 12646
rect 11242 12608 11244 12617
rect 11296 12608 11298 12617
rect 11242 12543 11298 12552
rect 11164 12430 11284 12458
rect 11060 11620 11112 11626
rect 11112 11580 11192 11608
rect 11060 11562 11112 11568
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10888 11036 11008 11064
rect 10796 10934 10916 10962
rect 10704 10798 10824 10826
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10138 10296 10194 10305
rect 10289 10288 10585 10308
rect 10138 10231 10194 10240
rect 10152 10198 10180 10231
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10140 9512 10192 9518
rect 9968 9438 10088 9466
rect 10140 9454 10192 9460
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9862 9072 9918 9081
rect 9862 9007 9918 9016
rect 9876 8090 9904 9007
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7478 9904 7822
rect 9864 7472 9916 7478
rect 9600 7398 9720 7426
rect 9770 7440 9826 7449
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 4078 9352 5510
rect 9416 5234 9444 6394
rect 9508 5914 9536 6598
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9416 4826 9444 5170
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9416 4146 9444 4762
rect 9600 4457 9628 7398
rect 9864 7414 9916 7420
rect 9770 7375 9826 7384
rect 9784 7342 9812 7375
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6798 9720 7142
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9692 5642 9720 6734
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 6225 9812 6598
rect 9770 6216 9826 6225
rect 9770 6151 9826 6160
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9678 5536 9734 5545
rect 9678 5471 9734 5480
rect 9692 4622 9720 5471
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9784 4554 9812 5782
rect 9862 4856 9918 4865
rect 9862 4791 9918 4800
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9586 4448 9642 4457
rect 9586 4383 9642 4392
rect 9494 4312 9550 4321
rect 9494 4247 9550 4256
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9508 4010 9536 4247
rect 9876 4146 9904 4791
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9968 4026 9996 9318
rect 10060 8498 10088 9438
rect 10152 9353 10180 9454
rect 10244 9450 10272 9998
rect 10428 9926 10456 9998
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10520 9518 10548 10066
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10600 9920 10652 9926
rect 10704 9897 10732 9998
rect 10600 9862 10652 9868
rect 10690 9888 10746 9897
rect 10612 9722 10640 9862
rect 10690 9823 10746 9832
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10138 9344 10194 9353
rect 10138 9279 10194 9288
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10060 7274 10088 8026
rect 10152 8022 10180 8230
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10152 7546 10180 7958
rect 10414 7576 10470 7585
rect 10140 7540 10192 7546
rect 10414 7511 10470 7520
rect 10140 7482 10192 7488
rect 10428 7342 10456 7511
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10704 6984 10732 9386
rect 10796 7857 10824 10798
rect 10888 9738 10916 10934
rect 10980 10810 11008 11036
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10980 10266 11008 10474
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11072 9994 11100 11290
rect 11164 9994 11192 11580
rect 11256 10282 11284 12430
rect 11440 12306 11468 12718
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11348 11218 11376 11834
rect 11440 11626 11468 12242
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11348 10742 11376 11154
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11336 10464 11388 10470
rect 11334 10432 11336 10441
rect 11388 10432 11390 10441
rect 11334 10367 11390 10376
rect 11256 10254 11376 10282
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 10888 9710 11008 9738
rect 10876 9648 10928 9654
rect 10874 9616 10876 9625
rect 10928 9616 10930 9625
rect 10874 9551 10930 9560
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10888 8430 10916 9046
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10782 7848 10838 7857
rect 10782 7783 10838 7792
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10612 6956 10732 6984
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 5370 10088 6802
rect 10612 6322 10640 6956
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5846 10732 6598
rect 10796 5846 10824 7482
rect 10888 7478 10916 8230
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10888 6458 10916 6734
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10796 5166 10824 5782
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10048 4752 10100 4758
rect 10046 4720 10048 4729
rect 10100 4720 10102 4729
rect 10046 4655 10102 4664
rect 10152 4282 10180 4966
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10782 4856 10838 4865
rect 10782 4791 10838 4800
rect 10796 4758 10824 4791
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10244 4622 10272 4694
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10244 4214 10272 4558
rect 10796 4214 10824 4694
rect 10888 4690 10916 6258
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10980 4146 11008 9710
rect 11072 9602 11100 9930
rect 11072 9574 11192 9602
rect 11058 9480 11114 9489
rect 11058 9415 11114 9424
rect 11072 8974 11100 9415
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8634 11100 8910
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11164 8299 11192 9574
rect 11348 9110 11376 10254
rect 11440 10044 11468 10746
rect 11532 10146 11560 13654
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12850 11652 13262
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11624 10810 11652 11698
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11532 10118 11652 10146
rect 11440 10016 11560 10044
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11440 9761 11468 9862
rect 11426 9752 11482 9761
rect 11426 9687 11482 9696
rect 11440 9586 11468 9687
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11150 8290 11206 8299
rect 11150 8225 11206 8234
rect 11058 7984 11114 7993
rect 11058 7919 11114 7928
rect 11072 7546 11100 7919
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11058 6624 11114 6633
rect 11058 6559 11114 6568
rect 11072 6322 11100 6559
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 5030 11100 5510
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9876 3998 9996 4026
rect 10048 4004 10100 4010
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 3505 9812 3538
rect 9494 3496 9550 3505
rect 9770 3496 9826 3505
rect 9494 3431 9496 3440
rect 9548 3431 9550 3440
rect 9600 3454 9770 3482
rect 9496 3402 9548 3408
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9232 2650 9260 2994
rect 9324 2990 9352 3334
rect 9600 3194 9628 3454
rect 9770 3431 9826 3440
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9496 2984 9548 2990
rect 9548 2932 9720 2938
rect 9496 2926 9720 2932
rect 9508 2922 9720 2926
rect 9508 2916 9732 2922
rect 9508 2910 9680 2916
rect 9680 2858 9732 2864
rect 9876 2666 9904 3998
rect 10048 3946 10100 3952
rect 10060 3777 10088 3946
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10046 3768 10102 3777
rect 10289 3760 10585 3780
rect 10980 3738 11008 4082
rect 10046 3703 10102 3712
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10782 3360 10838 3369
rect 10782 3295 10838 3304
rect 10138 2952 10194 2961
rect 10138 2887 10194 2896
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9692 2638 9904 2666
rect 9692 480 9720 2638
rect 10152 480 10180 2887
rect 10692 2848 10744 2854
rect 10796 2825 10824 3295
rect 10876 2848 10928 2854
rect 10692 2790 10744 2796
rect 10782 2816 10838 2825
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2689 10732 2790
rect 10876 2790 10928 2796
rect 10782 2751 10838 2760
rect 10690 2680 10746 2689
rect 10888 2650 10916 2790
rect 10690 2615 10746 2624
rect 10876 2644 10928 2650
rect 10322 2544 10378 2553
rect 10322 2479 10324 2488
rect 10376 2479 10378 2488
rect 10324 2450 10376 2456
rect 10704 2394 10732 2615
rect 10876 2586 10928 2592
rect 10980 2530 11008 3470
rect 11072 2854 11100 3470
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10980 2514 11100 2530
rect 10980 2508 11112 2514
rect 10980 2502 11060 2508
rect 11060 2450 11112 2456
rect 10520 2366 10732 2394
rect 10520 2281 10548 2366
rect 10506 2272 10562 2281
rect 10506 2207 10562 2216
rect 10690 2272 10746 2281
rect 10690 2207 10746 2216
rect 10704 480 10732 2207
rect 11164 2009 11192 7686
rect 11256 6934 11284 7754
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 6458 11284 6734
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11348 6361 11376 8774
rect 11532 7154 11560 10016
rect 11624 9382 11652 10118
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11624 7546 11652 9114
rect 11716 7750 11744 13903
rect 11808 13410 11836 17326
rect 11900 16697 11928 19740
rect 11992 19553 12020 21286
rect 12268 21146 12296 21966
rect 12348 21480 12400 21486
rect 12452 21468 12480 22374
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12728 21690 12756 21830
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12728 21486 12756 21626
rect 12400 21440 12480 21468
rect 12716 21480 12768 21486
rect 12348 21422 12400 21428
rect 12716 21422 12768 21428
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12268 20874 12296 21082
rect 12256 20868 12308 20874
rect 12256 20810 12308 20816
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 11978 19544 12034 19553
rect 11978 19479 12034 19488
rect 12084 19145 12112 20538
rect 12360 20534 12388 21422
rect 12714 21040 12770 21049
rect 12440 21004 12492 21010
rect 12714 20975 12770 20984
rect 12440 20946 12492 20952
rect 12452 20602 12480 20946
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12348 20528 12400 20534
rect 12348 20470 12400 20476
rect 12360 20380 12388 20470
rect 12544 20398 12572 20878
rect 12624 20800 12676 20806
rect 12622 20768 12624 20777
rect 12676 20768 12678 20777
rect 12622 20703 12678 20712
rect 12440 20392 12492 20398
rect 12360 20352 12440 20380
rect 12440 20334 12492 20340
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12622 20360 12678 20369
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12360 19990 12388 20198
rect 12348 19984 12400 19990
rect 12348 19926 12400 19932
rect 12348 19848 12400 19854
rect 12346 19816 12348 19825
rect 12400 19816 12402 19825
rect 12452 19786 12480 20334
rect 12622 20295 12678 20304
rect 12346 19751 12402 19760
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 19496 12296 19654
rect 12268 19468 12388 19496
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12070 19136 12126 19145
rect 12070 19071 12126 19080
rect 11978 19000 12034 19009
rect 11978 18935 12034 18944
rect 11886 16688 11942 16697
rect 11886 16623 11942 16632
rect 11900 15978 11928 16623
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11900 14414 11928 14758
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11900 13734 11928 14350
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11808 13382 11928 13410
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11808 12986 11836 13262
rect 11900 12986 11928 13382
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11992 11744 12020 18935
rect 12268 18834 12296 19314
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12268 18630 12296 18770
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 12084 17202 12112 17750
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12176 17270 12204 17546
rect 12164 17264 12216 17270
rect 12162 17232 12164 17241
rect 12216 17232 12218 17241
rect 12072 17196 12124 17202
rect 12162 17167 12218 17176
rect 12072 17138 12124 17144
rect 12070 17096 12126 17105
rect 12360 17066 12388 19468
rect 12438 19000 12494 19009
rect 12636 18986 12664 20295
rect 12728 19310 12756 20975
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12820 19174 12848 23423
rect 12912 20058 12940 24142
rect 13096 23730 13124 24618
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13082 22264 13138 22273
rect 12992 22228 13044 22234
rect 13082 22199 13138 22208
rect 12992 22170 13044 22176
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12912 19446 12940 19858
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12636 18958 12848 18986
rect 12438 18935 12494 18944
rect 12452 18737 12480 18935
rect 12438 18728 12494 18737
rect 12622 18728 12678 18737
rect 12438 18663 12494 18672
rect 12544 18686 12622 18714
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12452 17184 12480 18566
rect 12544 18057 12572 18686
rect 12622 18663 12678 18672
rect 12716 18624 12768 18630
rect 12622 18592 12678 18601
rect 12716 18566 12768 18572
rect 12622 18527 12678 18536
rect 12636 18358 12664 18527
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12530 18048 12586 18057
rect 12530 17983 12586 17992
rect 12530 17776 12586 17785
rect 12530 17711 12586 17720
rect 12544 17338 12572 17711
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12452 17156 12572 17184
rect 12070 17031 12126 17040
rect 12348 17060 12400 17066
rect 12084 15722 12112 17031
rect 12348 17002 12400 17008
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12452 16969 12480 17002
rect 12438 16960 12494 16969
rect 12438 16895 12494 16904
rect 12544 16810 12572 17156
rect 12452 16782 12572 16810
rect 12162 16552 12218 16561
rect 12162 16487 12218 16496
rect 12176 16250 12204 16487
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12176 15910 12204 16186
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12084 15694 12204 15722
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12084 14618 12112 14894
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12084 12238 12112 14214
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12084 11762 12112 12038
rect 11900 11716 12020 11744
rect 12072 11756 12124 11762
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11808 9178 11836 11494
rect 11900 11354 11928 11716
rect 12072 11698 12124 11704
rect 11980 11620 12032 11626
rect 11980 11562 12032 11568
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11900 9722 11928 9862
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11440 7126 11560 7154
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11334 6352 11390 6361
rect 11334 6287 11390 6296
rect 11440 5846 11468 7126
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11256 4826 11284 5646
rect 11440 5370 11468 5782
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11150 2000 11206 2009
rect 11150 1935 11206 1944
rect 11256 480 11284 4626
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11348 2009 11376 3878
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11440 2922 11468 3130
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 11440 2650 11468 2858
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11532 2038 11560 6054
rect 11624 5817 11652 6598
rect 11610 5808 11666 5817
rect 11610 5743 11666 5752
rect 11610 5672 11666 5681
rect 11610 5607 11666 5616
rect 11624 5370 11652 5607
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11716 5273 11744 7142
rect 11808 6497 11836 8774
rect 11900 7721 11928 9658
rect 11992 9654 12020 11562
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10538 12112 10950
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 12070 10296 12126 10305
rect 12070 10231 12126 10240
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 12084 9160 12112 10231
rect 11992 9132 12112 9160
rect 11992 8430 12020 9132
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11886 7712 11942 7721
rect 11886 7647 11942 7656
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11794 6488 11850 6497
rect 11794 6423 11850 6432
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11808 5681 11836 5782
rect 11794 5672 11850 5681
rect 11794 5607 11850 5616
rect 11702 5264 11758 5273
rect 11612 5228 11664 5234
rect 11702 5199 11758 5208
rect 11612 5170 11664 5176
rect 11624 4826 11652 5170
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11794 4040 11850 4049
rect 11900 4010 11928 7482
rect 11794 3975 11850 3984
rect 11888 4004 11940 4010
rect 11610 3632 11666 3641
rect 11610 3567 11612 3576
rect 11664 3567 11666 3576
rect 11612 3538 11664 3544
rect 11520 2032 11572 2038
rect 11334 2000 11390 2009
rect 11520 1974 11572 1980
rect 11334 1935 11390 1944
rect 11808 480 11836 3975
rect 11888 3946 11940 3952
rect 11992 2972 12020 8366
rect 12084 8090 12112 8978
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 4842 12204 15694
rect 12452 15366 12480 16782
rect 12532 16176 12584 16182
rect 12530 16144 12532 16153
rect 12584 16144 12586 16153
rect 12530 16079 12586 16088
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 12268 13870 12296 14826
rect 12452 14482 12480 15302
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12268 7970 12296 12174
rect 12360 11665 12388 13330
rect 12544 12345 12572 15030
rect 12636 14804 12664 18294
rect 12728 17202 12756 18566
rect 12820 17921 12848 18958
rect 12912 18698 12940 19246
rect 12900 18692 12952 18698
rect 12900 18634 12952 18640
rect 12806 17912 12862 17921
rect 12806 17847 12862 17856
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12820 17082 12848 17750
rect 12728 17054 12848 17082
rect 12728 16658 12756 17054
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12728 16153 12756 16594
rect 12714 16144 12770 16153
rect 12714 16079 12770 16088
rect 12714 15192 12770 15201
rect 12714 15127 12770 15136
rect 12728 14929 12756 15127
rect 12912 15026 12940 17818
rect 13004 17626 13032 22170
rect 13096 18358 13124 22199
rect 13188 20369 13216 26386
rect 13360 26376 13412 26382
rect 13360 26318 13412 26324
rect 13372 26081 13400 26318
rect 13358 26072 13414 26081
rect 13358 26007 13414 26016
rect 13268 25424 13320 25430
rect 13268 25366 13320 25372
rect 13280 24138 13308 25366
rect 13360 25356 13412 25362
rect 13360 25298 13412 25304
rect 13372 24614 13400 25298
rect 13648 24886 13676 27520
rect 13912 25968 13964 25974
rect 13912 25910 13964 25916
rect 13726 25392 13782 25401
rect 13726 25327 13782 25336
rect 13636 24880 13688 24886
rect 13636 24822 13688 24828
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13268 24132 13320 24138
rect 13268 24074 13320 24080
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 13280 23322 13308 23530
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 13280 22438 13308 23258
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13372 22250 13400 24550
rect 13452 24336 13504 24342
rect 13452 24278 13504 24284
rect 13464 23662 13492 24278
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 13452 23656 13504 23662
rect 13450 23624 13452 23633
rect 13504 23624 13506 23633
rect 13556 23594 13584 24074
rect 13450 23559 13506 23568
rect 13544 23588 13596 23594
rect 13544 23530 13596 23536
rect 13452 23520 13504 23526
rect 13452 23462 13504 23468
rect 13464 22574 13492 23462
rect 13740 23168 13768 25327
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 13832 24886 13860 25094
rect 13820 24880 13872 24886
rect 13820 24822 13872 24828
rect 13924 24596 13952 25910
rect 14096 25492 14148 25498
rect 14096 25434 14148 25440
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 14016 24750 14044 25094
rect 14108 24818 14136 25434
rect 14292 25378 14320 27520
rect 14464 26240 14516 26246
rect 14464 26182 14516 26188
rect 14292 25362 14412 25378
rect 14188 25356 14240 25362
rect 14292 25356 14424 25362
rect 14292 25350 14372 25356
rect 14188 25298 14240 25304
rect 14372 25298 14424 25304
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14004 24744 14056 24750
rect 14002 24712 14004 24721
rect 14056 24712 14058 24721
rect 14002 24647 14058 24656
rect 14200 24614 14228 25298
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14384 24993 14412 25094
rect 14370 24984 14426 24993
rect 14370 24919 14426 24928
rect 14280 24676 14332 24682
rect 14280 24618 14332 24624
rect 14188 24608 14240 24614
rect 13924 24568 14044 24596
rect 13910 24304 13966 24313
rect 13910 24239 13966 24248
rect 13924 23186 13952 24239
rect 13556 23140 13768 23168
rect 13912 23180 13964 23186
rect 13556 22658 13584 23140
rect 13912 23122 13964 23128
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13556 22630 13676 22658
rect 13452 22568 13504 22574
rect 13452 22510 13504 22516
rect 13280 22222 13400 22250
rect 13174 20360 13230 20369
rect 13174 20295 13230 20304
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13188 17785 13216 19654
rect 13280 19009 13308 22222
rect 13544 22092 13596 22098
rect 13544 22034 13596 22040
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 13266 19000 13322 19009
rect 13266 18935 13322 18944
rect 13266 18456 13322 18465
rect 13266 18391 13322 18400
rect 13280 17814 13308 18391
rect 13372 18290 13400 21626
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13464 20262 13492 21422
rect 13556 21010 13584 22034
rect 13648 21690 13676 22630
rect 13740 22506 13768 22918
rect 13832 22817 13860 23054
rect 13818 22808 13874 22817
rect 14016 22794 14044 24568
rect 14188 24550 14240 24556
rect 14016 22766 14136 22794
rect 13818 22743 13874 22752
rect 13728 22500 13780 22506
rect 13780 22460 13860 22488
rect 13728 22442 13780 22448
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13634 21584 13690 21593
rect 13634 21519 13690 21528
rect 13740 21536 13768 21966
rect 13832 21690 13860 22460
rect 13912 22160 13964 22166
rect 13912 22102 13964 22108
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13544 21004 13596 21010
rect 13544 20946 13596 20952
rect 13542 20360 13598 20369
rect 13542 20295 13598 20304
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13464 19514 13492 19994
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13464 18426 13492 18838
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13372 17882 13400 18226
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13268 17808 13320 17814
rect 13174 17776 13230 17785
rect 13464 17762 13492 18362
rect 13556 17882 13584 20295
rect 13648 20074 13676 21519
rect 13740 21508 13860 21536
rect 13832 20534 13860 21508
rect 13924 21146 13952 22102
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13924 20874 13952 21082
rect 13912 20868 13964 20874
rect 13912 20810 13964 20816
rect 14016 20806 14044 21966
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13648 20046 13860 20074
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13648 19174 13676 19790
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13740 19242 13768 19722
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13636 19168 13688 19174
rect 13634 19136 13636 19145
rect 13688 19136 13690 19145
rect 13634 19071 13690 19080
rect 13648 17921 13676 19071
rect 13740 18970 13768 19178
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13634 17912 13690 17921
rect 13544 17876 13596 17882
rect 13634 17847 13690 17856
rect 13544 17818 13596 17824
rect 13268 17750 13320 17756
rect 13174 17711 13230 17720
rect 13372 17734 13492 17762
rect 13004 17598 13308 17626
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 17066 13032 17478
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13096 16794 13124 17002
rect 13188 16794 13216 17138
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13096 16250 13124 16526
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12714 14920 12770 14929
rect 12714 14855 12770 14864
rect 12636 14776 12756 14804
rect 12530 12336 12586 12345
rect 12530 12271 12586 12280
rect 12544 12073 12572 12271
rect 12530 12064 12586 12073
rect 12530 11999 12586 12008
rect 12346 11656 12402 11665
rect 12346 11591 12402 11600
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12360 10452 12388 10678
rect 12452 10606 12480 11086
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12360 10424 12480 10452
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12360 9654 12388 10134
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 8838 12388 9454
rect 12452 9110 12480 10424
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12452 8634 12480 9046
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12438 8256 12494 8265
rect 12438 8191 12494 8200
rect 12268 7942 12388 7970
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7546 12296 7822
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12254 7304 12310 7313
rect 12254 7239 12256 7248
rect 12308 7239 12310 7248
rect 12256 7210 12308 7216
rect 12360 6746 12388 7942
rect 12452 7410 12480 8191
rect 12544 8090 12572 8298
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12544 7818 12572 8026
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12268 6718 12388 6746
rect 12438 6760 12494 6769
rect 12268 6322 12296 6718
rect 12438 6695 12494 6704
rect 12452 6662 12480 6695
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12176 4814 12296 4842
rect 12162 4720 12218 4729
rect 12268 4690 12296 4814
rect 12162 4655 12218 4664
rect 12256 4684 12308 4690
rect 12176 4554 12204 4655
rect 12256 4626 12308 4632
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12176 3097 12204 4218
rect 12268 4146 12296 4626
rect 12360 4536 12388 6598
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5953 12480 6054
rect 12438 5944 12494 5953
rect 12636 5914 12664 11222
rect 12438 5879 12494 5888
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12438 4992 12494 5001
rect 12438 4927 12494 4936
rect 12452 4729 12480 4927
rect 12438 4720 12494 4729
rect 12438 4655 12494 4664
rect 12440 4548 12492 4554
rect 12360 4508 12440 4536
rect 12440 4490 12492 4496
rect 12544 4321 12572 5238
rect 12636 5030 12664 5850
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12622 4720 12678 4729
rect 12622 4655 12678 4664
rect 12636 4622 12664 4655
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12530 4312 12586 4321
rect 12636 4282 12664 4558
rect 12530 4247 12586 4256
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12162 3088 12218 3097
rect 12162 3023 12218 3032
rect 11992 2944 12112 2972
rect 12084 2666 12112 2944
rect 12452 2802 12480 3334
rect 12728 2836 12756 14776
rect 12912 14362 12940 14962
rect 13174 14784 13230 14793
rect 13174 14719 13230 14728
rect 12912 14334 13032 14362
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 6984 12848 11494
rect 12912 7546 12940 14010
rect 13004 12986 13032 14334
rect 13188 14278 13216 14719
rect 13176 14272 13228 14278
rect 13082 14240 13138 14249
rect 13176 14214 13228 14220
rect 13082 14175 13138 14184
rect 13096 14074 13124 14175
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13188 13802 13216 14214
rect 13176 13796 13228 13802
rect 13176 13738 13228 13744
rect 13188 13530 13216 13738
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 13096 12714 13124 13262
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 13096 12306 13124 12650
rect 13280 12646 13308 17598
rect 13372 14249 13400 17734
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13464 16726 13492 17614
rect 13556 17338 13584 17818
rect 13634 17640 13690 17649
rect 13634 17575 13690 17584
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13464 16114 13492 16662
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13464 15706 13492 16050
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13556 15314 13584 17002
rect 13648 16590 13676 17575
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13634 16280 13690 16289
rect 13634 16215 13690 16224
rect 13648 15434 13676 16215
rect 13740 15745 13768 18566
rect 13832 16726 13860 20046
rect 14016 19174 14044 20742
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13832 16250 13860 16662
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13726 15736 13782 15745
rect 13726 15671 13782 15680
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13556 15286 13676 15314
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13464 14385 13492 14962
rect 13450 14376 13506 14385
rect 13450 14311 13506 14320
rect 13452 14272 13504 14278
rect 13358 14240 13414 14249
rect 13452 14214 13504 14220
rect 13358 14175 13414 14184
rect 13464 14090 13492 14214
rect 13372 14062 13492 14090
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13096 12186 13124 12242
rect 13004 12158 13124 12186
rect 13004 11286 13032 12158
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 13004 10810 13032 11222
rect 13096 11218 13124 12038
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13188 11354 13216 11630
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13004 10674 13032 10746
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13004 10130 13032 10610
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13096 10062 13124 11154
rect 13188 10742 13216 11290
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 10266 13216 10474
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13280 10198 13308 10950
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12992 8424 13044 8430
rect 13096 8401 13124 9318
rect 13188 8945 13216 9454
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13174 8936 13230 8945
rect 13174 8871 13230 8880
rect 12992 8366 13044 8372
rect 13082 8392 13138 8401
rect 13004 8022 13032 8366
rect 13082 8327 13138 8336
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 13004 7478 13032 7958
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12820 6956 12940 6984
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12820 6458 12848 6802
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5545 12848 6054
rect 12806 5536 12862 5545
rect 12806 5471 12862 5480
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12820 4282 12848 4762
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12912 3913 12940 6956
rect 13004 6934 13032 7414
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 13004 6458 13032 6870
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13004 6186 13032 6394
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 13096 6066 13124 8230
rect 13174 7712 13230 7721
rect 13174 7647 13230 7656
rect 13004 6038 13124 6066
rect 13004 5409 13032 6038
rect 13188 5642 13216 7647
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12990 5400 13046 5409
rect 12990 5335 13046 5344
rect 13004 5234 13032 5335
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13096 5098 13124 5510
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 13096 4865 13124 5034
rect 13082 4856 13138 4865
rect 13082 4791 13138 4800
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 12898 3904 12954 3913
rect 12898 3839 12954 3848
rect 13004 3738 13032 4558
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12530 2816 12586 2825
rect 12452 2774 12530 2802
rect 12084 2638 12296 2666
rect 12268 480 12296 2638
rect 12452 2553 12480 2774
rect 12530 2751 12586 2760
rect 12719 2808 12756 2836
rect 12719 2666 12747 2808
rect 12719 2638 12848 2666
rect 12438 2544 12494 2553
rect 12438 2479 12494 2488
rect 12820 480 12848 2638
rect 13280 2582 13308 9318
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13280 2310 13308 2518
rect 12900 2304 12952 2310
rect 13268 2304 13320 2310
rect 12900 2246 12952 2252
rect 13266 2272 13268 2281
rect 13320 2272 13322 2281
rect 12912 1465 12940 2246
rect 13266 2207 13322 2216
rect 12898 1456 12954 1465
rect 12898 1391 12954 1400
rect 13372 480 13400 14062
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13556 12986 13584 13126
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13556 12782 13584 12922
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 9722 13492 10542
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13556 9178 13584 12582
rect 13544 9172 13596 9178
rect 13464 9132 13544 9160
rect 13464 2990 13492 9132
rect 13544 9114 13596 9120
rect 13542 7984 13598 7993
rect 13542 7919 13598 7928
rect 13556 7478 13584 7919
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13556 7002 13584 7142
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 13556 5234 13584 6122
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13648 4826 13676 15286
rect 13832 15162 13860 15574
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13726 13424 13782 13433
rect 13726 13359 13782 13368
rect 13740 13258 13768 13359
rect 13924 13326 13952 18702
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 14016 14385 14044 18566
rect 14108 17218 14136 22766
rect 14200 17626 14228 24550
rect 14292 23769 14320 24618
rect 14370 24168 14426 24177
rect 14370 24103 14426 24112
rect 14278 23760 14334 23769
rect 14278 23695 14334 23704
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14292 21010 14320 21830
rect 14384 21146 14412 24103
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14292 19145 14320 20946
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14384 20058 14412 20198
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14384 19310 14412 19994
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14278 19136 14334 19145
rect 14278 19071 14334 19080
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14292 17746 14320 18226
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14200 17598 14412 17626
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14200 17338 14228 17478
rect 14384 17338 14412 17598
rect 14476 17354 14504 26182
rect 14556 25832 14608 25838
rect 14740 25832 14792 25838
rect 14608 25780 14688 25786
rect 14556 25774 14688 25780
rect 14740 25774 14792 25780
rect 14568 25758 14688 25774
rect 14554 24304 14610 24313
rect 14660 24290 14688 25758
rect 14752 25498 14780 25774
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 14844 25430 14872 27520
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 14832 25424 14884 25430
rect 14832 25366 14884 25372
rect 14936 25242 14964 25434
rect 14844 25214 14964 25242
rect 14844 24857 14872 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14830 24848 14886 24857
rect 14830 24783 14886 24792
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 14660 24262 14872 24290
rect 14554 24239 14556 24248
rect 14608 24239 14610 24248
rect 14556 24210 14608 24216
rect 14740 24132 14792 24138
rect 14740 24074 14792 24080
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 14568 21457 14596 23802
rect 14752 23594 14780 24074
rect 14740 23588 14792 23594
rect 14740 23530 14792 23536
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14660 21593 14688 22918
rect 14752 22778 14780 23530
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14844 22574 14872 24262
rect 15212 24052 15240 24618
rect 15304 24562 15332 24754
rect 15396 24750 15424 27520
rect 15660 25968 15712 25974
rect 15660 25910 15712 25916
rect 15750 25936 15806 25945
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15580 25401 15608 25434
rect 15566 25392 15622 25401
rect 15476 25356 15528 25362
rect 15566 25327 15622 25336
rect 15476 25298 15528 25304
rect 15384 24744 15436 24750
rect 15384 24686 15436 24692
rect 15304 24534 15424 24562
rect 15212 24024 15332 24052
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23594 15332 24024
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15396 23474 15424 24534
rect 15488 24410 15516 25298
rect 15672 24886 15700 25910
rect 15750 25871 15806 25880
rect 15568 24880 15620 24886
rect 15568 24822 15620 24828
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15212 23446 15424 23474
rect 15106 23080 15162 23089
rect 15106 23015 15108 23024
rect 15160 23015 15162 23024
rect 15108 22986 15160 22992
rect 15212 22964 15240 23446
rect 15382 23352 15438 23361
rect 15382 23287 15438 23296
rect 15396 23050 15424 23287
rect 15488 23254 15516 24346
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15384 23044 15436 23050
rect 15384 22986 15436 22992
rect 15212 22936 15332 22964
rect 15304 22930 15332 22936
rect 15304 22902 15424 22930
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14832 22568 14884 22574
rect 14832 22510 14884 22516
rect 15396 22250 15424 22902
rect 15488 22778 15516 23190
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15304 22222 15424 22250
rect 15304 22137 15332 22222
rect 15290 22128 15346 22137
rect 15290 22063 15346 22072
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15108 22024 15160 22030
rect 15106 21992 15108 22001
rect 15160 21992 15162 22001
rect 15106 21927 15162 21936
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15396 21729 15424 22034
rect 15382 21720 15438 21729
rect 15382 21655 15384 21664
rect 15436 21655 15438 21664
rect 15384 21626 15436 21632
rect 14646 21584 14702 21593
rect 14646 21519 14702 21528
rect 14554 21448 14610 21457
rect 14554 21383 14610 21392
rect 14660 20942 14688 21519
rect 14832 21480 14884 21486
rect 14830 21448 14832 21457
rect 14884 21448 14886 21457
rect 14830 21383 14886 21392
rect 15014 21176 15070 21185
rect 15014 21111 15016 21120
rect 15068 21111 15070 21120
rect 15382 21176 15438 21185
rect 15382 21111 15438 21120
rect 15016 21082 15068 21088
rect 14832 21072 14884 21078
rect 14832 21014 14884 21020
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14738 20632 14794 20641
rect 14844 20602 14872 21014
rect 15290 20904 15346 20913
rect 15290 20839 15346 20848
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14738 20567 14794 20576
rect 14832 20596 14884 20602
rect 14646 20496 14702 20505
rect 14752 20466 14780 20567
rect 14832 20538 14884 20544
rect 14646 20431 14702 20440
rect 14740 20460 14792 20466
rect 14660 20058 14688 20431
rect 14740 20402 14792 20408
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 15304 19990 15332 20839
rect 15396 20466 15424 21111
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15488 20330 15516 22714
rect 15580 22098 15608 24822
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15672 23769 15700 24550
rect 15764 24290 15792 25871
rect 15844 25424 15896 25430
rect 15844 25366 15896 25372
rect 15856 24410 15884 25366
rect 15948 24954 15976 27520
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 16118 26344 16174 26353
rect 16040 25945 16068 26318
rect 16118 26279 16174 26288
rect 16026 25936 16082 25945
rect 16026 25871 16082 25880
rect 16028 25152 16080 25158
rect 16028 25094 16080 25100
rect 16040 24993 16068 25094
rect 16026 24984 16082 24993
rect 15936 24948 15988 24954
rect 16026 24919 16082 24928
rect 15936 24890 15988 24896
rect 16132 24886 16160 26279
rect 16120 24880 16172 24886
rect 16120 24822 16172 24828
rect 16396 24744 16448 24750
rect 16396 24686 16448 24692
rect 16026 24440 16082 24449
rect 15844 24404 15896 24410
rect 16026 24375 16082 24384
rect 16120 24404 16172 24410
rect 15844 24346 15896 24352
rect 15764 24262 15976 24290
rect 15750 23896 15806 23905
rect 15750 23831 15752 23840
rect 15804 23831 15806 23840
rect 15752 23802 15804 23808
rect 15658 23760 15714 23769
rect 15658 23695 15714 23704
rect 15752 23588 15804 23594
rect 15752 23530 15804 23536
rect 15658 22128 15714 22137
rect 15568 22092 15620 22098
rect 15658 22063 15714 22072
rect 15568 22034 15620 22040
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15580 21570 15608 21830
rect 15672 21690 15700 22063
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15580 21542 15700 21570
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 20324 15528 20330
rect 15476 20266 15528 20272
rect 15488 20058 15516 20266
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15292 19984 15344 19990
rect 14738 19952 14794 19961
rect 15292 19926 15344 19932
rect 14738 19887 14794 19896
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14568 19242 14596 19450
rect 14648 19440 14700 19446
rect 14646 19408 14648 19417
rect 14700 19408 14702 19417
rect 14646 19343 14702 19352
rect 14556 19236 14608 19242
rect 14556 19178 14608 19184
rect 14568 18426 14596 19178
rect 14752 18465 14780 19887
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15382 19544 15438 19553
rect 15382 19479 15438 19488
rect 15396 19446 15424 19479
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15382 19272 15438 19281
rect 15382 19207 15438 19216
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15106 18864 15162 18873
rect 15106 18799 15108 18808
rect 15160 18799 15162 18808
rect 15108 18770 15160 18776
rect 14830 18728 14886 18737
rect 15212 18714 15240 19110
rect 14886 18686 15240 18714
rect 15396 18698 15424 19207
rect 15384 18692 15436 18698
rect 14830 18663 14886 18672
rect 15384 18634 15436 18640
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14738 18456 14794 18465
rect 14556 18420 14608 18426
rect 14956 18448 15252 18468
rect 15382 18456 15438 18465
rect 14738 18391 14794 18400
rect 15292 18420 15344 18426
rect 14556 18362 14608 18368
rect 15382 18391 15438 18400
rect 15292 18362 15344 18368
rect 15304 18306 15332 18362
rect 15120 18278 15332 18306
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14568 17746 14596 18090
rect 15120 17882 15148 18278
rect 15396 18086 15424 18391
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14738 17504 14794 17513
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14372 17332 14424 17338
rect 14476 17326 14596 17354
rect 14372 17274 14424 17280
rect 14108 17190 14504 17218
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 14108 15706 14136 16458
rect 14200 16425 14228 16934
rect 14384 16454 14412 17002
rect 14372 16448 14424 16454
rect 14186 16416 14242 16425
rect 14372 16390 14424 16396
rect 14186 16351 14242 16360
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14094 15328 14150 15337
rect 14094 15263 14150 15272
rect 14108 15162 14136 15263
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14002 14376 14058 14385
rect 14002 14311 14058 14320
rect 14016 13530 14044 14311
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13910 13152 13966 13161
rect 13910 13087 13966 13096
rect 13924 12918 13952 13087
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13924 12714 13952 12854
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 14108 12594 14136 13398
rect 13924 12566 14136 12594
rect 13728 12368 13780 12374
rect 13780 12316 13860 12322
rect 13728 12310 13860 12316
rect 13740 12294 13860 12310
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 9994 13768 12174
rect 13832 10742 13860 12294
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13832 9874 13860 10134
rect 13740 9846 13860 9874
rect 13740 9382 13768 9846
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13728 9376 13780 9382
rect 13832 9353 13860 9454
rect 13728 9318 13780 9324
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13924 8945 13952 12566
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14016 11898 14044 12174
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 14200 11665 14228 16186
rect 14384 15881 14412 16186
rect 14370 15872 14426 15881
rect 14370 15807 14426 15816
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14292 14278 14320 14758
rect 14384 14346 14412 14826
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14370 12880 14426 12889
rect 14370 12815 14426 12824
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14292 12102 14320 12718
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14186 11656 14242 11665
rect 14016 11614 14186 11642
rect 13910 8936 13966 8945
rect 13910 8871 13966 8880
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13832 7970 13860 8502
rect 13740 7954 13860 7970
rect 13728 7948 13860 7954
rect 13780 7942 13860 7948
rect 14016 7936 14044 11614
rect 14292 11626 14320 12038
rect 14186 11591 14242 11600
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14108 9761 14136 9930
rect 14094 9752 14150 9761
rect 14094 9687 14150 9696
rect 13728 7890 13780 7896
rect 13924 7908 14044 7936
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13634 3496 13690 3505
rect 13634 3431 13636 3440
rect 13688 3431 13690 3440
rect 13636 3402 13688 3408
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13648 1601 13676 2246
rect 13634 1592 13690 1601
rect 13634 1527 13690 1536
rect 4434 368 4490 377
rect 4434 303 4490 312
rect 4894 0 4950 480
rect 5446 0 5502 480
rect 5998 0 6054 480
rect 6458 0 6514 480
rect 7010 0 7066 480
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8574 0 8630 480
rect 9126 0 9182 480
rect 9678 0 9734 480
rect 10138 0 10194 480
rect 10690 0 10746 480
rect 11242 0 11298 480
rect 11794 0 11850 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13740 241 13768 7482
rect 13832 6934 13860 7754
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6186 13860 6598
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13832 5914 13860 6122
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13832 4758 13860 5714
rect 13924 5710 13952 7908
rect 14108 7834 14136 9687
rect 14200 8820 14228 9998
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14292 9353 14320 9522
rect 14278 9344 14334 9353
rect 14278 9279 14334 9288
rect 14384 8922 14412 12815
rect 14476 12306 14504 17190
rect 14568 15638 14596 17326
rect 14660 16794 14688 17478
rect 14738 17439 14794 17448
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14660 15586 14688 15982
rect 14752 15706 14780 17439
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14568 14074 14596 15574
rect 14660 15558 14780 15586
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14660 15201 14688 15438
rect 14646 15192 14702 15201
rect 14646 15127 14702 15136
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14660 14113 14688 14826
rect 14752 14482 14780 15558
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14646 14104 14702 14113
rect 14556 14068 14608 14074
rect 14646 14039 14702 14048
rect 14556 14010 14608 14016
rect 14752 13841 14780 14214
rect 14738 13832 14794 13841
rect 14738 13767 14794 13776
rect 14740 13388 14792 13394
rect 14660 13348 14740 13376
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 12850 14596 13262
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14660 12764 14688 13348
rect 14740 13330 14792 13336
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14752 12889 14780 13194
rect 14738 12880 14794 12889
rect 14738 12815 14794 12824
rect 14660 12736 14780 12764
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14476 9654 14504 12242
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14568 11014 14596 11562
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14568 10606 14596 10950
rect 14646 10840 14702 10849
rect 14646 10775 14648 10784
rect 14700 10775 14702 10784
rect 14648 10746 14700 10752
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14568 10062 14596 10542
rect 14660 10470 14688 10746
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14568 9450 14596 9998
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14384 8894 14504 8922
rect 14568 8906 14596 9386
rect 14280 8832 14332 8838
rect 14200 8792 14280 8820
rect 14280 8774 14332 8780
rect 14370 8800 14426 8809
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14016 7806 14136 7834
rect 14016 7342 14044 7806
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14108 7154 14136 7686
rect 14016 7126 14136 7154
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13924 5370 13952 5646
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13912 5024 13964 5030
rect 14016 5001 14044 7126
rect 14096 6724 14148 6730
rect 14096 6666 14148 6672
rect 13912 4966 13964 4972
rect 14002 4992 14058 5001
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 13832 4146 13860 4490
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13924 3777 13952 4966
rect 14002 4927 14058 4936
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 4146 14044 4422
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 14108 4010 14136 6666
rect 14200 4282 14228 8298
rect 14292 7970 14320 8774
rect 14370 8735 14426 8744
rect 14384 8634 14412 8735
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14476 8090 14504 8894
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14648 8832 14700 8838
rect 14554 8800 14610 8809
rect 14648 8774 14700 8780
rect 14554 8735 14610 8744
rect 14568 8566 14596 8735
rect 14660 8673 14688 8774
rect 14646 8664 14702 8673
rect 14646 8599 14702 8608
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14292 7942 14504 7970
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14384 7002 14412 7278
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14370 6896 14426 6905
rect 14370 6831 14426 6840
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14096 4004 14148 4010
rect 14096 3946 14148 3952
rect 14200 3777 14228 4218
rect 13910 3768 13966 3777
rect 13910 3703 13966 3712
rect 14186 3768 14242 3777
rect 14186 3703 14242 3712
rect 13818 3632 13874 3641
rect 13818 3567 13874 3576
rect 13832 2854 13860 3567
rect 14096 3528 14148 3534
rect 13910 3496 13966 3505
rect 13910 3431 13966 3440
rect 14094 3496 14096 3505
rect 14148 3496 14150 3505
rect 14094 3431 14150 3440
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13924 480 13952 3431
rect 14292 2650 14320 6666
rect 14384 6458 14412 6831
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14384 5370 14412 5714
rect 14476 5556 14504 7942
rect 14568 5846 14596 8502
rect 14752 6730 14780 12736
rect 14844 11642 14872 17274
rect 14922 17232 14978 17241
rect 14922 17167 14978 17176
rect 14936 16658 14964 17167
rect 15014 16960 15070 16969
rect 15014 16895 15070 16904
rect 15028 16794 15056 16895
rect 15488 16833 15516 18566
rect 15474 16824 15530 16833
rect 15016 16788 15068 16794
rect 15474 16759 15530 16768
rect 15016 16730 15068 16736
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15382 16280 15438 16289
rect 15382 16215 15438 16224
rect 15396 16046 15424 16215
rect 15474 16144 15530 16153
rect 15474 16079 15530 16088
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 14924 15972 14976 15978
rect 14924 15914 14976 15920
rect 14936 15881 14964 15914
rect 15200 15904 15252 15910
rect 14922 15872 14978 15881
rect 15200 15846 15252 15852
rect 14922 15807 14978 15816
rect 14936 15570 14964 15807
rect 15212 15638 15240 15846
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15198 15056 15254 15065
rect 15198 14991 15254 15000
rect 15212 14550 15240 14991
rect 15396 14822 15424 15506
rect 15384 14816 15436 14822
rect 15382 14784 15384 14793
rect 15436 14784 15438 14793
rect 15382 14719 15438 14728
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15200 14340 15252 14346
rect 15252 14300 15332 14328
rect 15200 14282 15252 14288
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15106 12608 15162 12617
rect 15106 12543 15162 12552
rect 14924 12232 14976 12238
rect 14922 12200 14924 12209
rect 15120 12209 15148 12543
rect 14976 12200 14978 12209
rect 14922 12135 14978 12144
rect 15106 12200 15162 12209
rect 15106 12135 15162 12144
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14844 11614 14964 11642
rect 14830 11520 14886 11529
rect 14830 11455 14886 11464
rect 14844 10538 14872 11455
rect 14936 11082 14964 11614
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14844 9926 14872 10474
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14752 5914 14780 6394
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14556 5840 14608 5846
rect 14556 5782 14608 5788
rect 14476 5528 14688 5556
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14476 4826 14504 5102
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14476 4214 14504 4490
rect 14568 4282 14596 4626
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14464 4208 14516 4214
rect 14660 4162 14688 5528
rect 14752 5098 14780 5850
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14844 4978 14872 8026
rect 14922 7848 14978 7857
rect 14922 7783 14924 7792
rect 14976 7783 14978 7792
rect 14924 7754 14976 7760
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7562 15332 14300
rect 15396 13734 15424 14418
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15396 10674 15424 11766
rect 15488 11234 15516 16079
rect 15580 11626 15608 20402
rect 15672 20369 15700 21542
rect 15764 21078 15792 23530
rect 15948 23322 15976 24262
rect 15936 23316 15988 23322
rect 15936 23258 15988 23264
rect 15844 23248 15896 23254
rect 15844 23190 15896 23196
rect 15856 22438 15884 23190
rect 15936 22976 15988 22982
rect 15936 22918 15988 22924
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15856 21146 15884 22374
rect 15948 21894 15976 22918
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15752 21072 15804 21078
rect 15752 21014 15804 21020
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15658 20360 15714 20369
rect 15658 20295 15714 20304
rect 15764 20262 15792 20878
rect 15856 20602 15884 21082
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15948 20482 15976 21558
rect 15856 20454 15976 20482
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 20058 15792 20198
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15750 19952 15806 19961
rect 15750 19887 15806 19896
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15672 17678 15700 18770
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15672 15910 15700 16458
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15658 15736 15714 15745
rect 15658 15671 15714 15680
rect 15672 15638 15700 15671
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 15658 15328 15714 15337
rect 15658 15263 15714 15272
rect 15672 15026 15700 15263
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15672 13394 15700 14486
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15764 13258 15792 19887
rect 15856 18737 15884 20454
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15948 19514 15976 19790
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 15948 18834 15976 19246
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15842 18728 15898 18737
rect 15842 18663 15898 18672
rect 15948 18426 15976 18770
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16040 17882 16068 24375
rect 16120 24346 16172 24352
rect 16132 21622 16160 24346
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16224 23526 16252 24142
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16212 23520 16264 23526
rect 16210 23488 16212 23497
rect 16264 23488 16266 23497
rect 16210 23423 16266 23432
rect 16212 23316 16264 23322
rect 16212 23258 16264 23264
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16132 20346 16160 21286
rect 16224 20466 16252 23258
rect 16316 21457 16344 24006
rect 16408 21865 16436 24686
rect 16500 24585 16528 27520
rect 17052 26110 17080 27520
rect 17604 26858 17632 27520
rect 17592 26852 17644 26858
rect 17592 26794 17644 26800
rect 17314 26480 17370 26489
rect 17314 26415 17370 26424
rect 17040 26104 17092 26110
rect 17040 26046 17092 26052
rect 16672 25288 16724 25294
rect 17328 25265 17356 26415
rect 17868 25968 17920 25974
rect 17788 25928 17868 25956
rect 16672 25230 16724 25236
rect 17314 25256 17370 25265
rect 16486 24576 16542 24585
rect 16486 24511 16542 24520
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16500 22778 16528 23598
rect 16592 23322 16620 24210
rect 16684 23905 16712 25230
rect 17314 25191 17370 25200
rect 17500 25220 17552 25226
rect 17500 25162 17552 25168
rect 17512 24954 17540 25162
rect 17500 24948 17552 24954
rect 17500 24890 17552 24896
rect 16762 24848 16818 24857
rect 16762 24783 16818 24792
rect 16670 23896 16726 23905
rect 16670 23831 16726 23840
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16500 21962 16528 22442
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16394 21856 16450 21865
rect 16394 21791 16450 21800
rect 16302 21448 16358 21457
rect 16302 21383 16358 21392
rect 16316 21078 16344 21383
rect 16408 21185 16436 21791
rect 16500 21690 16528 21898
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16592 21486 16620 23258
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16486 21312 16542 21321
rect 16486 21247 16542 21256
rect 16394 21176 16450 21185
rect 16394 21111 16450 21120
rect 16304 21072 16356 21078
rect 16304 21014 16356 21020
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16394 20360 16450 20369
rect 16132 20318 16344 20346
rect 16210 20224 16266 20233
rect 16210 20159 16266 20168
rect 16120 19712 16172 19718
rect 16120 19654 16172 19660
rect 16132 19417 16160 19654
rect 16224 19514 16252 20159
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16118 19408 16174 19417
rect 16118 19343 16120 19352
rect 16172 19343 16174 19352
rect 16120 19314 16172 19320
rect 16132 19283 16160 19314
rect 16212 18896 16264 18902
rect 16212 18838 16264 18844
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 15842 17776 15898 17785
rect 15842 17711 15898 17720
rect 15856 16794 15884 17711
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 15948 17270 15976 17546
rect 16026 17368 16082 17377
rect 16026 17303 16082 17312
rect 15936 17264 15988 17270
rect 15934 17232 15936 17241
rect 15988 17232 15990 17241
rect 15934 17167 15990 17176
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 16040 16454 16068 17303
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 16040 16250 16068 16390
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15856 15473 15884 15574
rect 15842 15464 15898 15473
rect 15842 15399 15898 15408
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15672 12442 15700 12786
rect 15764 12442 15792 12922
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15856 12238 15884 13670
rect 15936 13456 15988 13462
rect 15934 13424 15936 13433
rect 15988 13424 15990 13433
rect 15934 13359 15990 13368
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16040 12986 16068 13262
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15844 12232 15896 12238
rect 15658 12200 15714 12209
rect 15844 12174 15896 12180
rect 15658 12135 15714 12144
rect 15672 11665 15700 12135
rect 15752 11688 15804 11694
rect 15658 11656 15714 11665
rect 15568 11620 15620 11626
rect 15856 11676 15884 12174
rect 15804 11648 15884 11676
rect 15752 11630 15804 11636
rect 15658 11591 15714 11600
rect 15568 11562 15620 11568
rect 15856 11354 15884 11648
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15488 11206 15700 11234
rect 15476 11144 15528 11150
rect 15474 11112 15476 11121
rect 15528 11112 15530 11121
rect 15474 11047 15530 11056
rect 15568 11008 15620 11014
rect 15474 10976 15530 10985
rect 15568 10950 15620 10956
rect 15474 10911 15530 10920
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15396 9042 15424 10066
rect 15488 9994 15516 10911
rect 15580 10538 15608 10950
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 10198 15608 10474
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15568 9920 15620 9926
rect 15566 9888 15568 9897
rect 15620 9888 15622 9897
rect 15566 9823 15622 9832
rect 15580 9518 15608 9823
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15384 9036 15436 9042
rect 15488 9024 15516 9454
rect 15568 9036 15620 9042
rect 15488 8996 15568 9024
rect 15384 8978 15436 8984
rect 15568 8978 15620 8984
rect 15580 8634 15608 8978
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15304 7534 15608 7562
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 14922 7032 14978 7041
rect 14922 6967 14978 6976
rect 14936 6934 14964 6967
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 15120 6882 15148 7142
rect 15212 7002 15240 7210
rect 15384 7200 15436 7206
rect 15382 7168 15384 7177
rect 15436 7168 15438 7177
rect 15382 7103 15438 7112
rect 15200 6996 15252 7002
rect 15252 6956 15332 6984
rect 15200 6938 15252 6944
rect 15120 6854 15240 6882
rect 15212 6798 15240 6854
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14844 4950 15240 4978
rect 15212 4826 15240 4950
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 14752 4282 14780 4762
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14464 4150 14516 4156
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14384 3194 14412 3470
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14384 480 14412 2994
rect 14476 1601 14504 4150
rect 14568 4134 14688 4162
rect 14568 3058 14596 4134
rect 14752 4078 14780 4218
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14646 3632 14702 3641
rect 14646 3567 14648 3576
rect 14700 3567 14702 3576
rect 14648 3538 14700 3544
rect 14752 3194 14780 4014
rect 15304 3942 15332 6956
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 6118 15424 6802
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15488 6361 15516 6598
rect 15474 6352 15530 6361
rect 15474 6287 15530 6296
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 4758 15424 4966
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15396 3738 15424 4694
rect 15474 3904 15530 3913
rect 15474 3839 15530 3848
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14554 2952 14610 2961
rect 14554 2887 14610 2896
rect 14568 2854 14596 2887
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14752 2582 14780 3130
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14646 2136 14702 2145
rect 14646 2071 14648 2080
rect 14700 2071 14702 2080
rect 14648 2042 14700 2048
rect 14752 1737 14780 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14554 1728 14610 1737
rect 14554 1663 14610 1672
rect 14738 1728 14794 1737
rect 14738 1663 14794 1672
rect 14462 1592 14518 1601
rect 14568 1578 14596 1663
rect 14568 1550 15056 1578
rect 14462 1527 14518 1536
rect 14922 1456 14978 1465
rect 15028 1442 15056 1550
rect 15106 1456 15162 1465
rect 15028 1414 15106 1442
rect 14922 1391 14978 1400
rect 15106 1391 15162 1400
rect 14936 480 14964 1391
rect 15304 1193 15332 3334
rect 15396 2922 15424 3674
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15290 1184 15346 1193
rect 15290 1119 15346 1128
rect 15488 480 15516 3839
rect 13726 232 13782 241
rect 13726 167 13782 176
rect 13910 0 13966 480
rect 14370 0 14426 480
rect 14922 0 14978 480
rect 15474 0 15530 480
rect 15580 377 15608 7534
rect 15672 5778 15700 11206
rect 15856 10810 15884 11290
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15764 8945 15792 10134
rect 15856 9450 15884 10746
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 16132 9382 16160 18226
rect 16224 18086 16252 18838
rect 16316 18290 16344 20318
rect 16500 20346 16528 21247
rect 16500 20318 16620 20346
rect 16394 20295 16450 20304
rect 16408 20244 16436 20295
rect 16408 20216 16528 20244
rect 16500 19990 16528 20216
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16212 18080 16264 18086
rect 16210 18048 16212 18057
rect 16264 18048 16266 18057
rect 16210 17983 16266 17992
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16224 17338 16252 17682
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16408 16674 16436 19858
rect 16500 18970 16528 19926
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16592 17746 16620 20318
rect 16684 20262 16712 23462
rect 16776 22953 16804 24783
rect 16856 24676 16908 24682
rect 16856 24618 16908 24624
rect 16868 24410 16896 24618
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16948 24336 17000 24342
rect 16948 24278 17000 24284
rect 16854 23080 16910 23089
rect 16960 23050 16988 24278
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17604 23662 17632 24006
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 17408 23248 17460 23254
rect 17408 23190 17460 23196
rect 17590 23216 17646 23225
rect 16854 23015 16910 23024
rect 16948 23044 17000 23050
rect 16762 22944 16818 22953
rect 16762 22879 16818 22888
rect 16764 22704 16816 22710
rect 16764 22646 16816 22652
rect 16776 21418 16804 22646
rect 16868 22506 16896 23015
rect 16948 22986 17000 22992
rect 17420 22778 17448 23190
rect 17590 23151 17646 23160
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16776 20602 16804 21082
rect 16868 20874 16896 22442
rect 17224 22432 17276 22438
rect 17224 22374 17276 22380
rect 17236 22234 17264 22374
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17132 22092 17184 22098
rect 17132 22034 17184 22040
rect 17038 21992 17094 22001
rect 17038 21927 17094 21936
rect 16948 21684 17000 21690
rect 16948 21626 17000 21632
rect 16960 21486 16988 21626
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16868 20398 16896 20470
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16316 16646 16436 16674
rect 16488 16652 16540 16658
rect 16210 16008 16266 16017
rect 16210 15943 16266 15952
rect 16224 14006 16252 15943
rect 16316 14056 16344 16646
rect 16488 16594 16540 16600
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16408 15910 16436 16526
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16408 15570 16436 15846
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16500 15434 16528 16594
rect 16488 15428 16540 15434
rect 16488 15370 16540 15376
rect 16488 14068 16540 14074
rect 16316 14028 16436 14056
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16302 13968 16358 13977
rect 16302 13903 16304 13912
rect 16356 13903 16358 13912
rect 16304 13874 16356 13880
rect 16408 12374 16436 14028
rect 16592 14056 16620 17478
rect 16684 17134 16712 20198
rect 16960 20058 16988 21422
rect 17052 21350 17080 21927
rect 17144 21690 17172 22034
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 17236 21690 17264 21830
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17052 21049 17080 21286
rect 17038 21040 17094 21049
rect 17038 20975 17094 20984
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17144 19258 17172 21354
rect 17328 21078 17356 21830
rect 17316 21072 17368 21078
rect 17316 21014 17368 21020
rect 17328 20505 17356 21014
rect 17420 20924 17448 22714
rect 17500 22568 17552 22574
rect 17500 22510 17552 22516
rect 17512 21690 17540 22510
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17512 21078 17540 21422
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17420 20896 17540 20924
rect 17314 20496 17370 20505
rect 17314 20431 17370 20440
rect 16776 19230 17172 19258
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16776 16640 16804 19230
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16946 19136 17002 19145
rect 16684 16612 16804 16640
rect 16684 15502 16712 16612
rect 16762 16552 16818 16561
rect 16762 16487 16818 16496
rect 16776 15881 16804 16487
rect 16762 15872 16818 15881
rect 16762 15807 16818 15816
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16684 15026 16712 15302
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16540 14028 16620 14056
rect 16488 14010 16540 14016
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16500 13530 16528 13738
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16500 13297 16528 13330
rect 16486 13288 16542 13297
rect 16486 13223 16542 13232
rect 16500 12986 16528 13223
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16592 12646 16620 14028
rect 16684 13410 16712 14826
rect 16776 14618 16804 15807
rect 16868 15473 16896 19110
rect 16946 19071 17002 19080
rect 16960 18698 16988 19071
rect 17038 18728 17094 18737
rect 16948 18692 17000 18698
rect 17038 18663 17094 18672
rect 16948 18634 17000 18640
rect 17052 18426 17080 18663
rect 17130 18456 17186 18465
rect 17040 18420 17092 18426
rect 17130 18391 17186 18400
rect 17040 18362 17092 18368
rect 16946 17640 17002 17649
rect 16946 17575 17002 17584
rect 16960 17066 16988 17575
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16854 15464 16910 15473
rect 16854 15399 16910 15408
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16762 14376 16818 14385
rect 16762 14311 16818 14320
rect 16776 14278 16804 14311
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16868 14113 16896 15302
rect 16960 15162 16988 17002
rect 17052 16697 17080 17070
rect 17038 16688 17094 16697
rect 17038 16623 17094 16632
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16946 14920 17002 14929
rect 16946 14855 16948 14864
rect 17000 14855 17002 14864
rect 16948 14826 17000 14832
rect 17052 14521 17080 14962
rect 17038 14512 17094 14521
rect 17038 14447 17094 14456
rect 16946 14376 17002 14385
rect 16946 14311 17002 14320
rect 16854 14104 16910 14113
rect 16854 14039 16910 14048
rect 16960 13938 16988 14311
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 17144 13802 17172 18391
rect 17236 17746 17264 19246
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17328 18068 17356 18702
rect 17420 18290 17448 18838
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17408 18080 17460 18086
rect 17328 18040 17408 18068
rect 17408 18022 17460 18028
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17236 17270 17264 17682
rect 17224 17264 17276 17270
rect 17276 17224 17356 17252
rect 17224 17206 17276 17212
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 17236 16250 17264 16662
rect 17328 16658 17356 17224
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17328 16250 17356 16594
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17420 15858 17448 18022
rect 17328 15830 17448 15858
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 13938 17264 14826
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16762 13560 16818 13569
rect 16762 13495 16764 13504
rect 16816 13495 16818 13504
rect 16764 13466 16816 13472
rect 16684 13382 16804 13410
rect 16868 13394 16896 13670
rect 17236 13462 17264 13874
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 16776 13161 16804 13382
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16762 13152 16818 13161
rect 16762 13087 16818 13096
rect 16776 12782 16804 13087
rect 17236 12918 17264 13398
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16304 11756 16356 11762
rect 16408 11744 16436 12310
rect 16356 11716 16436 11744
rect 16304 11698 16356 11704
rect 16394 11656 16450 11665
rect 16394 11591 16450 11600
rect 16408 10810 16436 11591
rect 16500 11286 16528 12378
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16500 11098 16528 11222
rect 16500 11070 16620 11098
rect 16592 10810 16620 11070
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16684 10606 16712 11562
rect 16856 11552 16908 11558
rect 16908 11512 16988 11540
rect 16856 11494 16908 11500
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 16408 10305 16436 10474
rect 16394 10296 16450 10305
rect 16868 10266 16896 10610
rect 16394 10231 16396 10240
rect 16448 10231 16450 10240
rect 16856 10260 16908 10266
rect 16396 10202 16448 10208
rect 16856 10202 16908 10208
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 15750 8936 15806 8945
rect 15750 8871 15806 8880
rect 15764 8634 15792 8871
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15948 7546 15976 8774
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 16040 7993 16068 8298
rect 16026 7984 16082 7993
rect 16026 7919 16082 7928
rect 16132 7834 16160 9318
rect 16500 9160 16528 10066
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16580 9172 16632 9178
rect 16500 9132 16580 9160
rect 16580 9114 16632 9120
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16210 8664 16266 8673
rect 16210 8599 16266 8608
rect 16224 8362 16252 8599
rect 16316 8498 16344 9046
rect 16672 8560 16724 8566
rect 16670 8528 16672 8537
rect 16724 8528 16726 8537
rect 16304 8492 16356 8498
rect 16670 8463 16726 8472
rect 16304 8434 16356 8440
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16316 8090 16344 8434
rect 16394 8392 16450 8401
rect 16394 8327 16450 8336
rect 16672 8356 16724 8362
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16132 7806 16252 7834
rect 16120 7744 16172 7750
rect 16118 7712 16120 7721
rect 16172 7712 16174 7721
rect 16118 7647 16174 7656
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15750 7168 15806 7177
rect 15750 7103 15806 7112
rect 15764 6458 15792 7103
rect 16224 6934 16252 7806
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15856 6458 15884 6802
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 16040 6254 16068 6734
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16302 6216 16358 6225
rect 16040 5914 16068 6190
rect 16302 6151 16358 6160
rect 16316 5914 16344 6151
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 15658 4992 15714 5001
rect 15658 4927 15714 4936
rect 15672 4758 15700 4927
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15658 3768 15714 3777
rect 15856 3738 15884 4490
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15658 3703 15714 3712
rect 15844 3732 15896 3738
rect 15672 3670 15700 3703
rect 15844 3674 15896 3680
rect 15948 3670 15976 3878
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15948 3194 15976 3606
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15660 2100 15712 2106
rect 15660 2042 15712 2048
rect 15672 1873 15700 2042
rect 15764 2009 15792 2450
rect 15750 2000 15806 2009
rect 15750 1935 15806 1944
rect 15658 1864 15714 1873
rect 15658 1799 15714 1808
rect 16040 480 16068 5510
rect 16316 4690 16344 5850
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16408 4321 16436 8327
rect 16672 8298 16724 8304
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16488 6792 16540 6798
rect 16486 6760 16488 6769
rect 16540 6760 16542 6769
rect 16486 6695 16542 6704
rect 16486 5672 16542 5681
rect 16486 5607 16488 5616
rect 16540 5607 16542 5616
rect 16488 5578 16540 5584
rect 16488 4616 16540 4622
rect 16592 4604 16620 7686
rect 16684 7206 16712 8298
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 4758 16712 7142
rect 16776 5778 16804 9590
rect 16868 9110 16896 9658
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16960 8022 16988 11512
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 17130 10704 17186 10713
rect 17130 10639 17186 10648
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17052 9761 17080 9862
rect 17038 9752 17094 9761
rect 17038 9687 17094 9696
rect 17144 9178 17172 10639
rect 17236 9897 17264 11018
rect 17222 9888 17278 9897
rect 17222 9823 17278 9832
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17038 9072 17094 9081
rect 17038 9007 17094 9016
rect 17052 8634 17080 9007
rect 17236 8974 17264 9823
rect 17328 9654 17356 15830
rect 17512 14793 17540 20896
rect 17604 17338 17632 23151
rect 17684 23112 17736 23118
rect 17682 23080 17684 23089
rect 17736 23080 17738 23089
rect 17682 23015 17738 23024
rect 17696 22710 17724 23015
rect 17684 22704 17736 22710
rect 17684 22646 17736 22652
rect 17788 22166 17816 25928
rect 17868 25910 17920 25916
rect 18156 24834 18184 27520
rect 18708 25770 18736 27520
rect 18880 26104 18932 26110
rect 18880 26046 18932 26052
rect 18696 25764 18748 25770
rect 18696 25706 18748 25712
rect 18788 25764 18840 25770
rect 18788 25706 18840 25712
rect 18800 25498 18828 25706
rect 18788 25492 18840 25498
rect 18788 25434 18840 25440
rect 18512 25356 18564 25362
rect 18512 25298 18564 25304
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 17972 24806 18184 24834
rect 17868 24676 17920 24682
rect 17868 24618 17920 24624
rect 17880 23338 17908 24618
rect 17972 23633 18000 24806
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 18064 24206 18092 24686
rect 18248 24206 18276 25094
rect 18524 24614 18552 25298
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18340 24342 18368 24550
rect 18328 24336 18380 24342
rect 18326 24304 18328 24313
rect 18380 24304 18382 24313
rect 18326 24239 18382 24248
rect 18052 24200 18104 24206
rect 18236 24200 18288 24206
rect 18052 24142 18104 24148
rect 18142 24168 18198 24177
rect 18236 24142 18288 24148
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 18142 24103 18198 24112
rect 18156 23866 18184 24103
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 17958 23624 18014 23633
rect 17958 23559 18014 23568
rect 18144 23588 18196 23594
rect 18144 23530 18196 23536
rect 17880 23310 18000 23338
rect 18156 23322 18184 23530
rect 17972 23254 18000 23310
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 17960 23248 18012 23254
rect 17960 23190 18012 23196
rect 18156 23066 18184 23258
rect 17972 23038 18184 23066
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 17776 22160 17828 22166
rect 17776 22102 17828 22108
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17696 20602 17724 21966
rect 17880 21690 17908 22374
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17866 20632 17922 20641
rect 17684 20596 17736 20602
rect 17866 20567 17868 20576
rect 17684 20538 17736 20544
rect 17920 20567 17922 20576
rect 17868 20538 17920 20544
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17590 17096 17646 17105
rect 17590 17031 17646 17040
rect 17604 15638 17632 17031
rect 17788 16998 17816 18702
rect 17880 17814 17908 19790
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 17880 17270 17908 17750
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17866 16144 17922 16153
rect 17866 16079 17922 16088
rect 17880 15706 17908 16079
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17592 15632 17644 15638
rect 17880 15586 17908 15642
rect 17592 15574 17644 15580
rect 17604 15162 17632 15574
rect 17788 15558 17908 15586
rect 17788 15162 17816 15558
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17880 14906 17908 15302
rect 17972 15026 18000 23038
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 18064 22098 18092 22918
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 18156 21554 18184 22918
rect 18248 22681 18276 24006
rect 18432 23730 18460 24142
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 18234 22672 18290 22681
rect 18234 22607 18290 22616
rect 18236 22500 18288 22506
rect 18236 22442 18288 22448
rect 18248 22234 18276 22442
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18248 21486 18276 22170
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18050 19272 18106 19281
rect 18050 19207 18106 19216
rect 18064 17882 18092 19207
rect 18156 18970 18184 20538
rect 18340 19854 18368 23598
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18340 19242 18368 19654
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18144 18964 18196 18970
rect 18196 18924 18276 18952
rect 18144 18906 18196 18912
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18064 16726 18092 17818
rect 18156 17785 18184 18294
rect 18248 18222 18276 18924
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18142 17776 18198 17785
rect 18142 17711 18198 17720
rect 18248 17377 18276 18158
rect 18234 17368 18290 17377
rect 18234 17303 18290 17312
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18142 16144 18198 16153
rect 18142 16079 18198 16088
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17880 14878 18000 14906
rect 17498 14784 17554 14793
rect 17498 14719 17554 14728
rect 17866 14784 17922 14793
rect 17866 14719 17922 14728
rect 17880 14550 17908 14719
rect 17972 14618 18000 14878
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 18064 14346 18092 15438
rect 18156 15337 18184 16079
rect 18142 15328 18198 15337
rect 18142 15263 18198 15272
rect 18248 14414 18276 16934
rect 18432 16794 18460 23666
rect 18524 23186 18552 24550
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 18696 24132 18748 24138
rect 18696 24074 18748 24080
rect 18602 23624 18658 23633
rect 18602 23559 18604 23568
rect 18656 23559 18658 23568
rect 18604 23530 18656 23536
rect 18602 23488 18658 23497
rect 18602 23423 18658 23432
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18524 22273 18552 23122
rect 18510 22264 18566 22273
rect 18510 22199 18566 22208
rect 18512 20800 18564 20806
rect 18510 20768 18512 20777
rect 18564 20768 18566 20777
rect 18510 20703 18566 20712
rect 18616 20534 18644 23423
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18602 18864 18658 18873
rect 18512 18828 18564 18834
rect 18602 18799 18658 18808
rect 18512 18770 18564 18776
rect 18524 18601 18552 18770
rect 18510 18592 18566 18601
rect 18510 18527 18566 18536
rect 18524 17882 18552 18527
rect 18616 18290 18644 18799
rect 18708 18358 18736 24074
rect 18800 23730 18828 24346
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18892 23338 18920 26046
rect 18970 25528 19026 25537
rect 18970 25463 19026 25472
rect 18984 23866 19012 25463
rect 19062 24712 19118 24721
rect 19062 24647 19118 24656
rect 19076 24614 19104 24647
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 19260 24449 19288 27520
rect 19432 26648 19484 26654
rect 19432 26590 19484 26596
rect 19338 26208 19394 26217
rect 19338 26143 19394 26152
rect 19246 24440 19302 24449
rect 19246 24375 19302 24384
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 18972 23860 19024 23866
rect 18972 23802 19024 23808
rect 18984 23662 19012 23802
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 18800 23310 18920 23338
rect 18800 22030 18828 23310
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 18972 23248 19024 23254
rect 19076 23236 19104 23734
rect 19168 23361 19196 24006
rect 19154 23352 19210 23361
rect 19352 23322 19380 26143
rect 19444 25158 19472 26590
rect 19812 26042 19840 27520
rect 19800 26036 19852 26042
rect 19800 25978 19852 25984
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19432 24608 19484 24614
rect 19536 24596 19564 25298
rect 20076 25152 20128 25158
rect 20076 25094 20128 25100
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 19484 24568 19564 24596
rect 19432 24550 19484 24556
rect 19154 23287 19210 23296
rect 19340 23316 19392 23322
rect 19024 23208 19104 23236
rect 18972 23190 19024 23196
rect 18892 22166 18920 23190
rect 18880 22160 18932 22166
rect 18880 22102 18932 22108
rect 18984 22098 19012 23190
rect 19168 22273 19196 23287
rect 19340 23258 19392 23264
rect 19444 23202 19472 24550
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19996 24410 20024 24890
rect 20088 24750 20116 25094
rect 20166 24984 20222 24993
rect 20166 24919 20222 24928
rect 20076 24744 20128 24750
rect 20076 24686 20128 24692
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19708 24268 19760 24274
rect 19708 24210 19760 24216
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19352 23174 19472 23202
rect 19352 23089 19380 23174
rect 19338 23080 19394 23089
rect 19338 23015 19394 23024
rect 19340 22976 19392 22982
rect 19338 22944 19340 22953
rect 19432 22976 19484 22982
rect 19392 22944 19394 22953
rect 19432 22918 19484 22924
rect 19338 22879 19394 22888
rect 19340 22704 19392 22710
rect 19338 22672 19340 22681
rect 19392 22672 19394 22681
rect 19338 22607 19394 22616
rect 19340 22568 19392 22574
rect 19338 22536 19340 22545
rect 19392 22536 19394 22545
rect 19338 22471 19394 22480
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19154 22264 19210 22273
rect 19154 22199 19210 22208
rect 18972 22092 19024 22098
rect 18972 22034 19024 22040
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18972 21072 19024 21078
rect 18972 21014 19024 21020
rect 18788 20868 18840 20874
rect 18788 20810 18840 20816
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18616 17649 18644 18226
rect 18800 18086 18828 20810
rect 18984 20641 19012 21014
rect 19064 20936 19116 20942
rect 19064 20878 19116 20884
rect 18970 20632 19026 20641
rect 19076 20602 19104 20878
rect 18970 20567 19026 20576
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 18880 20528 18932 20534
rect 19168 20482 19196 22034
rect 19352 21486 19380 22374
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19444 21321 19472 22918
rect 19536 22030 19564 24006
rect 19720 23866 19748 24210
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19984 23520 20036 23526
rect 20088 23497 20116 24550
rect 19984 23462 20036 23468
rect 20074 23488 20130 23497
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19800 23044 19852 23050
rect 19800 22986 19852 22992
rect 19812 22710 19840 22986
rect 19996 22982 20024 23462
rect 20074 23423 20130 23432
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19708 22704 19760 22710
rect 19706 22672 19708 22681
rect 19800 22704 19852 22710
rect 19760 22672 19762 22681
rect 19800 22646 19852 22652
rect 19706 22607 19762 22616
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19616 22160 19668 22166
rect 19614 22128 19616 22137
rect 19668 22128 19670 22137
rect 19614 22063 19670 22072
rect 19524 22024 19576 22030
rect 19524 21966 19576 21972
rect 19430 21312 19486 21321
rect 19430 21247 19486 21256
rect 19260 21010 19472 21026
rect 19248 21004 19472 21010
rect 19300 20998 19472 21004
rect 19248 20946 19300 20952
rect 19338 20904 19394 20913
rect 19338 20839 19394 20848
rect 18880 20470 18932 20476
rect 18892 19417 18920 20470
rect 19076 20454 19196 20482
rect 19248 20460 19300 20466
rect 18878 19408 18934 19417
rect 18878 19343 18934 19352
rect 18970 19000 19026 19009
rect 18970 18935 19026 18944
rect 18984 18902 19012 18935
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18984 18426 19012 18838
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18694 17912 18750 17921
rect 18694 17847 18750 17856
rect 18602 17640 18658 17649
rect 18602 17575 18658 17584
rect 18708 17218 18736 17847
rect 18800 17513 18828 18022
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18786 17504 18842 17513
rect 18786 17439 18842 17448
rect 18892 17354 18920 17614
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18616 17190 18736 17218
rect 18800 17326 18920 17354
rect 18800 17202 18828 17326
rect 18788 17196 18840 17202
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18340 16046 18368 16594
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18432 15910 18460 16730
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18432 15706 18460 15846
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18512 15496 18564 15502
rect 18326 15464 18382 15473
rect 18512 15438 18564 15444
rect 18326 15399 18382 15408
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18248 14249 18276 14350
rect 18234 14240 18290 14249
rect 18234 14175 18290 14184
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17512 12986 17540 13330
rect 18340 13274 18368 15399
rect 18524 15094 18552 15438
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18432 13938 18460 14350
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18524 13870 18552 14010
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18524 13394 18552 13806
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18340 13246 18552 13274
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 18340 12850 18368 13126
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17788 11257 17816 12038
rect 17774 11248 17830 11257
rect 17774 11183 17830 11192
rect 17880 10674 17908 12718
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 18064 12306 18092 12650
rect 18432 12374 18460 12854
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17774 10568 17830 10577
rect 17774 10503 17830 10512
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17420 9897 17448 9998
rect 17406 9888 17462 9897
rect 17406 9823 17462 9832
rect 17316 9648 17368 9654
rect 17512 9625 17540 10134
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17604 9722 17632 9998
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17788 9654 17816 10503
rect 17960 10192 18012 10198
rect 17958 10160 17960 10169
rect 18012 10160 18014 10169
rect 17958 10095 18014 10104
rect 17776 9648 17828 9654
rect 17316 9590 17368 9596
rect 17498 9616 17554 9625
rect 17776 9590 17828 9596
rect 17498 9551 17554 9560
rect 17314 9344 17370 9353
rect 17314 9279 17370 9288
rect 17328 9081 17356 9279
rect 17314 9072 17370 9081
rect 17314 9007 17370 9016
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17592 8832 17644 8838
rect 17512 8792 17592 8820
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17408 8560 17460 8566
rect 17406 8528 17408 8537
rect 17460 8528 17462 8537
rect 17406 8463 17462 8472
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16868 7426 16896 7754
rect 16960 7546 16988 7958
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17420 7449 17448 7686
rect 17406 7440 17462 7449
rect 16868 7398 16988 7426
rect 16960 7313 16988 7398
rect 17406 7375 17462 7384
rect 16946 7304 17002 7313
rect 16946 7239 17002 7248
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16868 6322 16896 6870
rect 16960 6662 16988 7239
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16960 6458 16988 6598
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 17052 5846 17080 6326
rect 17222 5944 17278 5953
rect 17222 5879 17278 5888
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16776 5098 16804 5714
rect 16764 5092 16816 5098
rect 16764 5034 16816 5040
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16540 4576 16620 4604
rect 16488 4558 16540 4564
rect 16394 4312 16450 4321
rect 16394 4247 16450 4256
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16316 3126 16344 4014
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16488 3392 16540 3398
rect 16486 3360 16488 3369
rect 16540 3360 16542 3369
rect 16486 3295 16542 3304
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16592 2553 16620 3402
rect 16670 2680 16726 2689
rect 16670 2615 16726 2624
rect 16578 2544 16634 2553
rect 16684 2514 16712 2615
rect 16776 2582 16804 5034
rect 17052 4457 17080 5782
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17038 4448 17094 4457
rect 17038 4383 17094 4392
rect 17038 4312 17094 4321
rect 17038 4247 17094 4256
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16868 3233 16896 3538
rect 16854 3224 16910 3233
rect 16854 3159 16910 3168
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 16578 2479 16634 2488
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16408 598 16528 626
rect 16408 513 16436 598
rect 16394 504 16450 513
rect 15566 368 15622 377
rect 15566 303 15622 312
rect 16026 0 16082 480
rect 16500 480 16528 598
rect 17052 480 17080 4247
rect 17144 4185 17172 4558
rect 17130 4176 17186 4185
rect 17130 4111 17186 4120
rect 17130 3768 17186 3777
rect 17130 3703 17132 3712
rect 17184 3703 17186 3712
rect 17132 3674 17184 3680
rect 17236 3670 17264 5879
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17328 5137 17356 5510
rect 17314 5128 17370 5137
rect 17314 5063 17370 5072
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17328 4185 17356 4966
rect 17420 4826 17448 5782
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17420 4282 17448 4762
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17314 4176 17370 4185
rect 17314 4111 17370 4120
rect 17420 3738 17448 4218
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17236 3194 17264 3606
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17420 2145 17448 2246
rect 17406 2136 17462 2145
rect 17406 2071 17462 2080
rect 17512 1329 17540 8792
rect 18064 8820 18092 12242
rect 18326 11792 18382 11801
rect 18326 11727 18382 11736
rect 18340 10266 18368 11727
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18340 9042 18368 9318
rect 18432 9178 18460 12310
rect 18524 11801 18552 13246
rect 18616 11937 18644 17190
rect 18788 17138 18840 17144
rect 18800 16425 18828 17138
rect 18984 16810 19012 17478
rect 18892 16782 19012 16810
rect 18786 16416 18842 16425
rect 18786 16351 18842 16360
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18800 14958 18828 15914
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18800 14278 18828 14894
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18800 14074 18828 14214
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18892 12753 18920 16782
rect 19076 16153 19104 20454
rect 19352 20448 19380 20839
rect 19444 20482 19472 20998
rect 19536 20602 19564 21966
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19444 20454 19564 20482
rect 19300 20420 19380 20448
rect 19248 20402 19300 20408
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19168 16250 19196 19858
rect 19260 19786 19288 20402
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19352 19689 19380 20198
rect 19444 20058 19472 20266
rect 19536 20262 19564 20454
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19432 20052 19484 20058
rect 19536 20040 19564 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19536 20012 19656 20040
rect 19432 19994 19484 20000
rect 19338 19680 19394 19689
rect 19260 19638 19338 19666
rect 19260 18698 19288 19638
rect 19338 19615 19394 19624
rect 19444 19514 19472 19994
rect 19432 19508 19484 19514
rect 19484 19468 19564 19496
rect 19432 19450 19484 19456
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19062 16144 19118 16153
rect 19062 16079 19118 16088
rect 19260 15978 19288 16934
rect 19352 16017 19380 19314
rect 19432 19236 19484 19242
rect 19432 19178 19484 19184
rect 19444 18970 19472 19178
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19444 18426 19472 18906
rect 19536 18902 19564 19468
rect 19628 19378 19656 20012
rect 19996 19990 20024 21286
rect 20088 20466 20116 23258
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19984 19984 20036 19990
rect 19984 19926 20036 19932
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19996 18970 20024 19926
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 20088 19174 20116 19654
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20088 19009 20116 19110
rect 20074 19000 20130 19009
rect 19984 18964 20036 18970
rect 20074 18935 20130 18944
rect 19984 18906 20036 18912
rect 19524 18896 19576 18902
rect 20076 18896 20128 18902
rect 19524 18838 19576 18844
rect 19614 18864 19670 18873
rect 20076 18838 20128 18844
rect 19614 18799 19670 18808
rect 19628 18748 19656 18799
rect 19536 18720 19656 18748
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19444 17746 19472 18362
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19444 16794 19472 17682
rect 19536 17377 19564 18720
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19996 18034 20024 18566
rect 20088 18222 20116 18838
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19996 18006 20116 18034
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19800 17808 19852 17814
rect 19800 17750 19852 17756
rect 19616 17604 19668 17610
rect 19616 17546 19668 17552
rect 19522 17368 19578 17377
rect 19522 17303 19578 17312
rect 19628 17202 19656 17546
rect 19812 17338 19840 17750
rect 19890 17368 19946 17377
rect 19800 17332 19852 17338
rect 19890 17303 19946 17312
rect 19800 17274 19852 17280
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19536 16522 19564 17138
rect 19904 17134 19932 17303
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19996 16658 20024 16934
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19522 16416 19578 16425
rect 19522 16351 19578 16360
rect 19338 16008 19394 16017
rect 19248 15972 19300 15978
rect 19338 15943 19394 15952
rect 19248 15914 19300 15920
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19062 15600 19118 15609
rect 19062 15535 19118 15544
rect 18972 15360 19024 15366
rect 18970 15328 18972 15337
rect 19024 15328 19026 15337
rect 18970 15263 19026 15272
rect 19076 15162 19104 15535
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 19260 14618 19288 15370
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 18984 13802 19012 14282
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 18984 13462 19012 13738
rect 19062 13696 19118 13705
rect 19062 13631 19118 13640
rect 18972 13456 19024 13462
rect 18972 13398 19024 13404
rect 18878 12744 18934 12753
rect 18878 12679 18934 12688
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18984 12442 19012 12582
rect 18972 12436 19024 12442
rect 18892 12396 18972 12424
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18602 11928 18658 11937
rect 18602 11863 18658 11872
rect 18510 11792 18566 11801
rect 18510 11727 18566 11736
rect 18512 11144 18564 11150
rect 18616 11132 18644 11863
rect 18708 11694 18736 12242
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18708 11286 18736 11630
rect 18696 11280 18748 11286
rect 18696 11222 18748 11228
rect 18616 11104 18736 11132
rect 18512 11086 18564 11092
rect 18524 10810 18552 11086
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18602 10568 18658 10577
rect 18602 10503 18658 10512
rect 18616 9994 18644 10503
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 17592 8774 17644 8780
rect 17696 8792 18092 8820
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7206 17632 7822
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17604 6866 17632 7142
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17604 6633 17632 6802
rect 17590 6624 17646 6633
rect 17590 6559 17646 6568
rect 17604 6254 17632 6559
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17604 5914 17632 6190
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17590 5536 17646 5545
rect 17590 5471 17646 5480
rect 17498 1320 17554 1329
rect 17498 1255 17554 1264
rect 17604 480 17632 5471
rect 17696 5370 17724 8792
rect 18340 8430 18368 8978
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18340 8294 18368 8366
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17788 6866 17816 7210
rect 17880 7206 17908 7890
rect 18234 7576 18290 7585
rect 18234 7511 18236 7520
rect 18288 7511 18290 7520
rect 18236 7482 18288 7488
rect 18340 7478 18368 8230
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 18340 7274 18368 7414
rect 18432 7313 18460 7822
rect 18512 7744 18564 7750
rect 18616 7721 18644 7958
rect 18512 7686 18564 7692
rect 18602 7712 18658 7721
rect 18418 7304 18474 7313
rect 18328 7268 18380 7274
rect 18524 7290 18552 7686
rect 18602 7647 18658 7656
rect 18616 7449 18644 7647
rect 18708 7546 18736 11104
rect 18800 9489 18828 11766
rect 18892 11744 18920 12396
rect 18972 12378 19024 12384
rect 18970 12200 19026 12209
rect 18970 12135 18972 12144
rect 19024 12135 19026 12144
rect 18972 12106 19024 12112
rect 19076 11762 19104 13631
rect 19246 13560 19302 13569
rect 19246 13495 19302 13504
rect 19260 13394 19288 13495
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19352 13274 19380 15846
rect 19432 15632 19484 15638
rect 19430 15600 19432 15609
rect 19484 15600 19486 15609
rect 19430 15535 19486 15544
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19444 14618 19472 14826
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19430 14512 19486 14521
rect 19430 14447 19486 14456
rect 19444 13530 19472 14447
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19260 13246 19380 13274
rect 19156 12912 19208 12918
rect 19154 12880 19156 12889
rect 19208 12880 19210 12889
rect 19260 12850 19288 13246
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 12889 19380 13126
rect 19444 12986 19472 13330
rect 19536 12986 19564 16351
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19996 15688 20024 16594
rect 20088 16289 20116 18006
rect 20074 16280 20130 16289
rect 20074 16215 20130 16224
rect 20088 15745 20116 16215
rect 19904 15660 20024 15688
rect 20074 15736 20130 15745
rect 20074 15671 20130 15680
rect 19904 14890 19932 15660
rect 19982 15056 20038 15065
rect 19982 14991 20038 15000
rect 19892 14884 19944 14890
rect 19892 14826 19944 14832
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14618 20024 14991
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19720 14074 19748 14418
rect 19982 14376 20038 14385
rect 19982 14311 20038 14320
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19720 13841 19748 14010
rect 19706 13832 19762 13841
rect 19706 13767 19762 13776
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19996 13308 20024 14311
rect 20088 13569 20116 14758
rect 20180 14482 20208 24919
rect 20260 24880 20312 24886
rect 20260 24822 20312 24828
rect 20272 24410 20300 24822
rect 20260 24404 20312 24410
rect 20260 24346 20312 24352
rect 20364 23712 20392 27520
rect 20812 26580 20864 26586
rect 20812 26522 20864 26528
rect 20444 26308 20496 26314
rect 20444 26250 20496 26256
rect 20272 23684 20392 23712
rect 20272 23225 20300 23684
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20364 23322 20392 23530
rect 20352 23316 20404 23322
rect 20352 23258 20404 23264
rect 20258 23216 20314 23225
rect 20258 23151 20314 23160
rect 20364 23050 20392 23258
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 20456 22794 20484 26250
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20640 24682 20668 25094
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 20534 23896 20590 23905
rect 20534 23831 20590 23840
rect 20548 22982 20576 23831
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20272 22766 20484 22794
rect 20272 14618 20300 22766
rect 20548 22574 20576 22918
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20444 22500 20496 22506
rect 20444 22442 20496 22448
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20364 21350 20392 21830
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20364 21146 20392 21286
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20364 20398 20392 20742
rect 20352 20392 20404 20398
rect 20350 20360 20352 20369
rect 20404 20360 20406 20369
rect 20350 20295 20406 20304
rect 20364 20269 20392 20295
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20364 18630 20392 19790
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20456 17746 20484 22442
rect 20536 21072 20588 21078
rect 20536 21014 20588 21020
rect 20548 19281 20576 21014
rect 20534 19272 20590 19281
rect 20534 19207 20590 19216
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20444 17740 20496 17746
rect 20444 17682 20496 17688
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20364 15706 20392 17138
rect 20456 16726 20484 17682
rect 20548 17542 20576 18838
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20548 17105 20576 17206
rect 20534 17096 20590 17105
rect 20534 17031 20590 17040
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20548 16794 20576 16934
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20456 15978 20484 16526
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20456 15026 20484 15506
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20444 14476 20496 14482
rect 20444 14418 20496 14424
rect 20166 14104 20222 14113
rect 20166 14039 20222 14048
rect 20350 14104 20406 14113
rect 20350 14039 20406 14048
rect 20180 13841 20208 14039
rect 20166 13832 20222 13841
rect 20166 13767 20222 13776
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20074 13560 20130 13569
rect 20074 13495 20130 13504
rect 20088 13462 20116 13495
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 19996 13280 20116 13308
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19338 12880 19394 12889
rect 19154 12815 19210 12824
rect 19248 12844 19300 12850
rect 19338 12815 19394 12824
rect 19798 12880 19854 12889
rect 19798 12815 19854 12824
rect 19248 12786 19300 12792
rect 19260 12730 19288 12786
rect 19260 12702 19472 12730
rect 19812 12714 19840 12815
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 12481 19380 12582
rect 19338 12472 19394 12481
rect 19338 12407 19394 12416
rect 19156 12232 19208 12238
rect 19154 12200 19156 12209
rect 19208 12200 19210 12209
rect 19154 12135 19210 12144
rect 19064 11756 19116 11762
rect 18892 11716 19012 11744
rect 18878 11656 18934 11665
rect 18878 11591 18880 11600
rect 18932 11591 18934 11600
rect 18880 11562 18932 11568
rect 18984 11257 19012 11716
rect 19064 11698 19116 11704
rect 19076 11354 19104 11698
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18970 11248 19026 11257
rect 18970 11183 19026 11192
rect 19168 11082 19196 12135
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 18972 10532 19024 10538
rect 18972 10474 19024 10480
rect 18786 9480 18842 9489
rect 18786 9415 18842 9424
rect 18800 9178 18828 9415
rect 18984 9382 19012 10474
rect 19076 10198 19104 10746
rect 19260 10470 19288 12038
rect 19444 11898 19472 12702
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19444 11694 19472 11834
rect 20088 11830 20116 13280
rect 20180 13190 20208 13670
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20180 12850 20208 13126
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20260 12368 20312 12374
rect 20258 12336 20260 12345
rect 20312 12336 20314 12345
rect 20258 12271 20314 12280
rect 20258 11928 20314 11937
rect 20258 11863 20314 11872
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19340 11552 19392 11558
rect 19338 11520 19340 11529
rect 19392 11520 19394 11529
rect 19338 11455 19394 11464
rect 19444 11218 19472 11630
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19708 11280 19760 11286
rect 19628 11228 19708 11234
rect 19628 11222 19760 11228
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19628 11206 19748 11222
rect 19340 10736 19392 10742
rect 19338 10704 19340 10713
rect 19444 10724 19472 11154
rect 19628 10742 19656 11206
rect 19616 10736 19668 10742
rect 19392 10704 19394 10713
rect 19444 10696 19564 10724
rect 19338 10639 19394 10648
rect 19248 10464 19300 10470
rect 19300 10412 19472 10418
rect 19248 10406 19472 10412
rect 19260 10390 19472 10406
rect 19064 10192 19116 10198
rect 19062 10160 19064 10169
rect 19116 10160 19118 10169
rect 19062 10095 19118 10104
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19168 9722 19196 9998
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19156 9716 19208 9722
rect 19076 9676 19156 9704
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18984 9178 19012 9318
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18800 8537 18828 8978
rect 18984 8634 19012 9114
rect 19076 8634 19104 9676
rect 19156 9658 19208 9664
rect 19260 8838 19288 9930
rect 19248 8832 19300 8838
rect 19300 8792 19380 8820
rect 19248 8774 19300 8780
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 18786 8528 18842 8537
rect 18786 8463 18842 8472
rect 18984 8430 19012 8570
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18984 8090 19012 8366
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18602 7440 18658 7449
rect 18602 7375 18658 7384
rect 18708 7342 18736 7482
rect 18696 7336 18748 7342
rect 18524 7262 18644 7290
rect 18696 7278 18748 7284
rect 19076 7274 19104 8570
rect 19248 8424 19300 8430
rect 19246 8392 19248 8401
rect 19300 8392 19302 8401
rect 19246 8327 19302 8336
rect 19246 8120 19302 8129
rect 19352 8090 19380 8792
rect 19444 8090 19472 10390
rect 19536 10266 19564 10696
rect 19616 10678 19668 10684
rect 19996 10606 20024 11766
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 20180 11132 20208 11494
rect 20272 11257 20300 11863
rect 20364 11626 20392 14039
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20258 11248 20314 11257
rect 20258 11183 20314 11192
rect 20352 11144 20404 11150
rect 20074 11112 20130 11121
rect 20180 11104 20300 11132
rect 20074 11047 20130 11056
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 20088 10538 20116 11047
rect 20168 10736 20220 10742
rect 20168 10678 20220 10684
rect 20076 10532 20128 10538
rect 20076 10474 20128 10480
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 20088 10198 20116 10474
rect 20076 10192 20128 10198
rect 20076 10134 20128 10140
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19536 9178 19564 9454
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19246 8055 19302 8064
rect 19340 8084 19392 8090
rect 19260 7970 19288 8055
rect 19340 8026 19392 8032
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19260 7942 19380 7970
rect 19352 7721 19380 7942
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19338 7712 19394 7721
rect 19338 7647 19394 7656
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 18418 7239 18474 7248
rect 18328 7210 18380 7216
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17788 6118 17816 6802
rect 17880 6662 17908 7142
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17788 5545 17816 6054
rect 17880 5846 17908 6598
rect 18510 6488 18566 6497
rect 18510 6423 18512 6432
rect 18564 6423 18566 6432
rect 18512 6394 18564 6400
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 18156 5846 18184 6326
rect 18616 6118 18644 7262
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 19076 6866 19104 7210
rect 19260 7177 19288 7278
rect 19246 7168 19302 7177
rect 19246 7103 19302 7112
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 6322 18736 6598
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18696 6180 18748 6186
rect 18696 6122 18748 6128
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 17868 5840 17920 5846
rect 18144 5840 18196 5846
rect 17868 5782 17920 5788
rect 18050 5808 18106 5817
rect 17960 5772 18012 5778
rect 18616 5817 18644 6054
rect 18708 5914 18736 6122
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18144 5782 18196 5788
rect 18602 5808 18658 5817
rect 18050 5743 18106 5752
rect 18602 5743 18658 5752
rect 17960 5714 18012 5720
rect 17774 5536 17830 5545
rect 17774 5471 17830 5480
rect 17972 5386 18000 5714
rect 17880 5370 18000 5386
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17868 5364 18000 5370
rect 17920 5358 18000 5364
rect 17868 5306 17920 5312
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17682 3904 17738 3913
rect 17682 3839 17738 3848
rect 17696 3194 17724 3839
rect 17788 3466 17816 5170
rect 17868 4480 17920 4486
rect 17920 4440 18000 4468
rect 17868 4422 17920 4428
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17880 1329 17908 3878
rect 17972 3058 18000 4440
rect 18064 3074 18092 5743
rect 18604 5704 18656 5710
rect 18418 5672 18474 5681
rect 18418 5607 18474 5616
rect 18602 5672 18604 5681
rect 18656 5672 18658 5681
rect 18602 5607 18658 5616
rect 18326 5536 18382 5545
rect 18326 5471 18382 5480
rect 18340 5302 18368 5471
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 18340 4690 18368 5238
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18156 4010 18184 4626
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18248 3942 18276 3973
rect 18236 3936 18288 3942
rect 18234 3904 18236 3913
rect 18288 3904 18290 3913
rect 18234 3839 18290 3848
rect 18248 3670 18276 3839
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18432 3505 18460 5607
rect 18510 5536 18566 5545
rect 18510 5471 18566 5480
rect 18524 5234 18552 5471
rect 18616 5370 18644 5607
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18708 5234 18736 5850
rect 18972 5840 19024 5846
rect 18972 5782 19024 5788
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18602 5128 18658 5137
rect 18602 5063 18604 5072
rect 18656 5063 18658 5072
rect 18604 5034 18656 5040
rect 18708 4758 18736 5170
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18708 3942 18736 4694
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18708 3738 18736 3878
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18142 3496 18198 3505
rect 18142 3431 18198 3440
rect 18418 3496 18474 3505
rect 18418 3431 18474 3440
rect 18156 3194 18184 3431
rect 18602 3360 18658 3369
rect 18602 3295 18658 3304
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 17960 3052 18012 3058
rect 18064 3046 18184 3074
rect 17960 2994 18012 3000
rect 17866 1320 17922 1329
rect 17866 1255 17922 1264
rect 18156 480 18184 3046
rect 18616 2922 18644 3295
rect 18694 3224 18750 3233
rect 18694 3159 18750 3168
rect 18708 3058 18736 3159
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 18708 2825 18736 2858
rect 18694 2816 18750 2825
rect 18694 2751 18750 2760
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 18892 2417 18920 2518
rect 18878 2408 18934 2417
rect 18878 2343 18934 2352
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18432 1873 18460 2246
rect 18604 2032 18656 2038
rect 18604 1974 18656 1980
rect 18418 1864 18474 1873
rect 18418 1799 18474 1808
rect 18616 480 18644 1974
rect 18984 1873 19012 5782
rect 19352 5778 19380 7647
rect 19444 6798 19472 7890
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19800 6928 19852 6934
rect 19800 6870 19852 6876
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19536 6458 19564 6802
rect 19812 6769 19840 6870
rect 19798 6760 19854 6769
rect 19798 6695 19854 6704
rect 19982 6760 20038 6769
rect 19982 6695 20038 6704
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19720 6225 19748 6326
rect 19706 6216 19762 6225
rect 19706 6151 19762 6160
rect 19812 6100 19840 6695
rect 19996 6361 20024 6695
rect 19982 6352 20038 6361
rect 19982 6287 20038 6296
rect 19996 6254 20024 6287
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19812 6072 20024 6100
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19260 5250 19288 5578
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19338 5264 19394 5273
rect 19260 5222 19338 5250
rect 19338 5199 19394 5208
rect 19430 4856 19486 4865
rect 19430 4791 19486 4800
rect 19444 4622 19472 4791
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19430 3768 19486 3777
rect 19430 3703 19432 3712
rect 19484 3703 19486 3712
rect 19432 3674 19484 3680
rect 19338 3632 19394 3641
rect 19338 3567 19394 3576
rect 19352 3466 19380 3567
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 19076 2990 19104 3334
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19076 2446 19104 2926
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19154 2272 19210 2281
rect 19154 2207 19210 2216
rect 18970 1864 19026 1873
rect 18970 1799 19026 1808
rect 19168 480 19196 2207
rect 19352 1465 19380 3062
rect 19536 2650 19564 5510
rect 19720 5370 19748 5714
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19996 5030 20024 6072
rect 20088 5778 20116 9590
rect 20180 8537 20208 10678
rect 20272 10033 20300 11104
rect 20352 11086 20404 11092
rect 20258 10024 20314 10033
rect 20258 9959 20314 9968
rect 20364 9908 20392 11086
rect 20272 9880 20392 9908
rect 20272 9489 20300 9880
rect 20258 9480 20314 9489
rect 20258 9415 20314 9424
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20364 9178 20392 9386
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20166 8528 20222 8537
rect 20166 8463 20222 8472
rect 20350 7712 20406 7721
rect 20350 7647 20406 7656
rect 20364 7410 20392 7647
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20272 6662 20300 7142
rect 20350 7032 20406 7041
rect 20350 6967 20406 6976
rect 20364 6934 20392 6967
rect 20352 6928 20404 6934
rect 20352 6870 20404 6876
rect 20456 6866 20484 14418
rect 20548 13258 20576 16458
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20536 12640 20588 12646
rect 20534 12608 20536 12617
rect 20588 12608 20590 12617
rect 20534 12543 20590 12552
rect 20640 12458 20668 24618
rect 20720 24064 20772 24070
rect 20720 24006 20772 24012
rect 20732 23322 20760 24006
rect 20824 23905 20852 26522
rect 20916 25498 20944 27520
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 21088 24336 21140 24342
rect 20902 24304 20958 24313
rect 21088 24278 21140 24284
rect 20902 24239 20958 24248
rect 20810 23896 20866 23905
rect 20810 23831 20866 23840
rect 20812 23792 20864 23798
rect 20812 23734 20864 23740
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20718 23216 20774 23225
rect 20718 23151 20774 23160
rect 20732 22522 20760 23151
rect 20824 23089 20852 23734
rect 20810 23080 20866 23089
rect 20810 23015 20866 23024
rect 20732 22494 20852 22522
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20732 22098 20760 22374
rect 20824 22234 20852 22494
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20916 22148 20944 24239
rect 21100 23526 21128 24278
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 21100 23361 21128 23462
rect 21086 23352 21142 23361
rect 21086 23287 21142 23296
rect 21192 23066 21220 27639
rect 21546 27520 21602 28000
rect 22098 27520 22154 28000
rect 22650 27520 22706 28000
rect 23202 27520 23258 28000
rect 23754 27520 23810 28000
rect 24306 27520 24362 28000
rect 24858 27520 24914 28000
rect 25410 27520 25466 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 21560 26178 21588 27520
rect 21548 26172 21600 26178
rect 21548 26114 21600 26120
rect 22112 25702 22140 27520
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 22466 25392 22522 25401
rect 21272 25356 21324 25362
rect 22466 25327 22522 25336
rect 21272 25298 21324 25304
rect 21284 24614 21312 25298
rect 22376 25220 22428 25226
rect 22376 25162 22428 25168
rect 21640 25152 21692 25158
rect 21640 25094 21692 25100
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21100 23038 21220 23066
rect 20996 22160 21048 22166
rect 20810 22128 20866 22137
rect 20720 22092 20772 22098
rect 20916 22120 20996 22148
rect 20996 22102 21048 22108
rect 21100 22098 21128 23038
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 20810 22063 20866 22072
rect 21088 22092 21140 22098
rect 20720 22034 20772 22040
rect 20732 21865 20760 22034
rect 20718 21856 20774 21865
rect 20718 21791 20774 21800
rect 20718 20632 20774 20641
rect 20718 20567 20774 20576
rect 20732 17542 20760 20567
rect 20824 17814 20852 22063
rect 21088 22034 21140 22040
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20916 21418 20944 21966
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 20904 21412 20956 21418
rect 20904 21354 20956 21360
rect 20916 20602 20944 21354
rect 21100 21078 21128 21898
rect 21088 21072 21140 21078
rect 20994 21040 21050 21049
rect 21088 21014 21140 21020
rect 20994 20975 21050 20984
rect 21008 20874 21036 20975
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20916 20369 20944 20402
rect 20902 20360 20958 20369
rect 20902 20295 20958 20304
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20916 19922 20944 20198
rect 20994 20088 21050 20097
rect 20994 20023 21050 20032
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20916 18766 20944 19654
rect 21008 19530 21036 20023
rect 21100 19718 21128 20878
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21086 19544 21142 19553
rect 21008 19502 21086 19530
rect 21086 19479 21142 19488
rect 20994 19136 21050 19145
rect 20994 19071 21050 19080
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20916 18272 20944 18702
rect 21008 18698 21036 19071
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20916 18244 21036 18272
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20916 17882 20944 18090
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20732 15473 20760 17274
rect 20718 15464 20774 15473
rect 20718 15399 20774 15408
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20732 14618 20760 15098
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20718 14512 20774 14521
rect 20718 14447 20720 14456
rect 20772 14447 20774 14456
rect 20720 14418 20772 14424
rect 20718 14240 20774 14249
rect 20718 14175 20774 14184
rect 20732 12986 20760 14175
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20548 12430 20668 12458
rect 20548 9722 20576 12430
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 11626 20668 12038
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20732 11354 20760 12174
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20640 10554 20668 11222
rect 20640 10538 20760 10554
rect 20640 10532 20772 10538
rect 20640 10526 20720 10532
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20640 9518 20668 10526
rect 20720 10474 20772 10480
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20732 9110 20760 10134
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20626 8392 20682 8401
rect 20626 8327 20682 8336
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20352 6724 20404 6730
rect 20352 6666 20404 6672
rect 20260 6656 20312 6662
rect 20258 6624 20260 6633
rect 20312 6624 20314 6633
rect 20258 6559 20314 6568
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 20076 5636 20128 5642
rect 20076 5578 20128 5584
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19904 2922 19932 3470
rect 19996 2990 20024 3878
rect 20088 3126 20116 5578
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20272 5166 20300 5510
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20272 4826 20300 5102
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20166 4040 20222 4049
rect 20166 3975 20168 3984
rect 20220 3975 20222 3984
rect 20168 3946 20220 3952
rect 20166 3632 20222 3641
rect 20166 3567 20222 3576
rect 20076 3120 20128 3126
rect 20076 3062 20128 3068
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 20088 2922 20116 3062
rect 20180 3058 20208 3567
rect 20258 3496 20314 3505
rect 20258 3431 20314 3440
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 20076 2916 20128 2922
rect 20076 2858 20128 2864
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2644 19576 2650
rect 19996 2632 20024 2790
rect 19524 2586 19576 2592
rect 19720 2604 20024 2632
rect 19338 1456 19394 1465
rect 19338 1391 19394 1400
rect 19720 480 19748 2604
rect 20076 2372 20128 2378
rect 20076 2314 20128 2320
rect 20088 1057 20116 2314
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 20180 1465 20208 2246
rect 20166 1456 20222 1465
rect 20166 1391 20222 1400
rect 20272 1306 20300 3431
rect 20364 3369 20392 6666
rect 20456 6458 20484 6802
rect 20640 6798 20668 8327
rect 20824 8090 20852 17274
rect 20916 10146 20944 17614
rect 21008 17270 21036 18244
rect 21100 18057 21128 19479
rect 21086 18048 21142 18057
rect 21086 17983 21142 17992
rect 21192 17678 21220 22918
rect 21284 22817 21312 24550
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 21364 23792 21416 23798
rect 21560 23769 21588 24006
rect 21364 23734 21416 23740
rect 21546 23760 21602 23769
rect 21376 23633 21404 23734
rect 21546 23695 21602 23704
rect 21652 23662 21680 25094
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22008 24676 22060 24682
rect 22008 24618 22060 24624
rect 21824 24608 21876 24614
rect 21744 24556 21824 24562
rect 21744 24550 21876 24556
rect 21744 24534 21864 24550
rect 21640 23656 21692 23662
rect 21362 23624 21418 23633
rect 21640 23598 21692 23604
rect 21362 23559 21418 23568
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21468 23225 21496 23258
rect 21454 23216 21510 23225
rect 21454 23151 21510 23160
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21270 22808 21326 22817
rect 21270 22743 21326 22752
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21284 22137 21312 22578
rect 21376 22506 21404 23054
rect 21560 22778 21588 23054
rect 21652 23050 21680 23598
rect 21640 23044 21692 23050
rect 21640 22986 21692 22992
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21454 22264 21510 22273
rect 21454 22199 21456 22208
rect 21508 22199 21510 22208
rect 21456 22170 21508 22176
rect 21270 22128 21326 22137
rect 21270 22063 21326 22072
rect 21270 21992 21326 22001
rect 21270 21927 21326 21936
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21100 17202 21128 17546
rect 21284 17338 21312 21927
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21560 21486 21588 21830
rect 21638 21720 21694 21729
rect 21638 21655 21694 21664
rect 21548 21480 21600 21486
rect 21468 21440 21548 21468
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21376 20262 21404 21082
rect 21364 20256 21416 20262
rect 21362 20224 21364 20233
rect 21416 20224 21418 20233
rect 21362 20159 21418 20168
rect 21468 19990 21496 21440
rect 21548 21422 21600 21428
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21560 21078 21588 21286
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21560 19990 21588 20538
rect 21456 19984 21508 19990
rect 21456 19926 21508 19932
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 21376 19514 21404 19858
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21468 19310 21496 19926
rect 21456 19304 21508 19310
rect 21376 19252 21456 19258
rect 21376 19246 21508 19252
rect 21376 19230 21496 19246
rect 21376 18601 21404 19230
rect 21560 18970 21588 19926
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 21456 18896 21508 18902
rect 21454 18864 21456 18873
rect 21508 18864 21510 18873
rect 21454 18799 21510 18808
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21362 18592 21418 18601
rect 21362 18527 21418 18536
rect 21376 18426 21404 18527
rect 21468 18465 21496 18702
rect 21454 18456 21510 18465
rect 21364 18420 21416 18426
rect 21454 18391 21456 18400
rect 21364 18362 21416 18368
rect 21508 18391 21510 18400
rect 21456 18362 21508 18368
rect 21468 18331 21496 18362
rect 21560 18154 21588 18906
rect 21548 18148 21600 18154
rect 21548 18090 21600 18096
rect 21546 18048 21602 18057
rect 21546 17983 21602 17992
rect 21560 17814 21588 17983
rect 21548 17808 21600 17814
rect 21376 17756 21548 17762
rect 21376 17750 21600 17756
rect 21376 17734 21588 17750
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 21008 16561 21036 16662
rect 20994 16552 21050 16561
rect 20994 16487 21050 16496
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 21008 15162 21036 15438
rect 21100 15162 21128 17138
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21192 16794 21220 17070
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21180 16652 21232 16658
rect 21232 16612 21312 16640
rect 21180 16594 21232 16600
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 16046 21220 16390
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21192 15706 21220 15982
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 21086 15056 21142 15065
rect 21086 14991 21142 15000
rect 20994 14784 21050 14793
rect 20994 14719 21050 14728
rect 21008 14346 21036 14719
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 21100 14074 21128 14991
rect 21192 14958 21220 15642
rect 21284 15638 21312 16612
rect 21272 15632 21324 15638
rect 21272 15574 21324 15580
rect 21284 15366 21312 15574
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 21178 13832 21234 13841
rect 21100 12442 21128 13806
rect 21178 13767 21234 13776
rect 21192 13462 21220 13767
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21192 12918 21220 13398
rect 21284 13308 21312 15302
rect 21376 15065 21404 17734
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21456 17128 21508 17134
rect 21454 17096 21456 17105
rect 21508 17096 21510 17105
rect 21454 17031 21510 17040
rect 21560 16998 21588 17614
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21560 16726 21588 16934
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 21652 16538 21680 21655
rect 21560 16510 21680 16538
rect 21456 15972 21508 15978
rect 21456 15914 21508 15920
rect 21468 15502 21496 15914
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21362 15056 21418 15065
rect 21362 14991 21418 15000
rect 21468 14822 21496 15438
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21376 14006 21404 14486
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21364 14000 21416 14006
rect 21362 13968 21364 13977
rect 21416 13968 21418 13977
rect 21362 13903 21418 13912
rect 21468 13530 21496 14010
rect 21560 13938 21588 16510
rect 21638 15056 21694 15065
rect 21638 14991 21640 15000
rect 21692 14991 21694 15000
rect 21640 14962 21692 14968
rect 21744 14618 21772 24534
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21836 23730 21864 24074
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21928 23322 21956 24142
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21836 21690 21864 23122
rect 21824 21684 21876 21690
rect 21824 21626 21876 21632
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21836 20913 21864 21490
rect 21822 20904 21878 20913
rect 21822 20839 21878 20848
rect 21836 20602 21864 20839
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21822 20496 21878 20505
rect 21822 20431 21878 20440
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21652 13938 21680 14486
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21456 13320 21508 13326
rect 21284 13280 21456 13308
rect 21456 13262 21508 13268
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 21284 11937 21312 13126
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21376 12170 21404 12582
rect 21468 12374 21496 13262
rect 21744 13190 21772 14350
rect 21836 13870 21864 20431
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21364 12164 21416 12170
rect 21364 12106 21416 12112
rect 21560 12102 21588 12650
rect 21638 12608 21694 12617
rect 21638 12543 21694 12552
rect 21548 12096 21600 12102
rect 21548 12038 21600 12044
rect 21270 11928 21326 11937
rect 21270 11863 21326 11872
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 20916 10118 21128 10146
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20916 9722 20944 9998
rect 20994 9888 21050 9897
rect 20994 9823 21050 9832
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20718 7576 20774 7585
rect 20718 7511 20774 7520
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20350 3360 20406 3369
rect 20350 3295 20406 3304
rect 20456 3097 20484 5850
rect 20548 4049 20576 6734
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20640 5370 20668 5510
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20534 4040 20590 4049
rect 20534 3975 20590 3984
rect 20640 3913 20668 4422
rect 20626 3904 20682 3913
rect 20626 3839 20682 3848
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20442 3088 20498 3097
rect 20442 3023 20498 3032
rect 20640 2922 20668 3538
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20180 1278 20300 1306
rect 20074 1048 20130 1057
rect 20074 983 20130 992
rect 20180 480 20208 1278
rect 20640 921 20668 2858
rect 20626 912 20682 921
rect 20626 847 20682 856
rect 20732 480 20760 7511
rect 20810 6896 20866 6905
rect 20810 6831 20812 6840
rect 20864 6831 20866 6840
rect 20812 6802 20864 6808
rect 20812 6180 20864 6186
rect 20812 6122 20864 6128
rect 20824 5914 20852 6122
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20916 4690 20944 9522
rect 21008 9081 21036 9823
rect 20994 9072 21050 9081
rect 20994 9007 21050 9016
rect 21008 8906 21036 9007
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 21100 7546 21128 10118
rect 21284 9976 21312 11630
rect 21560 11336 21588 12038
rect 21652 11898 21680 12543
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21640 11348 21692 11354
rect 21560 11308 21640 11336
rect 21640 11290 21692 11296
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21468 10810 21496 11086
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21652 10742 21680 11290
rect 21640 10736 21692 10742
rect 21640 10678 21692 10684
rect 21454 10432 21510 10441
rect 21454 10367 21510 10376
rect 21364 10192 21416 10198
rect 21364 10134 21416 10140
rect 21192 9948 21312 9976
rect 21192 9586 21220 9948
rect 21376 9761 21404 10134
rect 21362 9752 21418 9761
rect 21272 9716 21324 9722
rect 21468 9722 21496 10367
rect 21546 9888 21602 9897
rect 21546 9823 21602 9832
rect 21362 9687 21418 9696
rect 21456 9716 21508 9722
rect 21272 9658 21324 9664
rect 21456 9658 21508 9664
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21192 9178 21220 9318
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21180 9036 21232 9042
rect 21180 8978 21232 8984
rect 21192 8242 21220 8978
rect 21284 8634 21312 9658
rect 21560 9568 21588 9823
rect 21468 9540 21588 9568
rect 21468 9110 21496 9540
rect 21652 9500 21680 10678
rect 21928 9874 21956 23258
rect 22020 21026 22048 24618
rect 22204 24585 22232 24754
rect 22296 24682 22324 25094
rect 22284 24676 22336 24682
rect 22284 24618 22336 24624
rect 22190 24576 22246 24585
rect 22190 24511 22246 24520
rect 22100 24200 22152 24206
rect 22296 24188 22324 24618
rect 22100 24142 22152 24148
rect 22204 24160 22324 24188
rect 22112 23866 22140 24142
rect 22100 23860 22152 23866
rect 22100 23802 22152 23808
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 22112 23186 22140 23530
rect 22204 23526 22232 24160
rect 22192 23520 22244 23526
rect 22192 23462 22244 23468
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 22112 22794 22140 23122
rect 22204 22982 22232 23462
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22112 22766 22232 22794
rect 22098 22672 22154 22681
rect 22098 22607 22154 22616
rect 22112 22574 22140 22607
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 22204 22438 22232 22766
rect 22388 22642 22416 25162
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 22112 21554 22140 21626
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22100 21344 22152 21350
rect 22098 21312 22100 21321
rect 22152 21312 22154 21321
rect 22098 21247 22154 21256
rect 22020 20998 22140 21026
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 22020 20312 22048 20742
rect 22112 20602 22140 20998
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22100 20324 22152 20330
rect 22020 20284 22100 20312
rect 22100 20266 22152 20272
rect 22112 20233 22140 20266
rect 22098 20224 22154 20233
rect 22098 20159 22154 20168
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22112 19514 22140 19858
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22112 18970 22140 19450
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22020 18426 22048 18702
rect 22204 18442 22232 22374
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 18902 22324 21830
rect 22376 21480 22428 21486
rect 22374 21448 22376 21457
rect 22428 21448 22430 21457
rect 22374 21383 22430 21392
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22388 20466 22416 20742
rect 22480 20534 22508 25327
rect 22560 24064 22612 24070
rect 22664 24041 22692 27520
rect 23216 25906 23244 27520
rect 23204 25900 23256 25906
rect 23204 25842 23256 25848
rect 23768 25838 23796 27520
rect 24320 26110 24348 27520
rect 24766 27160 24822 27169
rect 24766 27095 24822 27104
rect 24780 26518 24808 27095
rect 24768 26512 24820 26518
rect 24768 26454 24820 26460
rect 24308 26104 24360 26110
rect 24214 26072 24270 26081
rect 24308 26046 24360 26052
rect 24214 26007 24270 26016
rect 23756 25832 23808 25838
rect 23756 25774 23808 25780
rect 23020 25356 23072 25362
rect 23020 25298 23072 25304
rect 24124 25356 24176 25362
rect 24124 25298 24176 25304
rect 23032 24886 23060 25298
rect 23664 25152 23716 25158
rect 23386 25120 23442 25129
rect 23664 25094 23716 25100
rect 23386 25055 23442 25064
rect 23020 24880 23072 24886
rect 23020 24822 23072 24828
rect 22928 24676 22980 24682
rect 22928 24618 22980 24624
rect 22836 24336 22888 24342
rect 22836 24278 22888 24284
rect 22560 24006 22612 24012
rect 22650 24032 22706 24041
rect 22572 23662 22600 24006
rect 22650 23967 22706 23976
rect 22848 23905 22876 24278
rect 22834 23896 22890 23905
rect 22834 23831 22836 23840
rect 22888 23831 22890 23840
rect 22836 23802 22888 23808
rect 22848 23771 22876 23802
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22572 21962 22600 23598
rect 22836 23588 22888 23594
rect 22836 23530 22888 23536
rect 22848 23497 22876 23530
rect 22834 23488 22890 23497
rect 22834 23423 22890 23432
rect 22834 23216 22890 23225
rect 22834 23151 22890 23160
rect 22652 23112 22704 23118
rect 22652 23054 22704 23060
rect 22664 22098 22692 23054
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22560 21956 22612 21962
rect 22560 21898 22612 21904
rect 22664 21690 22692 22034
rect 22756 22030 22784 22918
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22848 21894 22876 23151
rect 22940 22137 22968 24618
rect 23032 24410 23060 24822
rect 23296 24608 23348 24614
rect 23296 24550 23348 24556
rect 23020 24404 23072 24410
rect 23020 24346 23072 24352
rect 23308 24274 23336 24550
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 23400 24206 23428 25055
rect 23480 24744 23532 24750
rect 23480 24686 23532 24692
rect 23492 24614 23520 24686
rect 23676 24682 23704 25094
rect 24136 24750 24164 25298
rect 24228 24954 24256 26007
rect 24766 25528 24822 25537
rect 24766 25463 24768 25472
rect 24820 25463 24822 25472
rect 24768 25434 24820 25440
rect 24872 25430 24900 27520
rect 25228 26784 25280 26790
rect 25424 26738 25452 27520
rect 25228 26726 25280 26732
rect 24860 25424 24912 25430
rect 24860 25366 24912 25372
rect 25042 25392 25098 25401
rect 25042 25327 25098 25336
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24688 24993 24716 25162
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 24674 24984 24730 24993
rect 24216 24948 24268 24954
rect 24674 24919 24730 24928
rect 24216 24890 24268 24896
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 23664 24676 23716 24682
rect 23664 24618 23716 24624
rect 24308 24676 24360 24682
rect 24308 24618 24360 24624
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23110 23760 23166 23769
rect 23110 23695 23166 23704
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 22926 22128 22982 22137
rect 22926 22063 22982 22072
rect 23032 21978 23060 23462
rect 22940 21950 23060 21978
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 22558 21448 22614 21457
rect 22558 21383 22614 21392
rect 22572 20874 22600 21383
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 22742 21312 22798 21321
rect 22560 20868 22612 20874
rect 22560 20810 22612 20816
rect 22664 20754 22692 21286
rect 22742 21247 22798 21256
rect 22572 20726 22692 20754
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22388 18834 22416 20402
rect 22572 20346 22600 20726
rect 22650 20496 22706 20505
rect 22650 20431 22706 20440
rect 22480 20318 22600 20346
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22388 18714 22416 18770
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 22112 18414 22232 18442
rect 22296 18686 22416 18714
rect 22112 18306 22140 18414
rect 22020 18278 22140 18306
rect 22020 16946 22048 18278
rect 22100 18148 22152 18154
rect 22100 18090 22152 18096
rect 22112 17105 22140 18090
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22204 17270 22232 18022
rect 22296 17882 22324 18686
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22388 18222 22416 18566
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22098 17096 22154 17105
rect 22098 17031 22154 17040
rect 22020 16918 22140 16946
rect 22008 16788 22060 16794
rect 22008 16730 22060 16736
rect 22020 16232 22048 16730
rect 22112 16402 22140 16918
rect 22204 16697 22232 17206
rect 22388 17202 22416 18158
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22296 16794 22324 17070
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22376 16720 22428 16726
rect 22190 16688 22246 16697
rect 22376 16662 22428 16668
rect 22190 16623 22246 16632
rect 22112 16374 22232 16402
rect 22100 16244 22152 16250
rect 22020 16204 22100 16232
rect 22100 16186 22152 16192
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 22020 14890 22048 15302
rect 22008 14884 22060 14890
rect 22008 14826 22060 14832
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 22020 11626 22048 14554
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22020 10810 22048 11222
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 22020 10266 22048 10474
rect 22112 10470 22140 15846
rect 22204 13802 22232 16374
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 14074 22324 14214
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22282 13560 22338 13569
rect 22282 13495 22284 13504
rect 22336 13495 22338 13504
rect 22284 13466 22336 13472
rect 22296 12850 22324 13466
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22296 11762 22324 12786
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22296 11354 22324 11698
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22100 10464 22152 10470
rect 22152 10424 22232 10452
rect 22100 10406 22152 10412
rect 22098 10296 22154 10305
rect 22008 10260 22060 10266
rect 22098 10231 22154 10240
rect 22008 10202 22060 10208
rect 21836 9846 21956 9874
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 21836 9602 21864 9846
rect 21836 9574 21956 9602
rect 21560 9472 21680 9500
rect 21456 9104 21508 9110
rect 21456 9046 21508 9052
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21376 8634 21404 8774
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21468 8566 21496 9046
rect 21456 8560 21508 8566
rect 21456 8502 21508 8508
rect 21456 8288 21508 8294
rect 21270 8256 21326 8265
rect 21192 8214 21270 8242
rect 21456 8230 21508 8236
rect 21270 8191 21326 8200
rect 21284 8090 21312 8191
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20994 7304 21050 7313
rect 20994 7239 21050 7248
rect 21008 6905 21036 7239
rect 20994 6896 21050 6905
rect 20994 6831 21050 6840
rect 21008 6730 21036 6831
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20994 4584 21050 4593
rect 20994 4519 20996 4528
rect 21048 4519 21050 4528
rect 20996 4490 21048 4496
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20916 3913 20944 3946
rect 20902 3904 20958 3913
rect 20902 3839 20958 3848
rect 20810 3768 20866 3777
rect 21100 3738 21128 6394
rect 21192 5250 21220 7754
rect 21376 6610 21404 7958
rect 21468 7750 21496 8230
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21468 7313 21496 7686
rect 21454 7304 21510 7313
rect 21454 7239 21510 7248
rect 21560 7041 21588 9472
rect 21640 9104 21692 9110
rect 21640 9046 21692 9052
rect 21652 7954 21680 9046
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21730 8256 21786 8265
rect 21730 8191 21786 8200
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21546 7032 21602 7041
rect 21652 7002 21680 7686
rect 21744 7546 21772 8191
rect 21836 8090 21864 8774
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21836 7721 21864 7822
rect 21822 7712 21878 7721
rect 21822 7647 21878 7656
rect 21822 7576 21878 7585
rect 21732 7540 21784 7546
rect 21822 7511 21878 7520
rect 21732 7482 21784 7488
rect 21836 7342 21864 7511
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21546 6967 21602 6976
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21456 6792 21508 6798
rect 21508 6752 21588 6780
rect 21456 6734 21508 6740
rect 21560 6633 21588 6752
rect 21546 6624 21602 6633
rect 21376 6582 21496 6610
rect 21272 6384 21324 6390
rect 21270 6352 21272 6361
rect 21324 6352 21326 6361
rect 21270 6287 21326 6296
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 21376 5370 21404 5714
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21192 5222 21312 5250
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 20810 3703 20812 3712
rect 20864 3703 20866 3712
rect 21088 3732 21140 3738
rect 20812 3674 20864 3680
rect 21088 3674 21140 3680
rect 21192 3505 21220 4694
rect 21178 3496 21234 3505
rect 21178 3431 21180 3440
rect 21232 3431 21234 3440
rect 21180 3402 21232 3408
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 20916 2310 20944 2518
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 16394 439 16450 448
rect 16486 0 16542 480
rect 17038 0 17094 480
rect 17590 0 17646 480
rect 18142 0 18198 480
rect 18602 0 18658 480
rect 19154 0 19210 480
rect 19706 0 19762 480
rect 20166 0 20222 480
rect 20718 0 20774 480
rect 20916 105 20944 2246
rect 21284 480 21312 5222
rect 21376 4826 21404 5306
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 21376 3777 21404 4626
rect 21468 4321 21496 6582
rect 21602 6582 21680 6610
rect 21546 6559 21602 6568
rect 21546 6488 21602 6497
rect 21546 6423 21602 6432
rect 21560 5522 21588 6423
rect 21652 5914 21680 6582
rect 21744 6186 21772 6802
rect 21928 6730 21956 9574
rect 22020 9432 22048 9862
rect 22112 9738 22140 10231
rect 22204 9874 22232 10424
rect 22388 10305 22416 16662
rect 22480 12753 22508 20318
rect 22560 20256 22612 20262
rect 22560 20198 22612 20204
rect 22572 17626 22600 20198
rect 22664 18426 22692 20431
rect 22756 19802 22784 21247
rect 22848 21010 22876 21558
rect 22940 21418 22968 21950
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 22928 21412 22980 21418
rect 22928 21354 22980 21360
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 22836 21004 22888 21010
rect 22836 20946 22888 20952
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22848 19922 22876 20742
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22756 19774 22876 19802
rect 22744 19712 22796 19718
rect 22744 19654 22796 19660
rect 22756 19446 22784 19654
rect 22744 19440 22796 19446
rect 22744 19382 22796 19388
rect 22744 18896 22796 18902
rect 22744 18838 22796 18844
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22572 17598 22692 17626
rect 22560 17536 22612 17542
rect 22558 17504 22560 17513
rect 22612 17504 22614 17513
rect 22558 17439 22614 17448
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22572 16658 22600 17274
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22572 16250 22600 16594
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 22558 15600 22614 15609
rect 22558 15535 22614 15544
rect 22572 13734 22600 15535
rect 22664 14929 22692 17598
rect 22650 14920 22706 14929
rect 22650 14855 22706 14864
rect 22756 14822 22784 18838
rect 22848 18698 22876 19774
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 22836 17808 22888 17814
rect 22836 17750 22888 17756
rect 22848 17338 22876 17750
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22664 14414 22692 14758
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22664 13870 22692 14350
rect 22744 14272 22796 14278
rect 22848 14249 22876 16526
rect 22744 14214 22796 14220
rect 22834 14240 22890 14249
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22572 13569 22600 13670
rect 22558 13560 22614 13569
rect 22664 13530 22692 13806
rect 22558 13495 22614 13504
rect 22652 13524 22704 13530
rect 22572 13394 22600 13495
rect 22652 13466 22704 13472
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22466 12744 22522 12753
rect 22466 12679 22522 12688
rect 22664 12646 22692 13466
rect 22756 13433 22784 14214
rect 22834 14175 22890 14184
rect 22940 13920 22968 21082
rect 23032 20874 23060 21830
rect 23124 21026 23152 23695
rect 23216 21146 23244 24006
rect 23400 23594 23428 24142
rect 23492 23798 23520 24550
rect 23480 23792 23532 23798
rect 23480 23734 23532 23740
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 23492 23474 23520 23530
rect 23768 23497 23796 24550
rect 24320 24274 24348 24618
rect 24780 24449 24808 25094
rect 25056 24750 25084 25327
rect 25240 25140 25268 26726
rect 25332 26710 25452 26738
rect 25332 25294 25360 26710
rect 25410 26616 25466 26625
rect 25410 26551 25466 26560
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25240 25112 25360 25140
rect 25136 24880 25188 24886
rect 25136 24822 25188 24828
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 24766 24440 24822 24449
rect 24766 24375 24822 24384
rect 24308 24268 24360 24274
rect 24308 24210 24360 24216
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24320 24120 24348 24210
rect 24228 24092 24348 24120
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24032 23792 24084 23798
rect 24032 23734 24084 23740
rect 23940 23520 23992 23526
rect 23308 23446 23520 23474
rect 23754 23488 23810 23497
rect 23308 21729 23336 23446
rect 23940 23462 23992 23468
rect 23754 23423 23810 23432
rect 23572 23248 23624 23254
rect 23572 23190 23624 23196
rect 23386 22808 23442 22817
rect 23442 22752 23520 22760
rect 23386 22743 23388 22752
rect 23440 22732 23520 22752
rect 23388 22714 23440 22720
rect 23492 22438 23520 22732
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23400 22250 23428 22374
rect 23400 22222 23520 22250
rect 23388 22160 23440 22166
rect 23388 22102 23440 22108
rect 23294 21720 23350 21729
rect 23294 21655 23350 21664
rect 23400 21298 23428 22102
rect 23492 22030 23520 22222
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23584 21962 23612 23190
rect 23756 23044 23808 23050
rect 23756 22986 23808 22992
rect 23768 22710 23796 22986
rect 23952 22982 23980 23462
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23756 22704 23808 22710
rect 23756 22646 23808 22652
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23664 22500 23716 22506
rect 23664 22442 23716 22448
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23676 21894 23704 22442
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23664 21888 23716 21894
rect 23584 21836 23664 21842
rect 23584 21830 23716 21836
rect 23584 21814 23704 21830
rect 23400 21270 23520 21298
rect 23204 21140 23256 21146
rect 23204 21082 23256 21088
rect 23124 20998 23244 21026
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 23020 20868 23072 20874
rect 23020 20810 23072 20816
rect 23124 19990 23152 20878
rect 23112 19984 23164 19990
rect 23112 19926 23164 19932
rect 23020 19304 23072 19310
rect 23018 19272 23020 19281
rect 23072 19272 23074 19281
rect 23018 19207 23074 19216
rect 23112 19236 23164 19242
rect 23112 19178 23164 19184
rect 23020 18896 23072 18902
rect 23020 18838 23072 18844
rect 23032 18154 23060 18838
rect 23020 18148 23072 18154
rect 23020 18090 23072 18096
rect 23124 17814 23152 19178
rect 23112 17808 23164 17814
rect 23112 17750 23164 17756
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 23032 15910 23060 16934
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 23018 15328 23074 15337
rect 23018 15263 23074 15272
rect 23032 15162 23060 15263
rect 23020 15156 23072 15162
rect 23020 15098 23072 15104
rect 23032 14890 23060 15098
rect 23020 14884 23072 14890
rect 23020 14826 23072 14832
rect 23018 14104 23074 14113
rect 23018 14039 23020 14048
rect 23072 14039 23074 14048
rect 23020 14010 23072 14016
rect 22848 13892 22968 13920
rect 22742 13424 22798 13433
rect 22742 13359 22798 13368
rect 22848 12866 22876 13892
rect 22928 13796 22980 13802
rect 22928 13738 22980 13744
rect 22940 13462 22968 13738
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22756 12838 22876 12866
rect 22652 12640 22704 12646
rect 22466 12608 22522 12617
rect 22652 12582 22704 12588
rect 22466 12543 22522 12552
rect 22480 11506 22508 12543
rect 22664 12374 22692 12582
rect 22652 12368 22704 12374
rect 22652 12310 22704 12316
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22572 11801 22600 12242
rect 22664 11898 22692 12310
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22558 11792 22614 11801
rect 22756 11762 22784 12838
rect 22940 12442 22968 13398
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 22558 11727 22614 11736
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22480 11478 22692 11506
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22480 10538 22508 10950
rect 22468 10532 22520 10538
rect 22468 10474 22520 10480
rect 22374 10296 22430 10305
rect 22374 10231 22430 10240
rect 22468 10192 22520 10198
rect 22468 10134 22520 10140
rect 22480 10033 22508 10134
rect 22466 10024 22522 10033
rect 22466 9959 22522 9968
rect 22204 9846 22416 9874
rect 22112 9710 22232 9738
rect 22020 9404 22140 9432
rect 22006 9208 22062 9217
rect 22006 9143 22008 9152
rect 22060 9143 22062 9152
rect 22008 9114 22060 9120
rect 22112 9110 22140 9404
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 22008 8832 22060 8838
rect 22006 8800 22008 8809
rect 22060 8800 22062 8809
rect 22006 8735 22062 8744
rect 22020 8362 22048 8735
rect 22098 8392 22154 8401
rect 22008 8356 22060 8362
rect 22098 8327 22154 8336
rect 22008 8298 22060 8304
rect 22020 8022 22048 8298
rect 22008 8016 22060 8022
rect 22008 7958 22060 7964
rect 22008 7472 22060 7478
rect 22008 7414 22060 7420
rect 22020 6934 22048 7414
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21836 6322 21864 6598
rect 22008 6384 22060 6390
rect 22008 6326 22060 6332
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 22020 5574 22048 6326
rect 22112 6254 22140 8327
rect 22204 8022 22232 9710
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22296 9489 22324 9658
rect 22282 9480 22338 9489
rect 22282 9415 22338 9424
rect 22296 8294 22324 9415
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 22204 7546 22232 7958
rect 22282 7848 22338 7857
rect 22282 7783 22338 7792
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22190 7440 22246 7449
rect 22190 7375 22246 7384
rect 22204 7274 22232 7375
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22008 5568 22060 5574
rect 21560 5494 21772 5522
rect 22008 5510 22060 5516
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21454 4312 21510 4321
rect 21454 4247 21510 4256
rect 21560 4078 21588 4558
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21652 3890 21680 4218
rect 21560 3862 21680 3890
rect 21362 3768 21418 3777
rect 21362 3703 21418 3712
rect 21560 3670 21588 3862
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 21548 3664 21600 3670
rect 21548 3606 21600 3612
rect 21560 3534 21588 3606
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 21560 3126 21588 3470
rect 21548 3120 21600 3126
rect 21548 3062 21600 3068
rect 21560 2514 21588 3062
rect 21652 3058 21680 3674
rect 21640 3052 21692 3058
rect 21640 2994 21692 3000
rect 21744 2922 21772 5494
rect 22020 5370 22048 5510
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 22296 5234 22324 7783
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 21914 5128 21970 5137
rect 21914 5063 21970 5072
rect 22282 5128 22338 5137
rect 22388 5114 22416 9846
rect 22466 9752 22522 9761
rect 22466 9687 22522 9696
rect 22480 6202 22508 9687
rect 22572 8838 22600 11018
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22572 8673 22600 8774
rect 22558 8664 22614 8673
rect 22558 8599 22614 8608
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 22572 8129 22600 8230
rect 22558 8120 22614 8129
rect 22558 8055 22614 8064
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22572 7002 22600 7482
rect 22664 7018 22692 11478
rect 22834 11384 22890 11393
rect 23124 11370 23152 17750
rect 23216 16697 23244 20998
rect 23296 21004 23348 21010
rect 23296 20946 23348 20952
rect 23308 19922 23336 20946
rect 23492 20602 23520 21270
rect 23584 20641 23612 21814
rect 23676 21765 23704 21814
rect 23768 21554 23796 22170
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23756 21072 23808 21078
rect 23756 21014 23808 21020
rect 23662 20768 23718 20777
rect 23662 20703 23718 20712
rect 23570 20632 23626 20641
rect 23480 20596 23532 20602
rect 23570 20567 23626 20576
rect 23480 20538 23532 20544
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23296 19780 23348 19786
rect 23296 19722 23348 19728
rect 23202 16688 23258 16697
rect 23202 16623 23258 16632
rect 23308 16590 23336 19722
rect 23400 16726 23428 20334
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23492 20097 23520 20198
rect 23478 20088 23534 20097
rect 23478 20023 23534 20032
rect 23572 19984 23624 19990
rect 23572 19926 23624 19932
rect 23480 19848 23532 19854
rect 23478 19816 23480 19825
rect 23532 19816 23534 19825
rect 23478 19751 23534 19760
rect 23584 19666 23612 19926
rect 23492 19638 23612 19666
rect 23492 19174 23520 19638
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23492 18329 23520 19110
rect 23478 18320 23534 18329
rect 23478 18255 23534 18264
rect 23584 17105 23612 19314
rect 23676 19258 23704 20703
rect 23768 20097 23796 21014
rect 23754 20088 23810 20097
rect 23754 20023 23810 20032
rect 23768 19514 23796 20023
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 23860 19378 23888 22510
rect 23848 19372 23900 19378
rect 23848 19314 23900 19320
rect 23676 19230 23796 19258
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23676 18630 23704 19110
rect 23664 18624 23716 18630
rect 23662 18592 23664 18601
rect 23716 18592 23718 18601
rect 23662 18527 23718 18536
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23676 18193 23704 18362
rect 23662 18184 23718 18193
rect 23662 18119 23718 18128
rect 23662 18048 23718 18057
rect 23662 17983 23718 17992
rect 23676 17882 23704 17983
rect 23768 17882 23796 19230
rect 23848 19236 23900 19242
rect 23848 19178 23900 19184
rect 23860 18290 23888 19178
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23952 18034 23980 22918
rect 24044 21554 24072 23734
rect 24136 23594 24164 24006
rect 24228 23730 24256 24092
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 24124 23588 24176 23594
rect 24124 23530 24176 23536
rect 24780 23225 24808 24006
rect 24858 23624 24914 23633
rect 24858 23559 24914 23568
rect 24872 23322 24900 23559
rect 24964 23526 24992 24210
rect 24952 23520 25004 23526
rect 24950 23488 24952 23497
rect 25004 23488 25006 23497
rect 24950 23423 25006 23432
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24766 23216 24822 23225
rect 24766 23151 24822 23160
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24124 23044 24176 23050
rect 24124 22986 24176 22992
rect 24136 22642 24164 22986
rect 24676 22976 24728 22982
rect 24676 22918 24728 22924
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24216 22160 24268 22166
rect 24216 22102 24268 22108
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 24136 21486 24164 22034
rect 24124 21480 24176 21486
rect 24124 21422 24176 21428
rect 24032 21412 24084 21418
rect 24032 21354 24084 21360
rect 24044 20806 24072 21354
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 24136 20330 24164 20946
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 24124 20324 24176 20330
rect 24124 20266 24176 20272
rect 24044 19854 24072 20266
rect 24122 20224 24178 20233
rect 24122 20159 24178 20168
rect 24136 20058 24164 20159
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 24124 19712 24176 19718
rect 24124 19654 24176 19660
rect 24030 19544 24086 19553
rect 24030 19479 24086 19488
rect 24044 19378 24072 19479
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 24032 19236 24084 19242
rect 24032 19178 24084 19184
rect 24044 19145 24072 19178
rect 24030 19136 24086 19145
rect 24030 19071 24086 19080
rect 24044 18970 24072 19071
rect 24032 18964 24084 18970
rect 24032 18906 24084 18912
rect 24032 18692 24084 18698
rect 24032 18634 24084 18640
rect 24044 18222 24072 18634
rect 24136 18329 24164 19654
rect 24228 19496 24256 22102
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21162 24716 22918
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24780 22166 24808 22646
rect 24872 22522 24900 23122
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24964 22642 24992 23054
rect 25148 22778 25176 24822
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25332 22658 25360 25112
rect 25424 24614 25452 26551
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25516 23662 25544 26182
rect 25870 25800 25926 25809
rect 25870 25735 25926 25744
rect 25686 23896 25742 23905
rect 25686 23831 25688 23840
rect 25740 23831 25742 23840
rect 25688 23802 25740 23808
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 25148 22630 25360 22658
rect 25594 22672 25650 22681
rect 24872 22494 24992 22522
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24768 22160 24820 22166
rect 24768 22102 24820 22108
rect 24872 21978 24900 22374
rect 24964 22030 24992 22494
rect 24780 21962 24900 21978
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24768 21956 24900 21962
rect 24820 21950 24900 21956
rect 24768 21898 24820 21904
rect 24766 21720 24822 21729
rect 24766 21655 24768 21664
rect 24820 21655 24822 21664
rect 24768 21626 24820 21632
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 24858 21176 24914 21185
rect 24688 21134 24808 21162
rect 24676 21072 24728 21078
rect 24676 21014 24728 21020
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24308 20324 24360 20330
rect 24308 20266 24360 20272
rect 24320 19786 24348 20266
rect 24688 20262 24716 21014
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 24688 19961 24716 20198
rect 24674 19952 24730 19961
rect 24780 19938 24808 21134
rect 24858 21111 24860 21120
rect 24912 21111 24914 21120
rect 24860 21082 24912 21088
rect 25056 21078 25084 21490
rect 25044 21072 25096 21078
rect 25044 21014 25096 21020
rect 25044 20868 25096 20874
rect 25044 20810 25096 20816
rect 25056 20262 25084 20810
rect 25148 20754 25176 22630
rect 25594 22607 25650 22616
rect 25228 22568 25280 22574
rect 25228 22510 25280 22516
rect 25240 22137 25268 22510
rect 25320 22500 25372 22506
rect 25320 22442 25372 22448
rect 25226 22128 25282 22137
rect 25226 22063 25282 22072
rect 25332 21962 25360 22442
rect 25410 21992 25466 22001
rect 25320 21956 25372 21962
rect 25410 21927 25466 21936
rect 25320 21898 25372 21904
rect 25228 21888 25280 21894
rect 25228 21830 25280 21836
rect 25240 21486 25268 21830
rect 25228 21480 25280 21486
rect 25226 21448 25228 21457
rect 25280 21448 25282 21457
rect 25226 21383 25282 21392
rect 25332 21350 25360 21898
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25332 20874 25360 21286
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 25148 20726 25360 20754
rect 25134 20632 25190 20641
rect 25134 20567 25190 20576
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 24780 19910 24900 19938
rect 24674 19887 24730 19896
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24308 19780 24360 19786
rect 24308 19722 24360 19728
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24228 19468 24440 19496
rect 24214 19408 24270 19417
rect 24214 19343 24270 19352
rect 24308 19372 24360 19378
rect 24228 19242 24256 19343
rect 24308 19314 24360 19320
rect 24216 19236 24268 19242
rect 24216 19178 24268 19184
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24228 18426 24256 18702
rect 24320 18698 24348 19314
rect 24412 18698 24440 19468
rect 24582 19408 24638 19417
rect 24492 19372 24544 19378
rect 24582 19343 24638 19352
rect 24492 19314 24544 19320
rect 24504 19145 24532 19314
rect 24490 19136 24546 19145
rect 24490 19071 24546 19080
rect 24596 18986 24624 19343
rect 24688 19281 24716 19722
rect 24780 19530 24808 19790
rect 24872 19666 24900 19910
rect 24872 19638 24992 19666
rect 24780 19514 24900 19530
rect 24768 19508 24900 19514
rect 24820 19502 24900 19508
rect 24768 19450 24820 19456
rect 24780 19419 24808 19450
rect 24674 19272 24730 19281
rect 24674 19207 24676 19216
rect 24728 19207 24730 19216
rect 24676 19178 24728 19184
rect 24596 18958 24808 18986
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24308 18692 24360 18698
rect 24308 18634 24360 18640
rect 24400 18692 24452 18698
rect 24400 18634 24452 18640
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 24122 18320 24178 18329
rect 24122 18255 24178 18264
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 24136 18154 24164 18255
rect 24124 18148 24176 18154
rect 24124 18090 24176 18096
rect 24688 18086 24716 18838
rect 24676 18080 24728 18086
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23676 17202 23704 17818
rect 23754 17640 23810 17649
rect 23754 17575 23810 17584
rect 23768 17338 23796 17575
rect 23756 17332 23808 17338
rect 23756 17274 23808 17280
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23570 17096 23626 17105
rect 23570 17031 23626 17040
rect 23388 16720 23440 16726
rect 23388 16662 23440 16668
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23662 16552 23718 16561
rect 23662 16487 23718 16496
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23216 15706 23244 16390
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 23216 15162 23244 15642
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 23308 14958 23336 16390
rect 23478 16280 23534 16289
rect 23478 16215 23480 16224
rect 23532 16215 23534 16224
rect 23480 16186 23532 16192
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23400 15026 23428 16118
rect 23492 15910 23520 16186
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23584 15162 23612 15914
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23308 13433 23336 14758
rect 23400 14618 23428 14962
rect 23478 14648 23534 14657
rect 23388 14612 23440 14618
rect 23478 14583 23534 14592
rect 23388 14554 23440 14560
rect 23388 14476 23440 14482
rect 23492 14464 23520 14583
rect 23440 14436 23520 14464
rect 23388 14418 23440 14424
rect 23400 13530 23428 14418
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23294 13424 23350 13433
rect 23294 13359 23350 13368
rect 23492 12889 23520 13670
rect 23478 12880 23534 12889
rect 23478 12815 23534 12824
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 23308 12322 23336 12582
rect 22834 11319 22890 11328
rect 22940 11342 23152 11370
rect 23216 12294 23336 12322
rect 23388 12300 23440 12306
rect 22848 11286 22876 11319
rect 22836 11280 22888 11286
rect 22836 11222 22888 11228
rect 22848 10674 22876 11222
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22756 10305 22784 10610
rect 22836 10532 22888 10538
rect 22836 10474 22888 10480
rect 22742 10296 22798 10305
rect 22742 10231 22798 10240
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22756 9654 22784 9998
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22756 9042 22784 9590
rect 22848 9178 22876 10474
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22756 7721 22784 8978
rect 22742 7712 22798 7721
rect 22742 7647 22798 7656
rect 22756 7546 22784 7647
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22560 6996 22612 7002
rect 22664 6990 22784 7018
rect 22560 6938 22612 6944
rect 22572 6458 22600 6938
rect 22652 6928 22704 6934
rect 22652 6870 22704 6876
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22480 6174 22600 6202
rect 22572 5114 22600 6174
rect 22664 5914 22692 6870
rect 22652 5908 22704 5914
rect 22652 5850 22704 5856
rect 22756 5846 22784 6990
rect 22848 5953 22876 9114
rect 22834 5944 22890 5953
rect 22834 5879 22890 5888
rect 22744 5840 22796 5846
rect 22744 5782 22796 5788
rect 22834 5400 22890 5409
rect 22834 5335 22890 5344
rect 22388 5086 22508 5114
rect 22572 5086 22784 5114
rect 22282 5063 22284 5072
rect 21822 4176 21878 4185
rect 21822 4111 21878 4120
rect 21732 2916 21784 2922
rect 21732 2858 21784 2864
rect 21730 2680 21786 2689
rect 21730 2615 21786 2624
rect 21548 2508 21600 2514
rect 21548 2450 21600 2456
rect 21744 2446 21772 2615
rect 21732 2440 21784 2446
rect 21362 2408 21418 2417
rect 21732 2382 21784 2388
rect 21362 2343 21364 2352
rect 21416 2343 21418 2352
rect 21364 2314 21416 2320
rect 21836 480 21864 4111
rect 21928 2514 21956 5063
rect 22336 5063 22338 5072
rect 22284 5034 22336 5040
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 22020 3942 22048 4626
rect 22204 4282 22232 4626
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 22388 4185 22416 4966
rect 22480 4554 22508 5086
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22468 4548 22520 4554
rect 22468 4490 22520 4496
rect 22374 4176 22430 4185
rect 22284 4140 22336 4146
rect 22374 4111 22430 4120
rect 22284 4082 22336 4088
rect 22296 4049 22324 4082
rect 22376 4072 22428 4078
rect 22282 4040 22338 4049
rect 22376 4014 22428 4020
rect 22282 3975 22338 3984
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 22388 3738 22416 4014
rect 22480 3754 22508 4490
rect 22560 4480 22612 4486
rect 22560 4422 22612 4428
rect 22572 3942 22600 4422
rect 22560 3936 22612 3942
rect 22664 3913 22692 4966
rect 22756 4010 22784 5086
rect 22848 4758 22876 5335
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 22848 4214 22876 4694
rect 22836 4208 22888 4214
rect 22836 4150 22888 4156
rect 22744 4004 22796 4010
rect 22744 3946 22796 3952
rect 22560 3878 22612 3884
rect 22650 3904 22706 3913
rect 22650 3839 22706 3848
rect 22480 3738 22692 3754
rect 22376 3732 22428 3738
rect 22480 3732 22704 3738
rect 22480 3726 22652 3732
rect 22376 3674 22428 3680
rect 22652 3674 22704 3680
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22376 3460 22428 3466
rect 22376 3402 22428 3408
rect 22282 3360 22338 3369
rect 22282 3295 22338 3304
rect 21916 2508 21968 2514
rect 21916 2450 21968 2456
rect 22296 480 22324 3295
rect 22388 1737 22416 3402
rect 22480 2825 22508 3538
rect 22560 3392 22612 3398
rect 22560 3334 22612 3340
rect 22572 3233 22600 3334
rect 22558 3224 22614 3233
rect 22664 3194 22692 3674
rect 22742 3632 22798 3641
rect 22742 3567 22798 3576
rect 22558 3159 22614 3168
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22756 2961 22784 3567
rect 22940 3466 22968 11342
rect 23020 11280 23072 11286
rect 23018 11248 23020 11257
rect 23072 11248 23074 11257
rect 23018 11183 23074 11192
rect 23032 10810 23060 11183
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 23124 10266 23152 11086
rect 23216 10674 23244 12294
rect 23388 12242 23440 12248
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23204 10668 23256 10674
rect 23204 10610 23256 10616
rect 23204 10532 23256 10538
rect 23204 10474 23256 10480
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23020 9988 23072 9994
rect 23020 9930 23072 9936
rect 23032 8430 23060 9930
rect 23216 9926 23244 10474
rect 23204 9920 23256 9926
rect 23202 9888 23204 9897
rect 23256 9888 23258 9897
rect 23202 9823 23258 9832
rect 23308 9586 23336 11766
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 23124 8634 23152 9318
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 23112 8356 23164 8362
rect 23112 8298 23164 8304
rect 23018 8120 23074 8129
rect 23018 8055 23074 8064
rect 23032 6934 23060 8055
rect 23020 6928 23072 6934
rect 23020 6870 23072 6876
rect 23032 6186 23060 6870
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 23032 5302 23060 6122
rect 23020 5296 23072 5302
rect 23020 5238 23072 5244
rect 23020 4752 23072 4758
rect 23018 4720 23020 4729
rect 23072 4720 23074 4729
rect 23018 4655 23074 4664
rect 23032 4282 23060 4655
rect 23020 4276 23072 4282
rect 23020 4218 23072 4224
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 22928 3460 22980 3466
rect 22928 3402 22980 3408
rect 23032 3194 23060 3470
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 22834 3088 22890 3097
rect 23124 3074 23152 8298
rect 23216 7818 23244 9454
rect 23400 9058 23428 12242
rect 23492 11529 23520 12815
rect 23676 12186 23704 16487
rect 23756 15632 23808 15638
rect 23756 15574 23808 15580
rect 23768 12986 23796 15574
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23860 12306 23888 18022
rect 23952 18006 24256 18034
rect 24676 18022 24728 18028
rect 24122 17912 24178 17921
rect 24122 17847 24178 17856
rect 24030 17640 24086 17649
rect 24136 17610 24164 17847
rect 24030 17575 24086 17584
rect 24124 17604 24176 17610
rect 23938 17368 23994 17377
rect 23938 17303 23994 17312
rect 23952 16794 23980 17303
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 23952 15706 23980 16730
rect 24044 16153 24072 17575
rect 24124 17546 24176 17552
rect 24228 17184 24256 18006
rect 24398 17776 24454 17785
rect 24398 17711 24400 17720
rect 24452 17711 24454 17720
rect 24400 17682 24452 17688
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17270 24716 17614
rect 24676 17264 24728 17270
rect 24136 17156 24256 17184
rect 24674 17232 24676 17241
rect 24728 17232 24730 17241
rect 24674 17167 24730 17176
rect 24030 16144 24086 16153
rect 24030 16079 24086 16088
rect 24030 15872 24086 15881
rect 24030 15807 24086 15816
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 23938 15192 23994 15201
rect 24044 15178 24072 15807
rect 24136 15314 24164 17156
rect 24214 17096 24270 17105
rect 24214 17031 24270 17040
rect 24676 17060 24728 17066
rect 24228 16998 24256 17031
rect 24676 17002 24728 17008
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24216 16516 24268 16522
rect 24216 16458 24268 16464
rect 24228 16114 24256 16458
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24400 16176 24452 16182
rect 24400 16118 24452 16124
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24214 16008 24270 16017
rect 24214 15943 24270 15952
rect 24228 15434 24256 15943
rect 24412 15706 24440 16118
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 24688 15586 24716 17002
rect 24596 15570 24716 15586
rect 24584 15564 24716 15570
rect 24636 15558 24716 15564
rect 24584 15506 24636 15512
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24216 15428 24268 15434
rect 24216 15370 24268 15376
rect 24136 15286 24256 15314
rect 24044 15150 24164 15178
rect 23938 15127 23994 15136
rect 23952 13870 23980 15127
rect 24032 14884 24084 14890
rect 24032 14826 24084 14832
rect 24044 14793 24072 14826
rect 24030 14784 24086 14793
rect 24030 14719 24086 14728
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 24136 13569 24164 15150
rect 23938 13560 23994 13569
rect 23938 13495 23994 13504
rect 24122 13560 24178 13569
rect 24122 13495 24178 13504
rect 23952 13394 23980 13495
rect 24030 13424 24086 13433
rect 23940 13388 23992 13394
rect 24030 13359 24086 13368
rect 23940 13330 23992 13336
rect 24044 13002 24072 13359
rect 24124 13184 24176 13190
rect 24122 13152 24124 13161
rect 24176 13152 24178 13161
rect 24122 13087 24178 13096
rect 24044 12974 24164 13002
rect 24030 12744 24086 12753
rect 24030 12679 24086 12688
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23676 12158 23980 12186
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23846 12064 23902 12073
rect 23478 11520 23534 11529
rect 23478 11455 23534 11464
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23492 11218 23520 11290
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 23492 10810 23520 11154
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23570 10840 23626 10849
rect 23480 10804 23532 10810
rect 23570 10775 23626 10784
rect 23480 10746 23532 10752
rect 23478 10160 23534 10169
rect 23478 10095 23534 10104
rect 23492 9178 23520 10095
rect 23584 9518 23612 10775
rect 23676 10606 23704 10950
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23662 10160 23718 10169
rect 23662 10095 23718 10104
rect 23676 9722 23704 10095
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23768 9568 23796 12038
rect 23846 11999 23902 12008
rect 23676 9540 23796 9568
rect 23572 9512 23624 9518
rect 23572 9454 23624 9460
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23296 9036 23348 9042
rect 23400 9030 23520 9058
rect 23296 8978 23348 8984
rect 23204 7812 23256 7818
rect 23204 7754 23256 7760
rect 23308 7750 23336 8978
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23296 7744 23348 7750
rect 23202 7712 23258 7721
rect 23296 7686 23348 7692
rect 23202 7647 23258 7656
rect 23216 7449 23244 7647
rect 23202 7440 23258 7449
rect 23202 7375 23258 7384
rect 23216 6916 23244 7375
rect 23308 7313 23336 7686
rect 23400 7478 23428 8230
rect 23492 7721 23520 9030
rect 23584 7954 23612 9318
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23584 7857 23612 7890
rect 23570 7848 23626 7857
rect 23570 7783 23626 7792
rect 23478 7712 23534 7721
rect 23478 7647 23534 7656
rect 23478 7576 23534 7585
rect 23478 7511 23480 7520
rect 23532 7511 23534 7520
rect 23480 7482 23532 7488
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 23294 7304 23350 7313
rect 23294 7239 23350 7248
rect 23216 6888 23336 6916
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23216 6633 23244 6734
rect 23202 6624 23258 6633
rect 23202 6559 23258 6568
rect 23216 6118 23244 6559
rect 23308 6168 23336 6888
rect 23400 6390 23428 7414
rect 23478 7168 23534 7177
rect 23478 7103 23534 7112
rect 23492 6866 23520 7103
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23308 6140 23520 6168
rect 23204 6112 23256 6118
rect 23256 6072 23336 6100
rect 23204 6054 23256 6060
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 22834 3023 22890 3032
rect 23032 3046 23152 3074
rect 22742 2952 22798 2961
rect 22742 2887 22798 2896
rect 22466 2816 22522 2825
rect 22466 2751 22522 2760
rect 22480 2650 22508 2751
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22374 1728 22430 1737
rect 22374 1663 22430 1672
rect 22848 480 22876 3023
rect 22926 1184 22982 1193
rect 22926 1119 22982 1128
rect 22940 513 22968 1119
rect 23032 785 23060 3046
rect 23216 1057 23244 3130
rect 23202 1048 23258 1057
rect 23202 983 23258 992
rect 23308 921 23336 6072
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23400 5370 23428 5782
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23492 5166 23520 6140
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23492 4457 23520 4966
rect 23478 4448 23534 4457
rect 23478 4383 23534 4392
rect 23584 4162 23612 7414
rect 23400 4134 23612 4162
rect 23400 4078 23428 4134
rect 23388 4072 23440 4078
rect 23676 4026 23704 9540
rect 23860 8566 23888 11999
rect 23952 10674 23980 12158
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 23952 10441 23980 10474
rect 23938 10432 23994 10441
rect 23938 10367 23994 10376
rect 23952 10266 23980 10367
rect 23940 10260 23992 10266
rect 23940 10202 23992 10208
rect 23940 10124 23992 10130
rect 23940 10066 23992 10072
rect 23952 9654 23980 10066
rect 23940 9648 23992 9654
rect 23940 9590 23992 9596
rect 23952 8838 23980 9590
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23848 8560 23900 8566
rect 23848 8502 23900 8508
rect 23952 8378 23980 8774
rect 23860 8350 23980 8378
rect 23756 8016 23808 8022
rect 23756 7958 23808 7964
rect 23768 4282 23796 7958
rect 23756 4276 23808 4282
rect 23756 4218 23808 4224
rect 23756 4072 23808 4078
rect 23388 4014 23440 4020
rect 23492 3998 23704 4026
rect 23754 4040 23756 4049
rect 23808 4040 23810 4049
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23400 3670 23428 3878
rect 23388 3664 23440 3670
rect 23388 3606 23440 3612
rect 23386 3088 23442 3097
rect 23386 3023 23442 3032
rect 23294 912 23350 921
rect 23294 847 23350 856
rect 23018 776 23074 785
rect 23018 711 23074 720
rect 22926 504 22982 513
rect 20902 96 20958 105
rect 20902 31 20958 40
rect 21270 0 21326 480
rect 21822 0 21878 480
rect 22282 0 22338 480
rect 22834 0 22890 480
rect 23400 480 23428 3023
rect 23492 2446 23520 3998
rect 23754 3975 23810 3984
rect 23860 3890 23888 8350
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 23952 6474 23980 8230
rect 24044 6730 24072 12679
rect 24136 11082 24164 12974
rect 24228 12782 24256 15286
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 15438
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24780 13818 24808 18958
rect 24872 18766 24900 19502
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24872 17882 24900 18226
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24872 16794 24900 17682
rect 24964 16810 24992 19638
rect 25056 19446 25084 20198
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 25044 18896 25096 18902
rect 25042 18864 25044 18873
rect 25096 18864 25098 18873
rect 25042 18799 25098 18808
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25056 18426 25084 18702
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 25056 17746 25084 18158
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 24860 16788 24912 16794
rect 24964 16782 25084 16810
rect 25148 16794 25176 20567
rect 25228 20392 25280 20398
rect 25226 20360 25228 20369
rect 25280 20360 25282 20369
rect 25226 20295 25282 20304
rect 25226 19816 25282 19825
rect 25226 19751 25228 19760
rect 25280 19751 25282 19760
rect 25228 19722 25280 19728
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25240 19009 25268 19246
rect 25226 19000 25282 19009
rect 25226 18935 25282 18944
rect 25332 17354 25360 20726
rect 25424 19174 25452 21927
rect 25504 21412 25556 21418
rect 25504 21354 25556 21360
rect 25516 21049 25544 21354
rect 25502 21040 25558 21049
rect 25502 20975 25558 20984
rect 25502 19952 25558 19961
rect 25502 19887 25558 19896
rect 25412 19168 25464 19174
rect 25412 19110 25464 19116
rect 25240 17326 25360 17354
rect 24860 16730 24912 16736
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 24964 16250 24992 16594
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 24858 15736 24914 15745
rect 24858 15671 24914 15680
rect 24872 14929 24900 15671
rect 24858 14920 24914 14929
rect 24858 14855 24914 14864
rect 24872 13977 24900 14855
rect 24964 14804 24992 15982
rect 25056 14940 25084 16782
rect 25136 16788 25188 16794
rect 25136 16730 25188 16736
rect 25240 16182 25268 17326
rect 25320 17264 25372 17270
rect 25320 17206 25372 17212
rect 25228 16176 25280 16182
rect 25228 16118 25280 16124
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25148 15162 25176 15438
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25136 14952 25188 14958
rect 25056 14912 25136 14940
rect 25136 14894 25188 14900
rect 24964 14776 25176 14804
rect 24858 13968 24914 13977
rect 24858 13903 24914 13912
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24596 13530 24624 13670
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12986 24716 13806
rect 24780 13790 24900 13818
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 24228 11393 24256 12582
rect 24308 12232 24360 12238
rect 24306 12200 24308 12209
rect 24360 12200 24362 12209
rect 24306 12135 24362 12144
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24214 11384 24270 11393
rect 24214 11319 24270 11328
rect 24584 11348 24636 11354
rect 24688 11336 24716 12718
rect 24780 11626 24808 13670
rect 24872 13530 24900 13790
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24952 13320 25004 13326
rect 24950 13288 24952 13297
rect 25004 13288 25006 13297
rect 24950 13223 25006 13232
rect 25056 12918 25084 13330
rect 25044 12912 25096 12918
rect 25044 12854 25096 12860
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 25056 12481 25084 12582
rect 25042 12472 25098 12481
rect 25042 12407 25098 12416
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24858 11928 24914 11937
rect 24858 11863 24914 11872
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 24636 11308 24716 11336
rect 24584 11290 24636 11296
rect 24780 11286 24808 11562
rect 24768 11280 24820 11286
rect 24768 11222 24820 11228
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 24122 10840 24178 10849
rect 24228 10826 24256 11154
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24780 10826 24808 11222
rect 24178 10798 24256 10826
rect 24688 10798 24808 10826
rect 24122 10775 24124 10784
rect 24176 10775 24178 10784
rect 24124 10746 24176 10752
rect 24688 10674 24716 10798
rect 24768 10736 24820 10742
rect 24768 10678 24820 10684
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 24122 10432 24178 10441
rect 24122 10367 24178 10376
rect 24136 8294 24164 10367
rect 24228 9722 24256 10542
rect 24688 9994 24716 10610
rect 24676 9988 24728 9994
rect 24676 9930 24728 9936
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24674 9752 24730 9761
rect 24216 9716 24268 9722
rect 24674 9687 24730 9696
rect 24216 9658 24268 9664
rect 24688 9586 24716 9687
rect 24308 9580 24360 9586
rect 24228 9540 24308 9568
rect 24228 8514 24256 9540
rect 24308 9522 24360 9528
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24674 9344 24730 9353
rect 24674 9279 24730 9288
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24688 8634 24716 9279
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24228 8486 24348 8514
rect 24124 8288 24176 8294
rect 24124 8230 24176 8236
rect 24216 8084 24268 8090
rect 24216 8026 24268 8032
rect 24124 7812 24176 7818
rect 24124 7754 24176 7760
rect 24136 7274 24164 7754
rect 24228 7410 24256 8026
rect 24320 8022 24348 8486
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24400 8356 24452 8362
rect 24400 8298 24452 8304
rect 24308 8016 24360 8022
rect 24308 7958 24360 7964
rect 24412 7954 24440 8298
rect 24688 8242 24716 8434
rect 24780 8344 24808 10678
rect 24872 10169 24900 11863
rect 24964 10441 24992 12174
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25056 11801 25084 11834
rect 25042 11792 25098 11801
rect 25042 11727 25098 11736
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 24950 10432 25006 10441
rect 24950 10367 25006 10376
rect 24858 10160 24914 10169
rect 24858 10095 24914 10104
rect 24858 10024 24914 10033
rect 24858 9959 24914 9968
rect 24872 8974 24900 9959
rect 24952 9920 25004 9926
rect 24950 9888 24952 9897
rect 25004 9888 25006 9897
rect 24950 9823 25006 9832
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 25056 8650 25084 11086
rect 25148 9217 25176 14776
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25240 14074 25268 14214
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25226 13696 25282 13705
rect 25226 13631 25282 13640
rect 25240 12889 25268 13631
rect 25226 12880 25282 12889
rect 25226 12815 25282 12824
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 25240 11150 25268 12174
rect 25332 11354 25360 17206
rect 25516 16250 25544 19887
rect 25608 18426 25636 22607
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 25686 21584 25742 21593
rect 25686 21519 25742 21528
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25594 17912 25650 17921
rect 25594 17847 25650 17856
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25410 16008 25466 16017
rect 25410 15943 25466 15952
rect 25424 14074 25452 15943
rect 25504 14884 25556 14890
rect 25504 14826 25556 14832
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25410 13968 25466 13977
rect 25410 13903 25466 13912
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25424 11234 25452 13903
rect 25516 12782 25544 14826
rect 25608 12986 25636 17847
rect 25700 17338 25728 21519
rect 25792 21146 25820 22170
rect 25780 21140 25832 21146
rect 25780 21082 25832 21088
rect 25780 20936 25832 20942
rect 25778 20904 25780 20913
rect 25832 20904 25834 20913
rect 25778 20839 25834 20848
rect 25780 20324 25832 20330
rect 25780 20266 25832 20272
rect 25792 18426 25820 20266
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25792 18222 25820 18362
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25884 17270 25912 25735
rect 25976 24721 26004 27520
rect 26528 26217 26556 27520
rect 26514 26208 26570 26217
rect 26514 26143 26570 26152
rect 26056 26036 26108 26042
rect 26056 25978 26108 25984
rect 25962 24712 26018 24721
rect 25962 24647 26018 24656
rect 25964 21344 26016 21350
rect 25962 21312 25964 21321
rect 26016 21312 26018 21321
rect 25962 21247 26018 21256
rect 25964 20868 26016 20874
rect 25964 20810 26016 20816
rect 25976 19825 26004 20810
rect 25962 19816 26018 19825
rect 25962 19751 26018 19760
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 25872 17264 25924 17270
rect 25872 17206 25924 17212
rect 25870 17096 25926 17105
rect 25870 17031 25926 17040
rect 25686 16552 25742 16561
rect 25686 16487 25742 16496
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25504 12776 25556 12782
rect 25504 12718 25556 12724
rect 25504 12368 25556 12374
rect 25504 12310 25556 12316
rect 25516 11558 25544 12310
rect 25596 11688 25648 11694
rect 25594 11656 25596 11665
rect 25648 11656 25650 11665
rect 25594 11591 25650 11600
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25332 11206 25452 11234
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 25228 10600 25280 10606
rect 25226 10568 25228 10577
rect 25280 10568 25282 10577
rect 25226 10503 25282 10512
rect 25228 9920 25280 9926
rect 25228 9862 25280 9868
rect 25240 9518 25268 9862
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25134 9208 25190 9217
rect 25134 9143 25190 9152
rect 25056 8622 25176 8650
rect 25044 8560 25096 8566
rect 25042 8528 25044 8537
rect 25096 8528 25098 8537
rect 25042 8463 25098 8472
rect 24780 8316 24900 8344
rect 24688 8214 24808 8242
rect 24400 7948 24452 7954
rect 24400 7890 24452 7896
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7546 24716 7686
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 24582 7032 24638 7041
rect 24582 6967 24638 6976
rect 24596 6934 24624 6967
rect 24584 6928 24636 6934
rect 24584 6870 24636 6876
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 24032 6724 24084 6730
rect 24032 6666 24084 6672
rect 23952 6446 24072 6474
rect 23940 5568 23992 5574
rect 23940 5510 23992 5516
rect 23952 4049 23980 5510
rect 23938 4040 23994 4049
rect 23938 3975 23994 3984
rect 23676 3862 23888 3890
rect 23938 3904 23994 3913
rect 23676 2650 23704 3862
rect 23938 3839 23994 3848
rect 23756 3120 23808 3126
rect 23756 3062 23808 3068
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23662 2544 23718 2553
rect 23768 2514 23796 3062
rect 23662 2479 23718 2488
rect 23756 2508 23808 2514
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23676 2310 23704 2479
rect 23756 2450 23808 2456
rect 23664 2304 23716 2310
rect 23664 2246 23716 2252
rect 23952 480 23980 3839
rect 24044 3466 24072 6446
rect 24228 6186 24256 6802
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 24492 6180 24544 6186
rect 24492 6122 24544 6128
rect 24504 5778 24532 6122
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24492 5772 24544 5778
rect 24492 5714 24544 5720
rect 24228 5114 24256 5714
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5166 24716 5646
rect 24676 5160 24728 5166
rect 24136 5086 24256 5114
rect 24504 5120 24676 5148
rect 24136 4826 24164 5086
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24124 4684 24176 4690
rect 24124 4626 24176 4632
rect 24136 4321 24164 4626
rect 24228 4554 24256 4966
rect 24504 4758 24532 5120
rect 24676 5102 24728 5108
rect 24492 4752 24544 4758
rect 24492 4694 24544 4700
rect 24584 4616 24636 4622
rect 24636 4564 24716 4570
rect 24584 4558 24716 4564
rect 24216 4548 24268 4554
rect 24596 4542 24716 4558
rect 24216 4490 24268 4496
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24122 4312 24178 4321
rect 24289 4304 24585 4324
rect 24122 4247 24178 4256
rect 24136 4214 24164 4247
rect 24124 4208 24176 4214
rect 24124 4150 24176 4156
rect 24584 4072 24636 4078
rect 24122 4040 24178 4049
rect 24584 4014 24636 4020
rect 24122 3975 24178 3984
rect 24216 4004 24268 4010
rect 24032 3460 24084 3466
rect 24032 3402 24084 3408
rect 24136 2961 24164 3975
rect 24216 3946 24268 3952
rect 24308 4004 24360 4010
rect 24308 3946 24360 3952
rect 24228 3602 24256 3946
rect 24320 3738 24348 3946
rect 24596 3913 24624 4014
rect 24688 3942 24716 4542
rect 24676 3936 24728 3942
rect 24582 3904 24638 3913
rect 24676 3878 24728 3884
rect 24582 3839 24638 3848
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24320 3466 24348 3674
rect 24582 3632 24638 3641
rect 24582 3567 24638 3576
rect 24596 3534 24624 3567
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24308 3460 24360 3466
rect 24228 3420 24308 3448
rect 24228 3194 24256 3420
rect 24308 3402 24360 3408
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24122 2952 24178 2961
rect 24122 2887 24178 2896
rect 24032 2372 24084 2378
rect 24032 2314 24084 2320
rect 24044 1170 24072 2314
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24122 2136 24178 2145
rect 24289 2128 24585 2148
rect 24122 2071 24124 2080
rect 24176 2071 24178 2080
rect 24124 2042 24176 2048
rect 24688 1329 24716 3878
rect 24780 2378 24808 8214
rect 24872 8090 24900 8316
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24872 7970 24900 8026
rect 24872 7942 24992 7970
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 24872 6662 24900 7822
rect 24964 7546 24992 7942
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24950 7304 25006 7313
rect 25148 7290 25176 8622
rect 25240 8566 25268 9454
rect 25228 8560 25280 8566
rect 25228 8502 25280 8508
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 25006 7262 25176 7290
rect 24950 7239 25006 7248
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24872 5370 24900 6598
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24858 3224 24914 3233
rect 24858 3159 24914 3168
rect 24872 3126 24900 3159
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 24964 3058 24992 7239
rect 25134 7032 25190 7041
rect 25134 6967 25190 6976
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 25056 5642 25084 6734
rect 25148 5914 25176 6967
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 25240 5778 25268 8230
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25136 5704 25188 5710
rect 25134 5672 25136 5681
rect 25188 5672 25190 5681
rect 25332 5658 25360 11206
rect 25410 10296 25466 10305
rect 25410 10231 25412 10240
rect 25464 10231 25466 10240
rect 25412 10202 25464 10208
rect 25412 9988 25464 9994
rect 25412 9930 25464 9936
rect 25424 8294 25452 9930
rect 25516 9761 25544 11494
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25608 10985 25636 11290
rect 25594 10976 25650 10985
rect 25594 10911 25650 10920
rect 25502 9752 25558 9761
rect 25502 9687 25558 9696
rect 25504 9444 25556 9450
rect 25504 9386 25556 9392
rect 25516 9042 25544 9386
rect 25504 9036 25556 9042
rect 25504 8978 25556 8984
rect 25608 8838 25636 10911
rect 25700 9194 25728 16487
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25792 10674 25820 13806
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25700 9166 25820 9194
rect 25884 9178 25912 17031
rect 25976 13734 26004 19654
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 25962 13560 26018 13569
rect 25962 13495 26018 13504
rect 25976 11898 26004 13495
rect 25964 11892 26016 11898
rect 25964 11834 26016 11840
rect 25962 11248 26018 11257
rect 25962 11183 26018 11192
rect 25976 9994 26004 11183
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 25962 9616 26018 9625
rect 25962 9551 25964 9560
rect 26016 9551 26018 9560
rect 25964 9522 26016 9528
rect 25688 9104 25740 9110
rect 25686 9072 25688 9081
rect 25740 9072 25742 9081
rect 25686 9007 25742 9016
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25596 8560 25648 8566
rect 25596 8502 25648 8508
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25412 8016 25464 8022
rect 25410 7984 25412 7993
rect 25464 7984 25466 7993
rect 25410 7919 25466 7928
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25410 6896 25466 6905
rect 25410 6831 25412 6840
rect 25464 6831 25466 6840
rect 25412 6802 25464 6808
rect 25412 6452 25464 6458
rect 25412 6394 25464 6400
rect 25044 5636 25096 5642
rect 25134 5607 25190 5616
rect 25240 5630 25360 5658
rect 25044 5578 25096 5584
rect 25240 5556 25268 5630
rect 25148 5528 25268 5556
rect 25320 5568 25372 5574
rect 25148 4826 25176 5528
rect 25320 5510 25372 5516
rect 25228 5160 25280 5166
rect 25226 5128 25228 5137
rect 25280 5128 25282 5137
rect 25226 5063 25282 5072
rect 25240 4826 25268 5063
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 25228 4820 25280 4826
rect 25228 4762 25280 4768
rect 25148 4078 25176 4762
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 25044 3528 25096 3534
rect 25042 3496 25044 3505
rect 25096 3496 25098 3505
rect 25042 3431 25098 3440
rect 25148 3097 25176 3878
rect 25134 3088 25190 3097
rect 24952 3052 25004 3058
rect 25134 3023 25190 3032
rect 24952 2994 25004 3000
rect 25228 2984 25280 2990
rect 25134 2952 25190 2961
rect 25228 2926 25280 2932
rect 25134 2887 25190 2896
rect 25148 2650 25176 2887
rect 25136 2644 25188 2650
rect 25136 2586 25188 2592
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 25240 2310 25268 2926
rect 25228 2304 25280 2310
rect 25228 2246 25280 2252
rect 24950 1456 25006 1465
rect 24950 1391 25006 1400
rect 24674 1320 24730 1329
rect 24674 1255 24730 1264
rect 24044 1142 24440 1170
rect 24412 480 24440 1142
rect 24964 480 24992 1391
rect 25332 1193 25360 5510
rect 25424 4570 25452 6394
rect 25516 5234 25544 7142
rect 25504 5228 25556 5234
rect 25504 5170 25556 5176
rect 25504 5092 25556 5098
rect 25504 5034 25556 5040
rect 25516 4865 25544 5034
rect 25502 4856 25558 4865
rect 25502 4791 25558 4800
rect 25424 4542 25544 4570
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 25424 4078 25452 4422
rect 25412 4072 25464 4078
rect 25412 4014 25464 4020
rect 25424 3058 25452 4014
rect 25516 4010 25544 4542
rect 25504 4004 25556 4010
rect 25504 3946 25556 3952
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25608 2854 25636 8502
rect 25686 8256 25742 8265
rect 25686 8191 25742 8200
rect 25700 8090 25728 8191
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25792 7546 25820 9166
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 25688 6928 25740 6934
rect 25688 6870 25740 6876
rect 25700 6118 25728 6870
rect 25780 6792 25832 6798
rect 25778 6760 25780 6769
rect 25832 6760 25834 6769
rect 25778 6695 25834 6704
rect 25884 6186 25912 8774
rect 25976 8634 26004 9114
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 25962 6352 26018 6361
rect 25962 6287 25964 6296
rect 26016 6287 26018 6296
rect 25964 6258 26016 6264
rect 25872 6180 25924 6186
rect 25872 6122 25924 6128
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 25870 6080 25926 6089
rect 25596 2848 25648 2854
rect 25596 2790 25648 2796
rect 25412 2440 25464 2446
rect 25410 2408 25412 2417
rect 25596 2440 25648 2446
rect 25464 2408 25466 2417
rect 25596 2382 25648 2388
rect 25410 2343 25466 2352
rect 25502 2000 25558 2009
rect 25502 1935 25558 1944
rect 25318 1184 25374 1193
rect 25318 1119 25374 1128
rect 25516 480 25544 1935
rect 25608 1601 25636 2382
rect 25594 1592 25650 1601
rect 25594 1527 25650 1536
rect 25700 1465 25728 6054
rect 25870 6015 25926 6024
rect 25884 5914 25912 6015
rect 25872 5908 25924 5914
rect 25872 5850 25924 5856
rect 25872 5772 25924 5778
rect 25872 5714 25924 5720
rect 25778 5400 25834 5409
rect 25884 5370 25912 5714
rect 25964 5636 26016 5642
rect 25964 5578 26016 5584
rect 25778 5335 25834 5344
rect 25872 5364 25924 5370
rect 25792 2106 25820 5335
rect 25872 5306 25924 5312
rect 25780 2100 25832 2106
rect 25780 2042 25832 2048
rect 25976 2009 26004 5578
rect 25962 2000 26018 2009
rect 25962 1935 26018 1944
rect 25686 1456 25742 1465
rect 25686 1391 25742 1400
rect 26068 480 26096 25978
rect 27080 25673 27108 27520
rect 27632 25770 27660 27520
rect 27620 25764 27672 25770
rect 27620 25706 27672 25712
rect 27066 25664 27122 25673
rect 27066 25599 27122 25608
rect 26330 22264 26386 22273
rect 26330 22199 26386 22208
rect 26344 21690 26372 22199
rect 26332 21684 26384 21690
rect 26332 21626 26384 21632
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26160 16046 26188 21422
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26344 20097 26372 20198
rect 26330 20088 26386 20097
rect 26330 20023 26386 20032
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 26240 18352 26292 18358
rect 26238 18320 26240 18329
rect 26292 18320 26294 18329
rect 26238 18255 26294 18264
rect 26344 16833 26372 19110
rect 26424 18692 26476 18698
rect 26424 18634 26476 18640
rect 26330 16824 26386 16833
rect 26330 16759 26386 16768
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26146 15056 26202 15065
rect 26146 14991 26202 15000
rect 26160 9178 26188 14991
rect 26332 11620 26384 11626
rect 26332 11562 26384 11568
rect 26240 10532 26292 10538
rect 26240 10474 26292 10480
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 26160 8634 26188 8978
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 26252 8090 26280 10474
rect 26344 9466 26372 11562
rect 26436 10441 26464 18634
rect 26516 11280 26568 11286
rect 26516 11222 26568 11228
rect 26422 10432 26478 10441
rect 26422 10367 26478 10376
rect 26344 9438 26464 9466
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26344 8945 26372 9318
rect 26330 8936 26386 8945
rect 26330 8871 26386 8880
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26252 6916 26280 8026
rect 26160 6888 26280 6916
rect 26160 2922 26188 6888
rect 26436 6866 26464 9438
rect 26424 6860 26476 6866
rect 26424 6802 26476 6808
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26344 5817 26372 6054
rect 26330 5808 26386 5817
rect 26330 5743 26386 5752
rect 26240 5568 26292 5574
rect 26240 5510 26292 5516
rect 26252 5273 26280 5510
rect 26238 5264 26294 5273
rect 26238 5199 26294 5208
rect 26332 5024 26384 5030
rect 26238 4992 26294 5001
rect 26332 4966 26384 4972
rect 26238 4927 26294 4936
rect 26252 4826 26280 4927
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 26344 4593 26372 4966
rect 26330 4584 26386 4593
rect 26330 4519 26386 4528
rect 26436 4162 26464 6802
rect 26344 4134 26464 4162
rect 26238 3904 26294 3913
rect 26238 3839 26294 3848
rect 26252 3738 26280 3839
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26344 3670 26372 4134
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26332 3664 26384 3670
rect 26332 3606 26384 3612
rect 26330 3224 26386 3233
rect 26330 3159 26332 3168
rect 26384 3159 26386 3168
rect 26332 3130 26384 3136
rect 26148 2916 26200 2922
rect 26148 2858 26200 2864
rect 26436 1873 26464 3878
rect 26528 2553 26556 11222
rect 26608 6248 26660 6254
rect 26608 6190 26660 6196
rect 26620 3097 26648 6190
rect 26700 5296 26752 5302
rect 26700 5238 26752 5244
rect 26606 3088 26662 3097
rect 26606 3023 26662 3032
rect 26514 2544 26570 2553
rect 26514 2479 26570 2488
rect 26422 1864 26478 1873
rect 26422 1799 26478 1808
rect 26436 598 26556 626
rect 22926 439 22982 448
rect 23386 0 23442 480
rect 23938 0 23994 480
rect 24398 0 24454 480
rect 24950 0 25006 480
rect 25502 0 25558 480
rect 26054 0 26110 480
rect 26436 377 26464 598
rect 26528 480 26556 598
rect 26422 368 26478 377
rect 26422 303 26478 312
rect 26514 0 26570 480
rect 26712 377 26740 5238
rect 27066 640 27122 649
rect 27066 575 27122 584
rect 27356 598 27660 626
rect 27080 480 27108 575
rect 26698 368 26754 377
rect 26698 303 26754 312
rect 27066 0 27122 480
rect 27356 241 27384 598
rect 27632 480 27660 598
rect 27342 232 27398 241
rect 27342 167 27398 176
rect 27618 0 27674 480
<< via2 >>
rect 21178 27648 21234 27704
rect 294 25880 350 25936
rect 1122 26968 1178 27024
rect 1398 26288 1454 26344
rect 1214 25744 1270 25800
rect 1582 25608 1638 25664
rect 1490 24928 1546 24984
rect 2134 26152 2190 26208
rect 1766 24928 1822 24984
rect 1582 24248 1638 24304
rect 1398 18808 1454 18864
rect 1398 16768 1454 16824
rect 1398 15988 1400 16008
rect 1400 15988 1452 16008
rect 1452 15988 1454 16008
rect 1398 15952 1454 15988
rect 1398 15564 1454 15600
rect 1398 15544 1400 15564
rect 1400 15544 1452 15564
rect 1452 15544 1454 15564
rect 1398 12824 1454 12880
rect 1398 12688 1454 12744
rect 1674 21528 1730 21584
rect 1582 20304 1638 20360
rect 1858 20440 1914 20496
rect 1766 20304 1822 20360
rect 2686 26016 2742 26072
rect 2686 24928 2742 24984
rect 3054 24792 3110 24848
rect 3606 24792 3662 24848
rect 2502 24384 2558 24440
rect 3698 24112 3754 24168
rect 2594 23568 2650 23624
rect 2410 23160 2466 23216
rect 2042 19216 2098 19272
rect 1950 19080 2006 19136
rect 2226 17992 2282 18048
rect 2042 17176 2098 17232
rect 2134 16632 2190 16688
rect 1490 12280 1546 12336
rect 1398 11348 1454 11384
rect 1398 11328 1400 11348
rect 1400 11328 1452 11348
rect 1452 11328 1454 11348
rect 1582 11056 1638 11112
rect 1398 9152 1454 9208
rect 1490 5752 1546 5808
rect 1950 9696 2006 9752
rect 1674 8472 1730 8528
rect 1766 6704 1822 6760
rect 2410 22208 2466 22264
rect 2686 22888 2742 22944
rect 2594 21120 2650 21176
rect 2410 20304 2466 20360
rect 2870 20576 2926 20632
rect 2502 20032 2558 20088
rect 2594 17856 2650 17912
rect 3054 22480 3110 22536
rect 3054 20596 3110 20632
rect 3054 20576 3056 20596
rect 3056 20576 3108 20596
rect 3108 20576 3110 20596
rect 2962 19080 3018 19136
rect 2870 18708 2872 18728
rect 2872 18708 2924 18728
rect 2924 18708 2926 18728
rect 2870 18672 2926 18708
rect 2778 17992 2834 18048
rect 2502 17720 2558 17776
rect 2870 16496 2926 16552
rect 2502 15680 2558 15736
rect 2134 11192 2190 11248
rect 2778 13504 2834 13560
rect 2502 12316 2504 12336
rect 2504 12316 2556 12336
rect 2556 12316 2558 12336
rect 2502 12280 2558 12316
rect 2870 12960 2926 13016
rect 2870 12552 2926 12608
rect 3054 17856 3110 17912
rect 3606 23024 3662 23080
rect 3330 20884 3332 20904
rect 3332 20884 3384 20904
rect 3384 20884 3386 20904
rect 3330 20848 3386 20884
rect 3238 19896 3294 19952
rect 3238 18128 3294 18184
rect 3146 17040 3202 17096
rect 3146 13368 3202 13424
rect 3422 18944 3478 19000
rect 3698 20712 3754 20768
rect 3698 20576 3754 20632
rect 3514 17876 3570 17912
rect 3514 17856 3516 17876
rect 3516 17856 3568 17876
rect 3568 17856 3570 17876
rect 4158 23432 4214 23488
rect 4066 21256 4122 21312
rect 4158 21120 4214 21176
rect 3974 20032 4030 20088
rect 3790 18944 3846 19000
rect 3790 18672 3846 18728
rect 3422 15408 3478 15464
rect 3238 12960 3294 13016
rect 2962 12144 3018 12200
rect 2962 11228 2964 11248
rect 2964 11228 3016 11248
rect 3016 11228 3018 11248
rect 2962 11192 3018 11228
rect 3330 12552 3386 12608
rect 3146 11872 3202 11928
rect 3054 10920 3110 10976
rect 2410 9968 2466 10024
rect 1582 3984 1638 4040
rect 1398 720 1454 776
rect 2134 7520 2190 7576
rect 2042 4664 2098 4720
rect 2134 4276 2190 4312
rect 2134 4256 2136 4276
rect 2136 4256 2188 4276
rect 2188 4256 2190 4276
rect 3054 10240 3110 10296
rect 2870 10104 2926 10160
rect 2778 9288 2834 9344
rect 2686 9016 2742 9072
rect 2318 7928 2374 7984
rect 2962 9424 3018 9480
rect 2134 1264 2190 1320
rect 2502 6840 2558 6896
rect 2870 8064 2926 8120
rect 3606 16904 3662 16960
rect 3606 15000 3662 15056
rect 3514 11736 3570 11792
rect 3238 10648 3294 10704
rect 3146 8336 3202 8392
rect 2778 5616 2834 5672
rect 3146 6296 3202 6352
rect 2962 5652 2964 5672
rect 2964 5652 3016 5672
rect 3016 5652 3018 5672
rect 2962 5616 3018 5652
rect 2962 4800 3018 4856
rect 2502 2796 2504 2816
rect 2504 2796 2556 2816
rect 2556 2796 2558 2816
rect 2502 2760 2558 2796
rect 2870 3848 2926 3904
rect 2962 2388 2964 2408
rect 2964 2388 3016 2408
rect 3016 2388 3018 2408
rect 2962 2352 3018 2388
rect 3514 9424 3570 9480
rect 3330 9016 3386 9072
rect 3514 7692 3516 7712
rect 3516 7692 3568 7712
rect 3568 7692 3570 7712
rect 3514 7656 3570 7692
rect 3238 3712 3294 3768
rect 3422 3440 3478 3496
rect 3146 1944 3202 2000
rect 3422 2508 3478 2544
rect 3422 2488 3424 2508
rect 3424 2488 3476 2508
rect 3476 2488 3478 2508
rect 4158 19252 4160 19272
rect 4160 19252 4212 19272
rect 4212 19252 4214 19272
rect 4158 19216 4214 19252
rect 4066 18264 4122 18320
rect 5814 25200 5870 25256
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4526 21528 4582 21584
rect 4434 20848 4490 20904
rect 4066 16632 4122 16688
rect 3790 13912 3846 13968
rect 4250 15952 4306 16008
rect 4342 14592 4398 14648
rect 4158 13776 4214 13832
rect 3882 12552 3938 12608
rect 3790 9696 3846 9752
rect 3790 9424 3846 9480
rect 4066 13096 4122 13152
rect 4250 13640 4306 13696
rect 4342 13268 4344 13288
rect 4344 13268 4396 13288
rect 4396 13268 4398 13288
rect 4342 13232 4398 13268
rect 4066 12280 4122 12336
rect 4434 12552 4490 12608
rect 4434 9152 4490 9208
rect 4066 8064 4122 8120
rect 3882 5208 3938 5264
rect 4158 5888 4214 5944
rect 3974 4936 4030 4992
rect 3882 4392 3938 4448
rect 3698 2216 3754 2272
rect 3790 1536 3846 1592
rect 3698 992 3754 1048
rect 4342 4120 4398 4176
rect 4710 21800 4766 21856
rect 4802 17060 4858 17096
rect 4802 17040 4804 17060
rect 4804 17040 4856 17060
rect 4856 17040 4858 17060
rect 4618 13504 4674 13560
rect 4618 11600 4674 11656
rect 4986 21956 5042 21992
rect 4986 21936 4988 21956
rect 4988 21936 5040 21956
rect 5040 21936 5042 21956
rect 5446 23432 5502 23488
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5630 23316 5686 23352
rect 5630 23296 5632 23316
rect 5632 23296 5684 23316
rect 5684 23296 5686 23316
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5722 22380 5724 22400
rect 5724 22380 5776 22400
rect 5776 22380 5778 22400
rect 5722 22344 5778 22380
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5998 21412 6054 21448
rect 5998 21392 6000 21412
rect 6000 21392 6052 21412
rect 6052 21392 6054 21412
rect 5630 20848 5686 20904
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5630 20440 5686 20496
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5262 19216 5318 19272
rect 5998 19080 6054 19136
rect 5998 18808 6054 18864
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5630 17040 5686 17096
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 4802 13368 4858 13424
rect 4802 12552 4858 12608
rect 4802 11872 4858 11928
rect 4710 11464 4766 11520
rect 5170 14764 5172 14784
rect 5172 14764 5224 14784
rect 5224 14764 5226 14784
rect 5170 14728 5226 14764
rect 4986 10784 5042 10840
rect 4618 9152 4674 9208
rect 4618 5072 4674 5128
rect 4894 10376 4950 10432
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5446 13368 5502 13424
rect 5262 12824 5318 12880
rect 5170 11600 5226 11656
rect 5262 10920 5318 10976
rect 5170 10648 5226 10704
rect 5262 10512 5318 10568
rect 5262 9596 5264 9616
rect 5264 9596 5316 9616
rect 5316 9596 5318 9616
rect 5262 9560 5318 9596
rect 5262 9016 5318 9072
rect 4894 7792 4950 7848
rect 4802 7384 4858 7440
rect 4986 7112 5042 7168
rect 5170 6976 5226 7032
rect 5078 6840 5134 6896
rect 4802 6160 4858 6216
rect 5078 6296 5134 6352
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 6550 23568 6606 23624
rect 6458 23024 6514 23080
rect 6366 22208 6422 22264
rect 6550 22380 6552 22400
rect 6552 22380 6604 22400
rect 6604 22380 6606 22400
rect 6550 22344 6606 22380
rect 6458 22072 6514 22128
rect 7194 25064 7250 25120
rect 7010 24656 7066 24712
rect 6734 23704 6790 23760
rect 6642 21936 6698 21992
rect 6642 18128 6698 18184
rect 6642 17720 6698 17776
rect 6642 17312 6698 17368
rect 7010 23976 7066 24032
rect 6826 23160 6882 23216
rect 7102 22380 7104 22400
rect 7104 22380 7156 22400
rect 7156 22380 7158 22400
rect 7102 22344 7158 22380
rect 7470 24112 7526 24168
rect 7654 25200 7710 25256
rect 6918 21936 6974 21992
rect 7010 21256 7066 21312
rect 7010 20984 7066 21040
rect 7194 20984 7250 21040
rect 7102 20848 7158 20904
rect 6826 19216 6882 19272
rect 7010 19216 7066 19272
rect 7010 18808 7066 18864
rect 7194 20032 7250 20088
rect 7378 20032 7434 20088
rect 7194 19488 7250 19544
rect 7194 18944 7250 19000
rect 6826 17720 6882 17776
rect 6090 15308 6092 15328
rect 6092 15308 6144 15328
rect 6144 15308 6146 15328
rect 6090 15272 6146 15308
rect 6182 14728 6238 14784
rect 6090 13504 6146 13560
rect 5998 12960 6054 13016
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5906 11348 5962 11384
rect 5906 11328 5908 11348
rect 5908 11328 5960 11348
rect 5960 11328 5962 11348
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5538 10240 5594 10296
rect 5722 10004 5724 10024
rect 5724 10004 5776 10024
rect 5776 10004 5778 10024
rect 5722 9968 5778 10004
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5446 8472 5502 8528
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5538 7928 5594 7984
rect 5446 7656 5502 7712
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5446 6704 5502 6760
rect 5170 5752 5226 5808
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5906 5752 5962 5808
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5078 4820 5134 4856
rect 5078 4800 5080 4820
rect 5080 4800 5132 4820
rect 5132 4800 5134 4820
rect 4986 4256 5042 4312
rect 4434 3576 4490 3632
rect 4894 3596 4950 3632
rect 4894 3576 4896 3596
rect 4896 3576 4948 3596
rect 4948 3576 4950 3596
rect 4434 1536 4490 1592
rect 3974 40 4030 96
rect 5262 4800 5318 4856
rect 6366 14592 6422 14648
rect 6918 16788 6974 16824
rect 6918 16768 6920 16788
rect 6920 16768 6972 16788
rect 6972 16768 6974 16788
rect 6918 16632 6974 16688
rect 6642 16360 6698 16416
rect 6734 15700 6790 15736
rect 6734 15680 6736 15700
rect 6736 15680 6788 15700
rect 6788 15680 6790 15700
rect 6642 15136 6698 15192
rect 6734 14728 6790 14784
rect 6734 14320 6790 14376
rect 6642 14068 6698 14104
rect 6642 14048 6644 14068
rect 6644 14048 6696 14068
rect 6696 14048 6698 14068
rect 6642 13812 6644 13832
rect 6644 13812 6696 13832
rect 6696 13812 6698 13832
rect 6642 13776 6698 13812
rect 6274 10784 6330 10840
rect 6642 11736 6698 11792
rect 6642 11328 6698 11384
rect 6642 10920 6698 10976
rect 6366 9424 6422 9480
rect 5262 3848 5318 3904
rect 5354 3032 5410 3088
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5998 4020 6000 4040
rect 6000 4020 6052 4040
rect 6052 4020 6054 4040
rect 5998 3984 6054 4020
rect 6550 9324 6552 9344
rect 6552 9324 6604 9344
rect 6604 9324 6606 9344
rect 6550 9288 6606 9324
rect 6366 5208 6422 5264
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6918 15000 6974 15056
rect 7102 15816 7158 15872
rect 7194 14220 7196 14240
rect 7196 14220 7248 14240
rect 7248 14220 7250 14240
rect 7194 14184 7250 14220
rect 7562 23860 7618 23896
rect 7562 23840 7564 23860
rect 7564 23840 7616 23860
rect 7616 23840 7618 23860
rect 7378 18536 7434 18592
rect 7838 22072 7894 22128
rect 7654 19216 7710 19272
rect 7746 18808 7802 18864
rect 7838 17992 7894 18048
rect 7378 15816 7434 15872
rect 7378 15408 7434 15464
rect 7562 15272 7618 15328
rect 7010 10512 7066 10568
rect 7102 10240 7158 10296
rect 6826 8744 6882 8800
rect 6918 8628 6974 8664
rect 6918 8608 6920 8628
rect 6920 8608 6972 8628
rect 6972 8608 6974 8628
rect 6734 8200 6790 8256
rect 6642 8064 6698 8120
rect 6642 7656 6698 7712
rect 6458 4528 6514 4584
rect 6366 4120 6422 4176
rect 6826 7520 6882 7576
rect 6918 6452 6974 6488
rect 6918 6432 6920 6452
rect 6920 6432 6972 6452
rect 6972 6432 6974 6452
rect 6918 5788 6920 5808
rect 6920 5788 6972 5808
rect 6972 5788 6974 5808
rect 6918 5752 6974 5788
rect 7010 4276 7066 4312
rect 7010 4256 7012 4276
rect 7012 4256 7064 4276
rect 7064 4256 7066 4276
rect 6550 3848 6606 3904
rect 5906 2372 5962 2408
rect 5906 2352 5908 2372
rect 5908 2352 5960 2372
rect 5960 2352 5962 2372
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7010 3984 7066 4040
rect 6918 3032 6974 3088
rect 7378 9832 7434 9888
rect 8022 24268 8078 24304
rect 8022 24248 8024 24268
rect 8024 24248 8076 24268
rect 8076 24248 8078 24268
rect 8114 23296 8170 23352
rect 8022 23024 8078 23080
rect 8114 22888 8170 22944
rect 8022 21936 8078 21992
rect 8206 22616 8262 22672
rect 8574 23196 8576 23216
rect 8576 23196 8628 23216
rect 8628 23196 8630 23216
rect 8574 23160 8630 23196
rect 8482 22752 8538 22808
rect 8758 24112 8814 24168
rect 8850 23160 8906 23216
rect 8298 21664 8354 21720
rect 8206 20848 8262 20904
rect 8390 19760 8446 19816
rect 8298 19352 8354 19408
rect 8666 22344 8722 22400
rect 8114 16904 8170 16960
rect 7838 15136 7894 15192
rect 8298 16496 8354 16552
rect 8482 18808 8538 18864
rect 8574 17992 8630 18048
rect 8390 14864 8446 14920
rect 7930 13368 7986 13424
rect 7930 13096 7986 13152
rect 8574 14456 8630 14512
rect 7838 11600 7894 11656
rect 7654 9424 7710 9480
rect 7654 8880 7710 8936
rect 7562 8744 7618 8800
rect 7378 6724 7434 6760
rect 7378 6704 7380 6724
rect 7380 6704 7432 6724
rect 7432 6704 7434 6724
rect 7746 4528 7802 4584
rect 7654 3576 7710 3632
rect 7746 3304 7802 3360
rect 7654 2896 7710 2952
rect 7378 2488 7434 2544
rect 7470 2216 7526 2272
rect 7562 2080 7618 2136
rect 8114 12416 8170 12472
rect 8206 12144 8262 12200
rect 8114 11736 8170 11792
rect 8022 11056 8078 11112
rect 8298 11464 8354 11520
rect 8298 10124 8354 10160
rect 8298 10104 8300 10124
rect 8300 10104 8352 10124
rect 8352 10104 8354 10124
rect 7930 9016 7986 9072
rect 7930 6976 7986 7032
rect 7930 6568 7986 6624
rect 8298 9152 8354 9208
rect 8206 8336 8262 8392
rect 8298 7792 8354 7848
rect 8482 11892 8538 11928
rect 8482 11872 8484 11892
rect 8484 11872 8536 11892
rect 8536 11872 8538 11892
rect 9402 25336 9458 25392
rect 9310 24384 9366 24440
rect 9310 22480 9366 22536
rect 8850 21664 8906 21720
rect 8850 19352 8906 19408
rect 8942 18264 8998 18320
rect 8942 17992 8998 18048
rect 8850 16904 8906 16960
rect 8850 14728 8906 14784
rect 8758 12144 8814 12200
rect 9218 22208 9274 22264
rect 9218 20576 9274 20632
rect 9586 24928 9642 24984
rect 10138 26424 10194 26480
rect 9954 26288 10010 26344
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10138 25472 10194 25528
rect 9770 24792 9826 24848
rect 9494 24520 9550 24576
rect 9586 24248 9642 24304
rect 9494 21800 9550 21856
rect 9402 21528 9458 21584
rect 9402 20712 9458 20768
rect 9862 23296 9918 23352
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 9862 21956 9918 21992
rect 9862 21936 9864 21956
rect 9864 21936 9916 21956
rect 9916 21936 9918 21956
rect 10046 21800 10102 21856
rect 9494 20440 9550 20496
rect 9678 20884 9680 20904
rect 9680 20884 9732 20904
rect 9732 20884 9734 20904
rect 9678 20848 9734 20884
rect 9770 20712 9826 20768
rect 9678 20204 9680 20224
rect 9680 20204 9732 20224
rect 9732 20204 9734 20224
rect 9678 20168 9734 20204
rect 9770 20032 9826 20088
rect 9494 18944 9550 19000
rect 9954 20032 10010 20088
rect 9770 19760 9826 19816
rect 9770 19080 9826 19136
rect 9034 12960 9090 13016
rect 9310 16360 9366 16416
rect 9402 15680 9458 15736
rect 9034 12300 9090 12336
rect 9034 12280 9036 12300
rect 9036 12280 9088 12300
rect 9088 12280 9090 12300
rect 8942 11620 8998 11656
rect 8942 11600 8944 11620
rect 8944 11600 8996 11620
rect 8996 11600 8998 11620
rect 8850 11464 8906 11520
rect 8666 9560 8722 9616
rect 8482 8200 8538 8256
rect 8482 8064 8538 8120
rect 8758 8880 8814 8936
rect 8666 7112 8722 7168
rect 8758 6840 8814 6896
rect 8666 6704 8722 6760
rect 8574 6160 8630 6216
rect 8666 5888 8722 5944
rect 8758 5092 8814 5128
rect 8758 5072 8760 5092
rect 8760 5072 8812 5092
rect 8812 5072 8814 5092
rect 8942 6704 8998 6760
rect 8114 3984 8170 4040
rect 8022 3304 8078 3360
rect 7930 1672 7986 1728
rect 7378 856 7434 912
rect 8758 4664 8814 4720
rect 9034 3984 9090 4040
rect 8942 1808 8998 1864
rect 9586 15680 9642 15736
rect 9494 15000 9550 15056
rect 9862 17584 9918 17640
rect 9862 16088 9918 16144
rect 9770 15952 9826 16008
rect 9770 15136 9826 15192
rect 9954 15544 10010 15600
rect 9954 15408 10010 15464
rect 9862 14320 9918 14376
rect 9494 14048 9550 14104
rect 9678 13912 9734 13968
rect 9770 13776 9826 13832
rect 9678 13640 9734 13696
rect 9678 12960 9734 13016
rect 9218 9832 9274 9888
rect 9402 9968 9458 10024
rect 9678 12416 9734 12472
rect 9678 12316 9680 12336
rect 9680 12316 9732 12336
rect 9732 12316 9734 12336
rect 9678 12280 9734 12316
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10782 23840 10838 23896
rect 11150 25744 11206 25800
rect 11150 25200 11206 25256
rect 11058 24112 11114 24168
rect 11242 22208 11298 22264
rect 10966 22072 11022 22128
rect 10690 21528 10746 21584
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 11150 21936 11206 21992
rect 11058 21836 11060 21856
rect 11060 21836 11112 21856
rect 11112 21836 11114 21856
rect 11058 21800 11114 21836
rect 11058 21664 11114 21720
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10874 19488 10930 19544
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10322 17756 10324 17776
rect 10324 17756 10376 17776
rect 10376 17756 10378 17776
rect 10322 17720 10378 17756
rect 11242 20576 11298 20632
rect 11334 20168 11390 20224
rect 11242 19216 11298 19272
rect 11334 19116 11336 19136
rect 11336 19116 11388 19136
rect 11388 19116 11390 19136
rect 11150 18400 11206 18456
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10322 16632 10378 16688
rect 10874 16632 10930 16688
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10874 15680 10930 15736
rect 10046 14592 10102 14648
rect 10046 14068 10102 14104
rect 10046 14048 10048 14068
rect 10048 14048 10100 14068
rect 10100 14048 10102 14068
rect 10046 13524 10102 13560
rect 10046 13504 10048 13524
rect 10048 13504 10100 13524
rect 10100 13504 10102 13524
rect 9862 12416 9918 12472
rect 9770 11328 9826 11384
rect 9770 10376 9826 10432
rect 9494 9832 9550 9888
rect 9218 7404 9274 7440
rect 9218 7384 9220 7404
rect 9220 7384 9272 7404
rect 9272 7384 9274 7404
rect 9586 7520 9642 7576
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 11334 19080 11390 19116
rect 11334 18128 11390 18184
rect 11334 17312 11390 17368
rect 10690 13232 10746 13288
rect 10598 12724 10600 12744
rect 10600 12724 10652 12744
rect 10652 12724 10654 12744
rect 10598 12688 10654 12724
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 11058 14728 11114 14784
rect 11058 13912 11114 13968
rect 11058 13504 11114 13560
rect 10690 11772 10692 11792
rect 10692 11772 10744 11792
rect 10744 11772 10746 11792
rect 10690 11736 10746 11772
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10322 11056 10378 11112
rect 10782 11464 10838 11520
rect 11794 24112 11850 24168
rect 12254 24656 12310 24712
rect 11886 23976 11942 24032
rect 11794 23568 11850 23624
rect 11978 23568 12034 23624
rect 11702 22208 11758 22264
rect 11702 20884 11704 20904
rect 11704 20884 11756 20904
rect 11756 20884 11758 20904
rect 11702 20848 11758 20884
rect 12530 24112 12586 24168
rect 13082 24812 13138 24848
rect 13082 24792 13084 24812
rect 13084 24792 13136 24812
rect 13136 24792 13138 24812
rect 12162 22516 12164 22536
rect 12164 22516 12216 22536
rect 12216 22516 12218 22536
rect 12162 22480 12218 22516
rect 12806 23432 12862 23488
rect 12530 22480 12586 22536
rect 12346 22072 12402 22128
rect 11886 20168 11942 20224
rect 11610 18264 11666 18320
rect 11702 13912 11758 13968
rect 11242 12588 11244 12608
rect 11244 12588 11296 12608
rect 11296 12588 11298 12608
rect 11242 12552 11298 12588
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10138 10240 10194 10296
rect 9862 9016 9918 9072
rect 9770 7384 9826 7440
rect 9770 6160 9826 6216
rect 9678 5480 9734 5536
rect 9862 4800 9918 4856
rect 9586 4392 9642 4448
rect 9494 4256 9550 4312
rect 10690 9832 10746 9888
rect 10138 9288 10194 9344
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10414 7520 10470 7576
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 11334 10412 11336 10432
rect 11336 10412 11388 10432
rect 11388 10412 11390 10432
rect 11334 10376 11390 10412
rect 10874 9596 10876 9616
rect 10876 9596 10928 9616
rect 10928 9596 10930 9616
rect 10874 9560 10930 9596
rect 10782 7792 10838 7848
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10046 4700 10048 4720
rect 10048 4700 10100 4720
rect 10100 4700 10102 4720
rect 10046 4664 10102 4700
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10782 4800 10838 4856
rect 11058 9424 11114 9480
rect 11426 9696 11482 9752
rect 11150 8234 11206 8290
rect 11058 7928 11114 7984
rect 11058 6568 11114 6624
rect 9494 3460 9550 3496
rect 9494 3440 9496 3460
rect 9496 3440 9548 3460
rect 9548 3440 9550 3460
rect 9770 3440 9826 3496
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10046 3712 10102 3768
rect 10782 3304 10838 3360
rect 10138 2896 10194 2952
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10782 2760 10838 2816
rect 10690 2624 10746 2680
rect 10322 2508 10378 2544
rect 10322 2488 10324 2508
rect 10324 2488 10376 2508
rect 10376 2488 10378 2508
rect 10506 2216 10562 2272
rect 10690 2216 10746 2272
rect 11978 19488 12034 19544
rect 12714 20984 12770 21040
rect 12622 20748 12624 20768
rect 12624 20748 12676 20768
rect 12676 20748 12678 20768
rect 12622 20712 12678 20748
rect 12346 19796 12348 19816
rect 12348 19796 12400 19816
rect 12400 19796 12402 19816
rect 12346 19760 12402 19796
rect 12622 20304 12678 20360
rect 12070 19080 12126 19136
rect 11978 18944 12034 19000
rect 11886 16632 11942 16688
rect 12162 17212 12164 17232
rect 12164 17212 12216 17232
rect 12216 17212 12218 17232
rect 12162 17176 12218 17212
rect 12070 17040 12126 17096
rect 12438 18944 12494 19000
rect 13082 22208 13138 22264
rect 12438 18672 12494 18728
rect 12622 18672 12678 18728
rect 12622 18536 12678 18592
rect 12530 17992 12586 18048
rect 12530 17720 12586 17776
rect 12438 16904 12494 16960
rect 12162 16496 12218 16552
rect 11334 6296 11390 6352
rect 11150 1944 11206 2000
rect 11610 5752 11666 5808
rect 11610 5616 11666 5672
rect 12070 10240 12126 10296
rect 11886 7656 11942 7712
rect 11794 6432 11850 6488
rect 11794 5616 11850 5672
rect 11702 5208 11758 5264
rect 11794 3984 11850 4040
rect 11610 3596 11666 3632
rect 11610 3576 11612 3596
rect 11612 3576 11664 3596
rect 11664 3576 11666 3596
rect 11334 1944 11390 2000
rect 12530 16124 12532 16144
rect 12532 16124 12584 16144
rect 12584 16124 12586 16144
rect 12530 16088 12586 16124
rect 12806 17856 12862 17912
rect 12714 16088 12770 16144
rect 12714 15136 12770 15192
rect 13358 26016 13414 26072
rect 13726 25336 13782 25392
rect 13450 23604 13452 23624
rect 13452 23604 13504 23624
rect 13504 23604 13506 23624
rect 13450 23568 13506 23604
rect 14002 24692 14004 24712
rect 14004 24692 14056 24712
rect 14056 24692 14058 24712
rect 14002 24656 14058 24692
rect 14370 24928 14426 24984
rect 13910 24248 13966 24304
rect 13174 20304 13230 20360
rect 13266 18944 13322 19000
rect 13266 18400 13322 18456
rect 13818 22752 13874 22808
rect 13634 21528 13690 21584
rect 13542 20304 13598 20360
rect 13174 17720 13230 17776
rect 13634 19116 13636 19136
rect 13636 19116 13688 19136
rect 13688 19116 13690 19136
rect 13634 19080 13690 19116
rect 13634 17856 13690 17912
rect 12714 14864 12770 14920
rect 12530 12280 12586 12336
rect 12530 12008 12586 12064
rect 12346 11600 12402 11656
rect 12438 8200 12494 8256
rect 12254 7268 12310 7304
rect 12254 7248 12256 7268
rect 12256 7248 12308 7268
rect 12308 7248 12310 7268
rect 12438 6704 12494 6760
rect 12162 4664 12218 4720
rect 12438 5888 12494 5944
rect 12438 4936 12494 4992
rect 12438 4664 12494 4720
rect 12622 4664 12678 4720
rect 12530 4256 12586 4312
rect 12162 3032 12218 3088
rect 13174 14728 13230 14784
rect 13082 14184 13138 14240
rect 13634 17584 13690 17640
rect 13634 16224 13690 16280
rect 13726 15680 13782 15736
rect 13450 14320 13506 14376
rect 13358 14184 13414 14240
rect 13174 8880 13230 8936
rect 13082 8336 13138 8392
rect 12806 5480 12862 5536
rect 13174 7656 13230 7712
rect 12990 5344 13046 5400
rect 13082 4800 13138 4856
rect 12898 3848 12954 3904
rect 12530 2760 12586 2816
rect 12438 2488 12494 2544
rect 13266 2252 13268 2272
rect 13268 2252 13320 2272
rect 13320 2252 13322 2272
rect 13266 2216 13322 2252
rect 12898 1400 12954 1456
rect 13542 7928 13598 7984
rect 13726 13368 13782 13424
rect 14370 24112 14426 24168
rect 14278 23704 14334 23760
rect 14278 19080 14334 19136
rect 14554 24268 14610 24304
rect 14554 24248 14556 24268
rect 14556 24248 14608 24268
rect 14608 24248 14610 24268
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14830 24792 14886 24848
rect 15566 25336 15622 25392
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15750 25880 15806 25936
rect 15106 23044 15162 23080
rect 15106 23024 15108 23044
rect 15108 23024 15160 23044
rect 15160 23024 15162 23044
rect 15382 23296 15438 23352
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15290 22072 15346 22128
rect 15106 21972 15108 21992
rect 15108 21972 15160 21992
rect 15160 21972 15162 21992
rect 15106 21936 15162 21972
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15382 21684 15438 21720
rect 15382 21664 15384 21684
rect 15384 21664 15436 21684
rect 15436 21664 15438 21684
rect 14646 21528 14702 21584
rect 14554 21392 14610 21448
rect 14830 21428 14832 21448
rect 14832 21428 14884 21448
rect 14884 21428 14886 21448
rect 14830 21392 14886 21428
rect 15014 21140 15070 21176
rect 15014 21120 15016 21140
rect 15016 21120 15068 21140
rect 15068 21120 15070 21140
rect 15382 21120 15438 21176
rect 14738 20576 14794 20632
rect 15290 20848 15346 20904
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14646 20440 14702 20496
rect 16118 26288 16174 26344
rect 16026 25880 16082 25936
rect 16026 24928 16082 24984
rect 16026 24384 16082 24440
rect 15750 23860 15806 23896
rect 15750 23840 15752 23860
rect 15752 23840 15804 23860
rect 15804 23840 15806 23860
rect 15658 23704 15714 23760
rect 15658 22072 15714 22128
rect 14738 19896 14794 19952
rect 14646 19388 14648 19408
rect 14648 19388 14700 19408
rect 14700 19388 14702 19408
rect 14646 19352 14702 19388
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15382 19488 15438 19544
rect 15382 19216 15438 19272
rect 15106 18828 15162 18864
rect 15106 18808 15108 18828
rect 15108 18808 15160 18828
rect 15160 18808 15162 18828
rect 14830 18672 14886 18728
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14738 18400 14794 18456
rect 15382 18400 15438 18456
rect 14186 16360 14242 16416
rect 14094 15272 14150 15328
rect 14002 14320 14058 14376
rect 13910 13096 13966 13152
rect 13818 9288 13874 9344
rect 14370 15816 14426 15872
rect 14370 12824 14426 12880
rect 13910 8880 13966 8936
rect 14186 11600 14242 11656
rect 14094 9696 14150 9752
rect 13634 3460 13690 3496
rect 13634 3440 13636 3460
rect 13636 3440 13688 3460
rect 13688 3440 13690 3460
rect 13634 1536 13690 1592
rect 4434 312 4490 368
rect 14278 9288 14334 9344
rect 14738 17448 14794 17504
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14646 15136 14702 15192
rect 14646 14048 14702 14104
rect 14738 13776 14794 13832
rect 14738 12824 14794 12880
rect 14646 10804 14702 10840
rect 14646 10784 14648 10804
rect 14648 10784 14700 10804
rect 14700 10784 14702 10804
rect 14002 4936 14058 4992
rect 14370 8744 14426 8800
rect 14554 8744 14610 8800
rect 14646 8608 14702 8664
rect 14370 6840 14426 6896
rect 13910 3712 13966 3768
rect 14186 3712 14242 3768
rect 13818 3576 13874 3632
rect 13910 3440 13966 3496
rect 14094 3476 14096 3496
rect 14096 3476 14148 3496
rect 14148 3476 14150 3496
rect 14094 3440 14150 3476
rect 14922 17176 14978 17232
rect 15014 16904 15070 16960
rect 15474 16768 15530 16824
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15382 16224 15438 16280
rect 15474 16088 15530 16144
rect 14922 15816 14978 15872
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15198 15000 15254 15056
rect 15382 14764 15384 14784
rect 15384 14764 15436 14784
rect 15436 14764 15438 14784
rect 15382 14728 15438 14764
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15106 12552 15162 12608
rect 14922 12180 14924 12200
rect 14924 12180 14976 12200
rect 14976 12180 14978 12200
rect 14922 12144 14978 12180
rect 15106 12144 15162 12200
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14830 11464 14886 11520
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14922 7812 14978 7848
rect 14922 7792 14924 7812
rect 14924 7792 14976 7812
rect 14976 7792 14978 7812
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15658 20304 15714 20360
rect 15750 19896 15806 19952
rect 15658 15680 15714 15736
rect 15658 15272 15714 15328
rect 15842 18672 15898 18728
rect 16210 23468 16212 23488
rect 16212 23468 16264 23488
rect 16264 23468 16266 23488
rect 16210 23432 16266 23468
rect 17314 26424 17370 26480
rect 16486 24520 16542 24576
rect 17314 25200 17370 25256
rect 16762 24792 16818 24848
rect 16670 23840 16726 23896
rect 16394 21800 16450 21856
rect 16302 21392 16358 21448
rect 16486 21256 16542 21312
rect 16394 21120 16450 21176
rect 16210 20168 16266 20224
rect 16118 19372 16174 19408
rect 16118 19352 16120 19372
rect 16120 19352 16172 19372
rect 16172 19352 16174 19372
rect 15842 17720 15898 17776
rect 16026 17312 16082 17368
rect 15934 17212 15936 17232
rect 15936 17212 15988 17232
rect 15988 17212 15990 17232
rect 15934 17176 15990 17212
rect 15842 15408 15898 15464
rect 15934 13404 15936 13424
rect 15936 13404 15988 13424
rect 15988 13404 15990 13424
rect 15934 13368 15990 13404
rect 15658 12144 15714 12200
rect 15658 11600 15714 11656
rect 15474 11092 15476 11112
rect 15476 11092 15528 11112
rect 15528 11092 15530 11112
rect 15474 11056 15530 11092
rect 15474 10920 15530 10976
rect 15566 9868 15568 9888
rect 15568 9868 15620 9888
rect 15620 9868 15622 9888
rect 15566 9832 15622 9868
rect 14922 6976 14978 7032
rect 15382 7148 15384 7168
rect 15384 7148 15436 7168
rect 15436 7148 15438 7168
rect 15382 7112 15438 7148
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14646 3596 14702 3632
rect 14646 3576 14648 3596
rect 14648 3576 14700 3596
rect 14700 3576 14702 3596
rect 15474 6296 15530 6352
rect 15474 3848 15530 3904
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14554 2896 14610 2952
rect 14646 2100 14702 2136
rect 14646 2080 14648 2100
rect 14648 2080 14700 2100
rect 14700 2080 14702 2100
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14554 1672 14610 1728
rect 14738 1672 14794 1728
rect 14462 1536 14518 1592
rect 14922 1400 14978 1456
rect 15106 1400 15162 1456
rect 15290 1128 15346 1184
rect 13726 176 13782 232
rect 16394 20304 16450 20360
rect 16210 18028 16212 18048
rect 16212 18028 16264 18048
rect 16264 18028 16266 18048
rect 16210 17992 16266 18028
rect 16854 23024 16910 23080
rect 16762 22888 16818 22944
rect 17590 23160 17646 23216
rect 17038 21936 17094 21992
rect 16210 15952 16266 16008
rect 16302 13932 16358 13968
rect 16302 13912 16304 13932
rect 16304 13912 16356 13932
rect 16356 13912 16358 13932
rect 17038 20984 17094 21040
rect 17314 20440 17370 20496
rect 16762 16496 16818 16552
rect 16762 15816 16818 15872
rect 16486 13232 16542 13288
rect 16946 19080 17002 19136
rect 17038 18672 17094 18728
rect 17130 18400 17186 18456
rect 16946 17584 17002 17640
rect 16854 15408 16910 15464
rect 16762 14320 16818 14376
rect 17038 16632 17094 16688
rect 16946 14884 17002 14920
rect 16946 14864 16948 14884
rect 16948 14864 17000 14884
rect 17000 14864 17002 14884
rect 17038 14456 17094 14512
rect 16946 14320 17002 14376
rect 16854 14048 16910 14104
rect 16762 13524 16818 13560
rect 16762 13504 16764 13524
rect 16764 13504 16816 13524
rect 16816 13504 16818 13524
rect 16762 13096 16818 13152
rect 16394 11600 16450 11656
rect 16394 10260 16450 10296
rect 16394 10240 16396 10260
rect 16396 10240 16448 10260
rect 16448 10240 16450 10260
rect 15750 8880 15806 8936
rect 16026 7928 16082 7984
rect 16210 8608 16266 8664
rect 16670 8508 16672 8528
rect 16672 8508 16724 8528
rect 16724 8508 16726 8528
rect 16670 8472 16726 8508
rect 16394 8336 16450 8392
rect 16118 7692 16120 7712
rect 16120 7692 16172 7712
rect 16172 7692 16174 7712
rect 16118 7656 16174 7692
rect 15750 7112 15806 7168
rect 16302 6160 16358 6216
rect 15658 4936 15714 4992
rect 15658 3712 15714 3768
rect 15750 1944 15806 2000
rect 15658 1808 15714 1864
rect 16486 6740 16488 6760
rect 16488 6740 16540 6760
rect 16540 6740 16542 6760
rect 16486 6704 16542 6740
rect 16486 5636 16542 5672
rect 16486 5616 16488 5636
rect 16488 5616 16540 5636
rect 16540 5616 16542 5636
rect 17130 10648 17186 10704
rect 17038 9696 17094 9752
rect 17222 9832 17278 9888
rect 17038 9016 17094 9072
rect 17682 23060 17684 23080
rect 17684 23060 17736 23080
rect 17736 23060 17738 23080
rect 17682 23024 17738 23060
rect 18326 24284 18328 24304
rect 18328 24284 18380 24304
rect 18380 24284 18382 24304
rect 18326 24248 18382 24284
rect 18142 24112 18198 24168
rect 17958 23568 18014 23624
rect 17866 20596 17922 20632
rect 17866 20576 17868 20596
rect 17868 20576 17920 20596
rect 17920 20576 17922 20596
rect 17590 17040 17646 17096
rect 17866 16088 17922 16144
rect 18234 22616 18290 22672
rect 18050 19216 18106 19272
rect 18142 17720 18198 17776
rect 18234 17312 18290 17368
rect 18142 16088 18198 16144
rect 17498 14728 17554 14784
rect 17866 14728 17922 14784
rect 18142 15272 18198 15328
rect 18602 23588 18658 23624
rect 18602 23568 18604 23588
rect 18604 23568 18656 23588
rect 18656 23568 18658 23588
rect 18602 23432 18658 23488
rect 18510 22208 18566 22264
rect 18510 20748 18512 20768
rect 18512 20748 18564 20768
rect 18564 20748 18566 20768
rect 18510 20712 18566 20748
rect 18602 18808 18658 18864
rect 18510 18536 18566 18592
rect 18970 25472 19026 25528
rect 19062 24656 19118 24712
rect 19338 26152 19394 26208
rect 19246 24384 19302 24440
rect 19154 23296 19210 23352
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20166 24928 20222 24984
rect 19338 23024 19394 23080
rect 19338 22924 19340 22944
rect 19340 22924 19392 22944
rect 19392 22924 19394 22944
rect 19338 22888 19394 22924
rect 19338 22652 19340 22672
rect 19340 22652 19392 22672
rect 19392 22652 19394 22672
rect 19338 22616 19394 22652
rect 19338 22516 19340 22536
rect 19340 22516 19392 22536
rect 19392 22516 19394 22536
rect 19338 22480 19394 22516
rect 19154 22208 19210 22264
rect 18970 20576 19026 20632
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 20074 23432 20130 23488
rect 19706 22652 19708 22672
rect 19708 22652 19760 22672
rect 19760 22652 19762 22672
rect 19706 22616 19762 22652
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19614 22108 19616 22128
rect 19616 22108 19668 22128
rect 19668 22108 19670 22128
rect 19614 22072 19670 22108
rect 19430 21256 19486 21312
rect 19338 20848 19394 20904
rect 18878 19352 18934 19408
rect 18970 18944 19026 19000
rect 18694 17856 18750 17912
rect 18602 17584 18658 17640
rect 18786 17448 18842 17504
rect 18326 15408 18382 15464
rect 18234 14184 18290 14240
rect 17774 11192 17830 11248
rect 17774 10512 17830 10568
rect 17406 9832 17462 9888
rect 17958 10140 17960 10160
rect 17960 10140 18012 10160
rect 18012 10140 18014 10160
rect 17958 10104 18014 10140
rect 17498 9560 17554 9616
rect 17314 9288 17370 9344
rect 17314 9016 17370 9072
rect 17406 8508 17408 8528
rect 17408 8508 17460 8528
rect 17460 8508 17462 8528
rect 17406 8472 17462 8508
rect 17406 7384 17462 7440
rect 16946 7248 17002 7304
rect 17222 5888 17278 5944
rect 16394 4256 16450 4312
rect 16486 3340 16488 3360
rect 16488 3340 16540 3360
rect 16540 3340 16542 3360
rect 16486 3304 16542 3340
rect 16670 2624 16726 2680
rect 16578 2488 16634 2544
rect 17038 4392 17094 4448
rect 17038 4256 17094 4312
rect 16854 3168 16910 3224
rect 15566 312 15622 368
rect 16394 448 16450 504
rect 17130 4120 17186 4176
rect 17130 3732 17186 3768
rect 17130 3712 17132 3732
rect 17132 3712 17184 3732
rect 17184 3712 17186 3732
rect 17314 5072 17370 5128
rect 17314 4120 17370 4176
rect 17406 2080 17462 2136
rect 18326 11736 18382 11792
rect 18786 16360 18842 16416
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19338 19624 19394 19680
rect 19062 16088 19118 16144
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 20074 18944 20130 19000
rect 19614 18808 19670 18864
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19522 17312 19578 17368
rect 19890 17312 19946 17368
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19522 16360 19578 16416
rect 19338 15952 19394 16008
rect 19062 15544 19118 15600
rect 18970 15308 18972 15328
rect 18972 15308 19024 15328
rect 19024 15308 19026 15328
rect 18970 15272 19026 15308
rect 19062 13640 19118 13696
rect 18878 12688 18934 12744
rect 18602 11872 18658 11928
rect 18510 11736 18566 11792
rect 18602 10512 18658 10568
rect 17590 6568 17646 6624
rect 17590 5480 17646 5536
rect 17498 1264 17554 1320
rect 18234 7540 18290 7576
rect 18234 7520 18236 7540
rect 18236 7520 18288 7540
rect 18288 7520 18290 7540
rect 18418 7248 18474 7304
rect 18602 7656 18658 7712
rect 18970 12164 19026 12200
rect 18970 12144 18972 12164
rect 18972 12144 19024 12164
rect 19024 12144 19026 12164
rect 19246 13504 19302 13560
rect 19430 15580 19432 15600
rect 19432 15580 19484 15600
rect 19484 15580 19486 15600
rect 19430 15544 19486 15580
rect 19430 14456 19486 14512
rect 19154 12860 19156 12880
rect 19156 12860 19208 12880
rect 19208 12860 19210 12880
rect 19154 12824 19210 12860
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 20074 16224 20130 16280
rect 20074 15680 20130 15736
rect 19982 15000 20038 15056
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19982 14320 20038 14376
rect 19706 13776 19762 13832
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 20258 23160 20314 23216
rect 20534 23840 20590 23896
rect 20350 20340 20352 20360
rect 20352 20340 20404 20360
rect 20404 20340 20406 20360
rect 20350 20304 20406 20340
rect 20534 19216 20590 19272
rect 20534 17040 20590 17096
rect 20166 14048 20222 14104
rect 20350 14048 20406 14104
rect 20166 13776 20222 13832
rect 20074 13504 20130 13560
rect 19338 12824 19394 12880
rect 19798 12824 19854 12880
rect 19338 12416 19394 12472
rect 19154 12180 19156 12200
rect 19156 12180 19208 12200
rect 19208 12180 19210 12200
rect 19154 12144 19210 12180
rect 18878 11620 18934 11656
rect 18878 11600 18880 11620
rect 18880 11600 18932 11620
rect 18932 11600 18934 11620
rect 18970 11192 19026 11248
rect 18786 9424 18842 9480
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 20258 12316 20260 12336
rect 20260 12316 20312 12336
rect 20312 12316 20314 12336
rect 20258 12280 20314 12316
rect 20258 11872 20314 11928
rect 19338 11500 19340 11520
rect 19340 11500 19392 11520
rect 19392 11500 19394 11520
rect 19338 11464 19394 11500
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19338 10684 19340 10704
rect 19340 10684 19392 10704
rect 19392 10684 19394 10704
rect 19338 10648 19394 10684
rect 19062 10140 19064 10160
rect 19064 10140 19116 10160
rect 19116 10140 19118 10160
rect 19062 10104 19118 10140
rect 18786 8472 18842 8528
rect 18602 7384 18658 7440
rect 19246 8372 19248 8392
rect 19248 8372 19300 8392
rect 19300 8372 19302 8392
rect 19246 8336 19302 8372
rect 19246 8064 19302 8120
rect 20258 11192 20314 11248
rect 20074 11056 20130 11112
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19338 7656 19394 7712
rect 18510 6452 18566 6488
rect 18510 6432 18512 6452
rect 18512 6432 18564 6452
rect 18564 6432 18566 6452
rect 19246 7112 19302 7168
rect 18050 5752 18106 5808
rect 18602 5752 18658 5808
rect 17774 5480 17830 5536
rect 17682 3848 17738 3904
rect 18418 5616 18474 5672
rect 18602 5652 18604 5672
rect 18604 5652 18656 5672
rect 18656 5652 18658 5672
rect 18602 5616 18658 5652
rect 18326 5480 18382 5536
rect 18234 3884 18236 3904
rect 18236 3884 18288 3904
rect 18288 3884 18290 3904
rect 18234 3848 18290 3884
rect 18510 5480 18566 5536
rect 18602 5092 18658 5128
rect 18602 5072 18604 5092
rect 18604 5072 18656 5092
rect 18656 5072 18658 5092
rect 18142 3440 18198 3496
rect 18418 3440 18474 3496
rect 18602 3304 18658 3360
rect 17866 1264 17922 1320
rect 18694 3168 18750 3224
rect 18694 2760 18750 2816
rect 18878 2352 18934 2408
rect 18418 1808 18474 1864
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19798 6704 19854 6760
rect 19982 6704 20038 6760
rect 19706 6160 19762 6216
rect 19982 6296 20038 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19338 5208 19394 5264
rect 19430 4800 19486 4856
rect 19430 3732 19486 3768
rect 19430 3712 19432 3732
rect 19432 3712 19484 3732
rect 19484 3712 19486 3732
rect 19338 3576 19394 3632
rect 19154 2216 19210 2272
rect 18970 1808 19026 1864
rect 20258 9968 20314 10024
rect 20258 9424 20314 9480
rect 20166 8472 20222 8528
rect 20350 7656 20406 7712
rect 20350 6976 20406 7032
rect 20534 12588 20536 12608
rect 20536 12588 20588 12608
rect 20588 12588 20590 12608
rect 20534 12552 20590 12588
rect 20902 24248 20958 24304
rect 20810 23840 20866 23896
rect 20718 23160 20774 23216
rect 20810 23024 20866 23080
rect 21086 23296 21142 23352
rect 22466 25336 22522 25392
rect 20810 22072 20866 22128
rect 20718 21800 20774 21856
rect 20718 20576 20774 20632
rect 20994 20984 21050 21040
rect 20902 20304 20958 20360
rect 20994 20032 21050 20088
rect 21086 19488 21142 19544
rect 20994 19080 21050 19136
rect 20718 15408 20774 15464
rect 20718 14476 20774 14512
rect 20718 14456 20720 14476
rect 20720 14456 20772 14476
rect 20772 14456 20774 14476
rect 20718 14184 20774 14240
rect 20626 8336 20682 8392
rect 20258 6604 20260 6624
rect 20260 6604 20312 6624
rect 20312 6604 20314 6624
rect 20258 6568 20314 6604
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20166 4004 20222 4040
rect 20166 3984 20168 4004
rect 20168 3984 20220 4004
rect 20220 3984 20222 4004
rect 20166 3576 20222 3632
rect 20258 3440 20314 3496
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19338 1400 19394 1456
rect 20166 1400 20222 1456
rect 21086 17992 21142 18048
rect 21546 23704 21602 23760
rect 21362 23568 21418 23624
rect 21454 23160 21510 23216
rect 21270 22752 21326 22808
rect 21454 22228 21510 22264
rect 21454 22208 21456 22228
rect 21456 22208 21508 22228
rect 21508 22208 21510 22228
rect 21270 22072 21326 22128
rect 21270 21936 21326 21992
rect 21638 21664 21694 21720
rect 21362 20204 21364 20224
rect 21364 20204 21416 20224
rect 21416 20204 21418 20224
rect 21362 20168 21418 20204
rect 21454 18844 21456 18864
rect 21456 18844 21508 18864
rect 21508 18844 21510 18864
rect 21454 18808 21510 18844
rect 21362 18536 21418 18592
rect 21454 18420 21510 18456
rect 21454 18400 21456 18420
rect 21456 18400 21508 18420
rect 21508 18400 21510 18420
rect 21546 17992 21602 18048
rect 20994 16496 21050 16552
rect 21086 15000 21142 15056
rect 20994 14728 21050 14784
rect 21178 13776 21234 13832
rect 21454 17076 21456 17096
rect 21456 17076 21508 17096
rect 21508 17076 21510 17096
rect 21454 17040 21510 17076
rect 21362 15000 21418 15056
rect 21362 13948 21364 13968
rect 21364 13948 21416 13968
rect 21416 13948 21418 13968
rect 21362 13912 21418 13948
rect 21638 15020 21694 15056
rect 21638 15000 21640 15020
rect 21640 15000 21692 15020
rect 21692 15000 21694 15020
rect 21822 20848 21878 20904
rect 21822 20440 21878 20496
rect 21638 12552 21694 12608
rect 21270 11872 21326 11928
rect 20994 9832 21050 9888
rect 20718 7520 20774 7576
rect 20350 3304 20406 3360
rect 20534 3984 20590 4040
rect 20626 3848 20682 3904
rect 20442 3032 20498 3088
rect 20074 992 20130 1048
rect 20626 856 20682 912
rect 20810 6860 20866 6896
rect 20810 6840 20812 6860
rect 20812 6840 20864 6860
rect 20864 6840 20866 6860
rect 20994 9016 21050 9072
rect 21454 10376 21510 10432
rect 21362 9696 21418 9752
rect 21546 9832 21602 9888
rect 22190 24520 22246 24576
rect 22098 22616 22154 22672
rect 22098 21292 22100 21312
rect 22100 21292 22152 21312
rect 22152 21292 22154 21312
rect 22098 21256 22154 21292
rect 22098 20168 22154 20224
rect 22374 21428 22376 21448
rect 22376 21428 22428 21448
rect 22428 21428 22430 21448
rect 22374 21392 22430 21428
rect 24766 27104 24822 27160
rect 24214 26016 24270 26072
rect 23386 25064 23442 25120
rect 22650 23976 22706 24032
rect 22834 23860 22890 23896
rect 22834 23840 22836 23860
rect 22836 23840 22888 23860
rect 22888 23840 22890 23860
rect 22834 23432 22890 23488
rect 22834 23160 22890 23216
rect 24766 25492 24822 25528
rect 24766 25472 24768 25492
rect 24768 25472 24820 25492
rect 24820 25472 24822 25492
rect 25042 25336 25098 25392
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24674 24928 24730 24984
rect 23110 23704 23166 23760
rect 22926 22072 22982 22128
rect 22558 21392 22614 21448
rect 22742 21256 22798 21312
rect 22650 20440 22706 20496
rect 22098 17040 22154 17096
rect 22190 16632 22246 16688
rect 22282 13524 22338 13560
rect 22282 13504 22284 13524
rect 22284 13504 22336 13524
rect 22336 13504 22338 13524
rect 22098 10240 22154 10296
rect 21270 8200 21326 8256
rect 20994 7248 21050 7304
rect 20994 6840 21050 6896
rect 20994 4548 21050 4584
rect 20994 4528 20996 4548
rect 20996 4528 21048 4548
rect 21048 4528 21050 4548
rect 20902 3848 20958 3904
rect 20810 3732 20866 3768
rect 21454 7248 21510 7304
rect 21730 8200 21786 8256
rect 21546 6976 21602 7032
rect 21822 7656 21878 7712
rect 21822 7520 21878 7576
rect 21270 6332 21272 6352
rect 21272 6332 21324 6352
rect 21324 6332 21326 6352
rect 21270 6296 21326 6332
rect 20810 3712 20812 3732
rect 20812 3712 20864 3732
rect 20864 3712 20866 3732
rect 21178 3460 21234 3496
rect 21178 3440 21180 3460
rect 21180 3440 21232 3460
rect 21232 3440 21234 3460
rect 21546 6568 21602 6624
rect 21546 6432 21602 6488
rect 22558 17484 22560 17504
rect 22560 17484 22612 17504
rect 22612 17484 22614 17504
rect 22558 17448 22614 17484
rect 22558 15544 22614 15600
rect 22650 14864 22706 14920
rect 22558 13504 22614 13560
rect 22466 12688 22522 12744
rect 22834 14184 22890 14240
rect 25410 26560 25466 26616
rect 24766 24384 24822 24440
rect 23754 23432 23810 23488
rect 23386 22772 23442 22808
rect 23386 22752 23388 22772
rect 23388 22752 23440 22772
rect 23440 22752 23442 22772
rect 23294 21664 23350 21720
rect 23018 19252 23020 19272
rect 23020 19252 23072 19272
rect 23072 19252 23074 19272
rect 23018 19216 23074 19252
rect 23018 15272 23074 15328
rect 23018 14068 23074 14104
rect 23018 14048 23020 14068
rect 23020 14048 23072 14068
rect 23072 14048 23074 14068
rect 22742 13368 22798 13424
rect 22466 12552 22522 12608
rect 22558 11736 22614 11792
rect 22374 10240 22430 10296
rect 22466 9968 22522 10024
rect 22006 9172 22062 9208
rect 22006 9152 22008 9172
rect 22008 9152 22060 9172
rect 22060 9152 22062 9172
rect 22006 8780 22008 8800
rect 22008 8780 22060 8800
rect 22060 8780 22062 8800
rect 22006 8744 22062 8780
rect 22098 8336 22154 8392
rect 22282 9424 22338 9480
rect 22282 7792 22338 7848
rect 22190 7384 22246 7440
rect 21454 4256 21510 4312
rect 21362 3712 21418 3768
rect 21914 5072 21970 5128
rect 22282 5092 22338 5128
rect 22282 5072 22284 5092
rect 22284 5072 22336 5092
rect 22336 5072 22338 5092
rect 22466 9696 22522 9752
rect 22558 8608 22614 8664
rect 22558 8064 22614 8120
rect 22834 11328 22890 11384
rect 23662 20712 23718 20768
rect 23570 20576 23626 20632
rect 23202 16632 23258 16688
rect 23478 20032 23534 20088
rect 23478 19796 23480 19816
rect 23480 19796 23532 19816
rect 23532 19796 23534 19816
rect 23478 19760 23534 19796
rect 23478 18264 23534 18320
rect 23754 20032 23810 20088
rect 23662 18572 23664 18592
rect 23664 18572 23716 18592
rect 23716 18572 23718 18592
rect 23662 18536 23718 18572
rect 23662 18128 23718 18184
rect 23662 17992 23718 18048
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24858 23568 24914 23624
rect 24950 23468 24952 23488
rect 24952 23468 25004 23488
rect 25004 23468 25006 23488
rect 24950 23432 25006 23468
rect 24766 23160 24822 23216
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24122 20168 24178 20224
rect 24030 19488 24086 19544
rect 24030 19080 24086 19136
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 25870 25744 25926 25800
rect 25686 23860 25742 23896
rect 25686 23840 25688 23860
rect 25688 23840 25740 23860
rect 25740 23840 25742 23860
rect 24766 21684 24822 21720
rect 24766 21664 24768 21684
rect 24768 21664 24820 21684
rect 24820 21664 24822 21684
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24674 19896 24730 19952
rect 24858 21140 24914 21176
rect 24858 21120 24860 21140
rect 24860 21120 24912 21140
rect 24912 21120 24914 21140
rect 25594 22616 25650 22672
rect 25226 22072 25282 22128
rect 25410 21936 25466 21992
rect 25226 21428 25228 21448
rect 25228 21428 25280 21448
rect 25280 21428 25282 21448
rect 25226 21392 25282 21428
rect 25134 20576 25190 20632
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24214 19352 24270 19408
rect 24582 19352 24638 19408
rect 24490 19080 24546 19136
rect 24674 19236 24730 19272
rect 24674 19216 24676 19236
rect 24676 19216 24728 19236
rect 24728 19216 24730 19236
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24122 18264 24178 18320
rect 23754 17584 23810 17640
rect 23570 17040 23626 17096
rect 23662 16496 23718 16552
rect 23478 16244 23534 16280
rect 23478 16224 23480 16244
rect 23480 16224 23532 16244
rect 23532 16224 23534 16244
rect 23478 14592 23534 14648
rect 23294 13368 23350 13424
rect 23478 12824 23534 12880
rect 22742 10240 22798 10296
rect 22742 7656 22798 7712
rect 22834 5888 22890 5944
rect 22834 5344 22890 5400
rect 21822 4120 21878 4176
rect 21730 2624 21786 2680
rect 21362 2372 21418 2408
rect 21362 2352 21364 2372
rect 21364 2352 21416 2372
rect 21416 2352 21418 2372
rect 22374 4120 22430 4176
rect 22282 3984 22338 4040
rect 22650 3848 22706 3904
rect 22282 3304 22338 3360
rect 22558 3168 22614 3224
rect 22742 3576 22798 3632
rect 23018 11228 23020 11248
rect 23020 11228 23072 11248
rect 23072 11228 23074 11248
rect 23018 11192 23074 11228
rect 23202 9868 23204 9888
rect 23204 9868 23256 9888
rect 23256 9868 23258 9888
rect 23202 9832 23258 9868
rect 23018 8064 23074 8120
rect 23018 4700 23020 4720
rect 23020 4700 23072 4720
rect 23072 4700 23074 4720
rect 23018 4664 23074 4700
rect 22834 3032 22890 3088
rect 24122 17856 24178 17912
rect 24030 17584 24086 17640
rect 23938 17312 23994 17368
rect 24398 17740 24454 17776
rect 24398 17720 24400 17740
rect 24400 17720 24452 17740
rect 24452 17720 24454 17740
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24674 17212 24676 17232
rect 24676 17212 24728 17232
rect 24728 17212 24730 17232
rect 24674 17176 24730 17212
rect 24030 16088 24086 16144
rect 24030 15816 24086 15872
rect 23938 15136 23994 15192
rect 24214 17040 24270 17096
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24214 15952 24270 16008
rect 24030 14728 24086 14784
rect 23938 13504 23994 13560
rect 24122 13504 24178 13560
rect 24030 13368 24086 13424
rect 24122 13132 24124 13152
rect 24124 13132 24176 13152
rect 24176 13132 24178 13152
rect 24122 13096 24178 13132
rect 24030 12688 24086 12744
rect 23478 11464 23534 11520
rect 23570 10784 23626 10840
rect 23478 10104 23534 10160
rect 23662 10104 23718 10160
rect 23846 12008 23902 12064
rect 23202 7656 23258 7712
rect 23202 7384 23258 7440
rect 23570 7792 23626 7848
rect 23478 7656 23534 7712
rect 23478 7540 23534 7576
rect 23478 7520 23480 7540
rect 23480 7520 23532 7540
rect 23532 7520 23534 7540
rect 23294 7248 23350 7304
rect 23202 6568 23258 6624
rect 23478 7112 23534 7168
rect 22742 2896 22798 2952
rect 22466 2760 22522 2816
rect 22374 1672 22430 1728
rect 22926 1128 22982 1184
rect 23202 992 23258 1048
rect 23478 4392 23534 4448
rect 23938 10376 23994 10432
rect 23754 4020 23756 4040
rect 23756 4020 23808 4040
rect 23808 4020 23810 4040
rect 23386 3032 23442 3088
rect 23294 856 23350 912
rect 23018 720 23074 776
rect 20902 40 20958 96
rect 22926 448 22982 504
rect 23754 3984 23810 4020
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 25042 18844 25044 18864
rect 25044 18844 25096 18864
rect 25096 18844 25098 18864
rect 25042 18808 25098 18844
rect 25226 20340 25228 20360
rect 25228 20340 25280 20360
rect 25280 20340 25282 20360
rect 25226 20304 25282 20340
rect 25226 19780 25282 19816
rect 25226 19760 25228 19780
rect 25228 19760 25280 19780
rect 25280 19760 25282 19780
rect 25226 18944 25282 19000
rect 25502 20984 25558 21040
rect 25502 19896 25558 19952
rect 24858 15680 24914 15736
rect 24858 14864 24914 14920
rect 24858 13912 24914 13968
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24306 12180 24308 12200
rect 24308 12180 24360 12200
rect 24360 12180 24362 12200
rect 24306 12144 24362 12180
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24214 11328 24270 11384
rect 24950 13268 24952 13288
rect 24952 13268 25004 13288
rect 25004 13268 25006 13288
rect 24950 13232 25006 13268
rect 25042 12416 25098 12472
rect 24858 11872 24914 11928
rect 24122 10804 24178 10840
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24122 10784 24124 10804
rect 24124 10784 24176 10804
rect 24176 10784 24178 10804
rect 24122 10376 24178 10432
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24674 9696 24730 9752
rect 24674 9288 24730 9344
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 25042 11736 25098 11792
rect 24950 10376 25006 10432
rect 24858 10104 24914 10160
rect 24858 9968 24914 10024
rect 24950 9868 24952 9888
rect 24952 9868 25004 9888
rect 25004 9868 25006 9888
rect 24950 9832 25006 9868
rect 25226 13640 25282 13696
rect 25226 12824 25282 12880
rect 25686 21528 25742 21584
rect 25594 17856 25650 17912
rect 25410 15952 25466 16008
rect 25410 13912 25466 13968
rect 25778 20884 25780 20904
rect 25780 20884 25832 20904
rect 25832 20884 25834 20904
rect 25778 20848 25834 20884
rect 26514 26152 26570 26208
rect 25962 24656 26018 24712
rect 25962 21292 25964 21312
rect 25964 21292 26016 21312
rect 26016 21292 26018 21312
rect 25962 21256 26018 21292
rect 25962 19760 26018 19816
rect 25870 17040 25926 17096
rect 25686 16496 25742 16552
rect 25594 11636 25596 11656
rect 25596 11636 25648 11656
rect 25648 11636 25650 11656
rect 25594 11600 25650 11636
rect 25226 10548 25228 10568
rect 25228 10548 25280 10568
rect 25280 10548 25282 10568
rect 25226 10512 25282 10548
rect 25134 9152 25190 9208
rect 25042 8508 25044 8528
rect 25044 8508 25096 8528
rect 25096 8508 25098 8528
rect 25042 8472 25098 8508
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24582 6976 24638 7032
rect 23938 3984 23994 4040
rect 23938 3848 23994 3904
rect 23662 2488 23718 2544
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24122 4256 24178 4312
rect 24122 3984 24178 4040
rect 24582 3848 24638 3904
rect 24582 3576 24638 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24122 2896 24178 2952
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24122 2100 24178 2136
rect 24122 2080 24124 2100
rect 24124 2080 24176 2100
rect 24176 2080 24178 2100
rect 24950 7248 25006 7304
rect 24858 3168 24914 3224
rect 25134 6976 25190 7032
rect 25134 5652 25136 5672
rect 25136 5652 25188 5672
rect 25188 5652 25190 5672
rect 25410 10260 25466 10296
rect 25410 10240 25412 10260
rect 25412 10240 25464 10260
rect 25464 10240 25466 10260
rect 25594 10920 25650 10976
rect 25502 9696 25558 9752
rect 25962 13504 26018 13560
rect 25962 11192 26018 11248
rect 25962 9580 26018 9616
rect 25962 9560 25964 9580
rect 25964 9560 26016 9580
rect 26016 9560 26018 9580
rect 25686 9052 25688 9072
rect 25688 9052 25740 9072
rect 25740 9052 25742 9072
rect 25686 9016 25742 9052
rect 25410 7964 25412 7984
rect 25412 7964 25464 7984
rect 25464 7964 25466 7984
rect 25410 7928 25466 7964
rect 25410 6860 25466 6896
rect 25410 6840 25412 6860
rect 25412 6840 25464 6860
rect 25464 6840 25466 6860
rect 25134 5616 25190 5652
rect 25226 5108 25228 5128
rect 25228 5108 25280 5128
rect 25280 5108 25282 5128
rect 25226 5072 25282 5108
rect 25042 3476 25044 3496
rect 25044 3476 25096 3496
rect 25096 3476 25098 3496
rect 25042 3440 25098 3476
rect 25134 3032 25190 3088
rect 25134 2896 25190 2952
rect 24950 1400 25006 1456
rect 24674 1264 24730 1320
rect 25502 4800 25558 4856
rect 25686 8200 25742 8256
rect 25778 6740 25780 6760
rect 25780 6740 25832 6760
rect 25832 6740 25834 6760
rect 25778 6704 25834 6740
rect 25962 6316 26018 6352
rect 25962 6296 25964 6316
rect 25964 6296 26016 6316
rect 26016 6296 26018 6316
rect 25410 2388 25412 2408
rect 25412 2388 25464 2408
rect 25464 2388 25466 2408
rect 25410 2352 25466 2388
rect 25502 1944 25558 2000
rect 25318 1128 25374 1184
rect 25594 1536 25650 1592
rect 25870 6024 25926 6080
rect 25778 5344 25834 5400
rect 25962 1944 26018 2000
rect 25686 1400 25742 1456
rect 27066 25608 27122 25664
rect 26330 22208 26386 22264
rect 26330 20032 26386 20088
rect 26238 18300 26240 18320
rect 26240 18300 26292 18320
rect 26292 18300 26294 18320
rect 26238 18264 26294 18300
rect 26330 16768 26386 16824
rect 26146 15000 26202 15056
rect 26422 10376 26478 10432
rect 26330 8880 26386 8936
rect 26330 5752 26386 5808
rect 26238 5208 26294 5264
rect 26238 4936 26294 4992
rect 26330 4528 26386 4584
rect 26238 3848 26294 3904
rect 26330 3188 26386 3224
rect 26330 3168 26332 3188
rect 26332 3168 26384 3188
rect 26384 3168 26386 3188
rect 26606 3032 26662 3088
rect 26514 2488 26570 2544
rect 26422 1808 26478 1864
rect 26422 312 26478 368
rect 27066 584 27122 640
rect 26698 312 26754 368
rect 27342 176 27398 232
<< metal3 >>
rect 0 27706 480 27736
rect 3366 27706 3372 27708
rect 0 27646 3372 27706
rect 0 27616 480 27646
rect 3366 27644 3372 27646
rect 3436 27644 3442 27708
rect 21173 27706 21239 27709
rect 27520 27706 28000 27736
rect 21173 27704 28000 27706
rect 21173 27648 21178 27704
rect 21234 27648 28000 27704
rect 21173 27646 28000 27648
rect 21173 27643 21239 27646
rect 27520 27616 28000 27646
rect 24761 27162 24827 27165
rect 27520 27162 28000 27192
rect 24761 27160 28000 27162
rect 24761 27104 24766 27160
rect 24822 27104 28000 27160
rect 24761 27102 28000 27104
rect 24761 27099 24827 27102
rect 27520 27072 28000 27102
rect 0 27026 480 27056
rect 1117 27026 1183 27029
rect 0 27024 1183 27026
rect 0 26968 1122 27024
rect 1178 26968 1183 27024
rect 0 26966 1183 26968
rect 0 26936 480 26966
rect 1117 26963 1183 26966
rect 25405 26618 25471 26621
rect 27520 26618 28000 26648
rect 25405 26616 28000 26618
rect 25405 26560 25410 26616
rect 25466 26560 28000 26616
rect 25405 26558 28000 26560
rect 25405 26555 25471 26558
rect 27520 26528 28000 26558
rect 10133 26482 10199 26485
rect 17309 26482 17375 26485
rect 10133 26480 17375 26482
rect 10133 26424 10138 26480
rect 10194 26424 17314 26480
rect 17370 26424 17375 26480
rect 10133 26422 17375 26424
rect 10133 26419 10199 26422
rect 17309 26419 17375 26422
rect 0 26346 480 26376
rect 1393 26346 1459 26349
rect 0 26344 1459 26346
rect 0 26288 1398 26344
rect 1454 26288 1459 26344
rect 0 26286 1459 26288
rect 0 26256 480 26286
rect 1393 26283 1459 26286
rect 9949 26346 10015 26349
rect 16113 26346 16179 26349
rect 9949 26344 16179 26346
rect 9949 26288 9954 26344
rect 10010 26288 16118 26344
rect 16174 26288 16179 26344
rect 9949 26286 16179 26288
rect 9949 26283 10015 26286
rect 16113 26283 16179 26286
rect 2129 26210 2195 26213
rect 19333 26210 19399 26213
rect 2129 26208 19399 26210
rect 2129 26152 2134 26208
rect 2190 26152 19338 26208
rect 19394 26152 19399 26208
rect 2129 26150 19399 26152
rect 2129 26147 2195 26150
rect 19333 26147 19399 26150
rect 26366 26148 26372 26212
rect 26436 26210 26442 26212
rect 26509 26210 26575 26213
rect 26436 26208 26575 26210
rect 26436 26152 26514 26208
rect 26570 26152 26575 26208
rect 26436 26150 26575 26152
rect 26436 26148 26442 26150
rect 26509 26147 26575 26150
rect 2681 26074 2747 26077
rect 13353 26074 13419 26077
rect 2681 26072 13419 26074
rect 2681 26016 2686 26072
rect 2742 26016 13358 26072
rect 13414 26016 13419 26072
rect 2681 26014 13419 26016
rect 2681 26011 2747 26014
rect 13353 26011 13419 26014
rect 24209 26074 24275 26077
rect 27520 26074 28000 26104
rect 24209 26072 28000 26074
rect 24209 26016 24214 26072
rect 24270 26016 28000 26072
rect 24209 26014 28000 26016
rect 24209 26011 24275 26014
rect 27520 25984 28000 26014
rect 289 25938 355 25941
rect 15745 25938 15811 25941
rect 289 25936 15811 25938
rect 289 25880 294 25936
rect 350 25880 15750 25936
rect 15806 25880 15811 25936
rect 289 25878 15811 25880
rect 289 25875 355 25878
rect 15745 25875 15811 25878
rect 16021 25938 16087 25941
rect 20662 25938 20668 25940
rect 16021 25936 20668 25938
rect 16021 25880 16026 25936
rect 16082 25880 20668 25936
rect 16021 25878 20668 25880
rect 16021 25875 16087 25878
rect 20662 25876 20668 25878
rect 20732 25876 20738 25940
rect 1209 25802 1275 25805
rect 11145 25802 11211 25805
rect 25865 25802 25931 25805
rect 1209 25800 10794 25802
rect 1209 25744 1214 25800
rect 1270 25744 10794 25800
rect 1209 25742 10794 25744
rect 1209 25739 1275 25742
rect 0 25666 480 25696
rect 1577 25666 1643 25669
rect 0 25664 1643 25666
rect 0 25608 1582 25664
rect 1638 25608 1643 25664
rect 0 25606 1643 25608
rect 10734 25666 10794 25742
rect 11145 25800 25931 25802
rect 11145 25744 11150 25800
rect 11206 25744 25870 25800
rect 25926 25744 25931 25800
rect 11145 25742 25931 25744
rect 11145 25739 11211 25742
rect 25865 25739 25931 25742
rect 10734 25606 19258 25666
rect 0 25576 480 25606
rect 1577 25603 1643 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 5390 25468 5396 25532
rect 5460 25530 5466 25532
rect 10133 25530 10199 25533
rect 18965 25530 19031 25533
rect 5460 25528 10199 25530
rect 5460 25472 10138 25528
rect 10194 25472 10199 25528
rect 5460 25470 10199 25472
rect 5460 25468 5466 25470
rect 10133 25467 10199 25470
rect 10734 25528 19031 25530
rect 10734 25472 18970 25528
rect 19026 25472 19031 25528
rect 10734 25470 19031 25472
rect 9397 25394 9463 25397
rect 10734 25394 10794 25470
rect 18965 25467 19031 25470
rect 9397 25392 10794 25394
rect 9397 25336 9402 25392
rect 9458 25336 10794 25392
rect 9397 25334 10794 25336
rect 13721 25394 13787 25397
rect 15561 25394 15627 25397
rect 13721 25392 15627 25394
rect 13721 25336 13726 25392
rect 13782 25336 15566 25392
rect 15622 25336 15627 25392
rect 13721 25334 15627 25336
rect 19198 25394 19258 25606
rect 26918 25604 26924 25668
rect 26988 25666 26994 25668
rect 27061 25666 27127 25669
rect 26988 25664 27127 25666
rect 26988 25608 27066 25664
rect 27122 25608 27127 25664
rect 26988 25606 27127 25608
rect 26988 25604 26994 25606
rect 27061 25603 27127 25606
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24761 25530 24827 25533
rect 27520 25530 28000 25560
rect 24761 25528 28000 25530
rect 24761 25472 24766 25528
rect 24822 25472 28000 25528
rect 24761 25470 28000 25472
rect 24761 25467 24827 25470
rect 27520 25440 28000 25470
rect 22461 25394 22527 25397
rect 25037 25394 25103 25397
rect 19198 25392 25103 25394
rect 19198 25336 22466 25392
rect 22522 25336 25042 25392
rect 25098 25336 25103 25392
rect 19198 25334 25103 25336
rect 9397 25331 9463 25334
rect 13721 25331 13787 25334
rect 15561 25331 15627 25334
rect 22461 25331 22527 25334
rect 25037 25331 25103 25334
rect 5809 25258 5875 25261
rect 6310 25258 6316 25260
rect 5809 25256 6316 25258
rect 5809 25200 5814 25256
rect 5870 25200 6316 25256
rect 5809 25198 6316 25200
rect 5809 25195 5875 25198
rect 6310 25196 6316 25198
rect 6380 25196 6386 25260
rect 7649 25258 7715 25261
rect 11145 25258 11211 25261
rect 17309 25258 17375 25261
rect 21030 25258 21036 25260
rect 7649 25256 11211 25258
rect 7649 25200 7654 25256
rect 7710 25200 11150 25256
rect 11206 25200 11211 25256
rect 7649 25198 11211 25200
rect 7649 25195 7715 25198
rect 11145 25195 11211 25198
rect 14414 25198 15394 25258
rect 7189 25122 7255 25125
rect 14414 25122 14474 25198
rect 7189 25120 14474 25122
rect 7189 25064 7194 25120
rect 7250 25064 14474 25120
rect 7189 25062 14474 25064
rect 15334 25122 15394 25198
rect 17309 25256 21036 25258
rect 17309 25200 17314 25256
rect 17370 25200 21036 25256
rect 17309 25198 21036 25200
rect 17309 25195 17375 25198
rect 21030 25196 21036 25198
rect 21100 25196 21106 25260
rect 23381 25122 23447 25125
rect 15334 25120 23447 25122
rect 15334 25064 23386 25120
rect 23442 25064 23447 25120
rect 15334 25062 23447 25064
rect 7189 25059 7255 25062
rect 23381 25059 23447 25062
rect 5610 25056 5930 25057
rect 0 24986 480 25016
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 1485 24986 1551 24989
rect 0 24984 1551 24986
rect 0 24928 1490 24984
rect 1546 24928 1551 24984
rect 0 24926 1551 24928
rect 0 24896 480 24926
rect 1485 24923 1551 24926
rect 1761 24986 1827 24989
rect 2681 24986 2747 24989
rect 1761 24984 2747 24986
rect 1761 24928 1766 24984
rect 1822 24928 2686 24984
rect 2742 24928 2747 24984
rect 1761 24926 2747 24928
rect 1761 24923 1827 24926
rect 2681 24923 2747 24926
rect 9581 24986 9647 24989
rect 14365 24986 14431 24989
rect 9581 24984 14431 24986
rect 9581 24928 9586 24984
rect 9642 24928 14370 24984
rect 14426 24928 14431 24984
rect 9581 24926 14431 24928
rect 9581 24923 9647 24926
rect 14365 24923 14431 24926
rect 16021 24986 16087 24989
rect 20161 24986 20227 24989
rect 16021 24984 20227 24986
rect 16021 24928 16026 24984
rect 16082 24928 20166 24984
rect 20222 24928 20227 24984
rect 16021 24926 20227 24928
rect 16021 24923 16087 24926
rect 20161 24923 20227 24926
rect 24669 24986 24735 24989
rect 27520 24986 28000 25016
rect 24669 24984 28000 24986
rect 24669 24928 24674 24984
rect 24730 24928 28000 24984
rect 24669 24926 28000 24928
rect 24669 24923 24735 24926
rect 27520 24896 28000 24926
rect 3049 24852 3115 24853
rect 2998 24850 3004 24852
rect 2958 24790 3004 24850
rect 3068 24848 3115 24852
rect 3110 24792 3115 24848
rect 2998 24788 3004 24790
rect 3068 24788 3115 24792
rect 3182 24788 3188 24852
rect 3252 24850 3258 24852
rect 3601 24850 3667 24853
rect 3252 24848 3667 24850
rect 3252 24792 3606 24848
rect 3662 24792 3667 24848
rect 3252 24790 3667 24792
rect 3252 24788 3258 24790
rect 3049 24787 3115 24788
rect 3601 24787 3667 24790
rect 9765 24852 9831 24853
rect 9765 24848 9812 24852
rect 9876 24850 9882 24852
rect 13077 24850 13143 24853
rect 14825 24850 14891 24853
rect 16757 24850 16823 24853
rect 9765 24792 9770 24848
rect 9765 24788 9812 24792
rect 9876 24790 9922 24850
rect 13077 24848 16823 24850
rect 13077 24792 13082 24848
rect 13138 24792 14830 24848
rect 14886 24792 16762 24848
rect 16818 24792 16823 24848
rect 13077 24790 16823 24792
rect 9876 24788 9882 24790
rect 9765 24787 9831 24788
rect 13077 24787 13143 24790
rect 14825 24787 14891 24790
rect 16757 24787 16823 24790
rect 7005 24714 7071 24717
rect 12249 24714 12315 24717
rect 13997 24714 14063 24717
rect 7005 24712 10794 24714
rect 7005 24656 7010 24712
rect 7066 24656 10794 24712
rect 7005 24654 10794 24656
rect 7005 24651 7071 24654
rect 8702 24516 8708 24580
rect 8772 24578 8778 24580
rect 9489 24578 9555 24581
rect 8772 24576 9555 24578
rect 8772 24520 9494 24576
rect 9550 24520 9555 24576
rect 8772 24518 9555 24520
rect 10734 24578 10794 24654
rect 12249 24712 14063 24714
rect 12249 24656 12254 24712
rect 12310 24656 14002 24712
rect 14058 24656 14063 24712
rect 12249 24654 14063 24656
rect 12249 24651 12315 24654
rect 13997 24651 14063 24654
rect 19057 24714 19123 24717
rect 25957 24714 26023 24717
rect 19057 24712 26023 24714
rect 19057 24656 19062 24712
rect 19118 24656 25962 24712
rect 26018 24656 26023 24712
rect 19057 24654 26023 24656
rect 19057 24651 19123 24654
rect 25957 24651 26023 24654
rect 16481 24578 16547 24581
rect 10734 24576 16547 24578
rect 10734 24520 16486 24576
rect 16542 24520 16547 24576
rect 10734 24518 16547 24520
rect 8772 24516 8778 24518
rect 9489 24515 9555 24518
rect 16481 24515 16547 24518
rect 20294 24516 20300 24580
rect 20364 24578 20370 24580
rect 22185 24578 22251 24581
rect 20364 24576 22251 24578
rect 20364 24520 22190 24576
rect 22246 24520 22251 24576
rect 20364 24518 22251 24520
rect 20364 24516 20370 24518
rect 22185 24515 22251 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 2497 24442 2563 24445
rect 9305 24442 9371 24445
rect 2497 24440 9371 24442
rect 2497 24384 2502 24440
rect 2558 24384 9310 24440
rect 9366 24384 9371 24440
rect 2497 24382 9371 24384
rect 2497 24379 2563 24382
rect 9305 24379 9371 24382
rect 16021 24442 16087 24445
rect 19241 24442 19307 24445
rect 16021 24440 19307 24442
rect 16021 24384 16026 24440
rect 16082 24384 19246 24440
rect 19302 24384 19307 24440
rect 16021 24382 19307 24384
rect 16021 24379 16087 24382
rect 19241 24379 19307 24382
rect 24761 24442 24827 24445
rect 27520 24442 28000 24472
rect 24761 24440 28000 24442
rect 24761 24384 24766 24440
rect 24822 24384 28000 24440
rect 24761 24382 28000 24384
rect 24761 24379 24827 24382
rect 27520 24352 28000 24382
rect 0 24306 480 24336
rect 1577 24306 1643 24309
rect 0 24304 1643 24306
rect 0 24248 1582 24304
rect 1638 24248 1643 24304
rect 0 24246 1643 24248
rect 0 24216 480 24246
rect 1577 24243 1643 24246
rect 8017 24306 8083 24309
rect 9438 24306 9444 24308
rect 8017 24304 9444 24306
rect 8017 24248 8022 24304
rect 8078 24248 9444 24304
rect 8017 24246 9444 24248
rect 8017 24243 8083 24246
rect 9438 24244 9444 24246
rect 9508 24244 9514 24308
rect 9581 24306 9647 24309
rect 13905 24306 13971 24309
rect 14549 24306 14615 24309
rect 9581 24304 14615 24306
rect 9581 24248 9586 24304
rect 9642 24248 13910 24304
rect 13966 24248 14554 24304
rect 14610 24248 14615 24304
rect 9581 24246 14615 24248
rect 9581 24243 9647 24246
rect 13905 24243 13971 24246
rect 14549 24243 14615 24246
rect 18321 24306 18387 24309
rect 20897 24306 20963 24309
rect 18321 24304 20963 24306
rect 18321 24248 18326 24304
rect 18382 24248 20902 24304
rect 20958 24248 20963 24304
rect 18321 24246 20963 24248
rect 18321 24243 18387 24246
rect 20897 24243 20963 24246
rect 3693 24170 3759 24173
rect 7465 24170 7531 24173
rect 8753 24170 8819 24173
rect 11053 24170 11119 24173
rect 3693 24168 7531 24170
rect 3693 24112 3698 24168
rect 3754 24112 7470 24168
rect 7526 24112 7531 24168
rect 3693 24110 7531 24112
rect 3693 24107 3759 24110
rect 7465 24107 7531 24110
rect 7606 24168 11119 24170
rect 7606 24112 8758 24168
rect 8814 24112 11058 24168
rect 11114 24112 11119 24168
rect 7606 24110 11119 24112
rect 7005 24034 7071 24037
rect 7606 24034 7666 24110
rect 8753 24107 8819 24110
rect 11053 24107 11119 24110
rect 11789 24170 11855 24173
rect 12525 24170 12591 24173
rect 11789 24168 12591 24170
rect 11789 24112 11794 24168
rect 11850 24112 12530 24168
rect 12586 24112 12591 24168
rect 11789 24110 12591 24112
rect 11789 24107 11855 24110
rect 12525 24107 12591 24110
rect 14365 24170 14431 24173
rect 18137 24170 18203 24173
rect 22318 24170 22324 24172
rect 14365 24168 15394 24170
rect 14365 24112 14370 24168
rect 14426 24112 15394 24168
rect 14365 24110 15394 24112
rect 14365 24107 14431 24110
rect 7005 24032 7666 24034
rect 7005 23976 7010 24032
rect 7066 23976 7666 24032
rect 7005 23974 7666 23976
rect 7005 23971 7071 23974
rect 8150 23972 8156 24036
rect 8220 24034 8226 24036
rect 11881 24034 11947 24037
rect 8220 24032 11947 24034
rect 8220 23976 11886 24032
rect 11942 23976 11947 24032
rect 8220 23974 11947 23976
rect 15334 24034 15394 24110
rect 18137 24168 22324 24170
rect 18137 24112 18142 24168
rect 18198 24112 22324 24168
rect 18137 24110 22324 24112
rect 18137 24107 18203 24110
rect 22318 24108 22324 24110
rect 22388 24108 22394 24172
rect 22645 24034 22711 24037
rect 15334 24032 22711 24034
rect 15334 23976 22650 24032
rect 22706 23976 22711 24032
rect 15334 23974 22711 23976
rect 8220 23972 8226 23974
rect 11881 23971 11947 23974
rect 22645 23971 22711 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 7557 23898 7623 23901
rect 10777 23898 10843 23901
rect 7557 23896 10843 23898
rect 7557 23840 7562 23896
rect 7618 23840 10782 23896
rect 10838 23840 10843 23896
rect 7557 23838 10843 23840
rect 7557 23835 7623 23838
rect 10777 23835 10843 23838
rect 15745 23898 15811 23901
rect 16665 23898 16731 23901
rect 20529 23898 20595 23901
rect 20805 23900 20871 23901
rect 20805 23898 20852 23900
rect 15745 23896 20595 23898
rect 15745 23840 15750 23896
rect 15806 23840 16670 23896
rect 16726 23840 20534 23896
rect 20590 23840 20595 23896
rect 15745 23838 20595 23840
rect 20760 23896 20852 23898
rect 20760 23840 20810 23896
rect 20760 23838 20852 23840
rect 15745 23835 15811 23838
rect 16665 23835 16731 23838
rect 20529 23835 20595 23838
rect 20805 23836 20852 23838
rect 20916 23836 20922 23900
rect 21950 23836 21956 23900
rect 22020 23898 22026 23900
rect 22829 23898 22895 23901
rect 22020 23896 22895 23898
rect 22020 23840 22834 23896
rect 22890 23840 22895 23896
rect 22020 23838 22895 23840
rect 22020 23836 22026 23838
rect 20805 23835 20871 23836
rect 22829 23835 22895 23838
rect 25681 23898 25747 23901
rect 27520 23898 28000 23928
rect 25681 23896 28000 23898
rect 25681 23840 25686 23896
rect 25742 23840 28000 23896
rect 25681 23838 28000 23840
rect 25681 23835 25747 23838
rect 27520 23808 28000 23838
rect 6729 23762 6795 23765
rect 14273 23762 14339 23765
rect 6729 23760 14339 23762
rect 6729 23704 6734 23760
rect 6790 23704 14278 23760
rect 14334 23704 14339 23760
rect 6729 23702 14339 23704
rect 6729 23699 6795 23702
rect 14273 23699 14339 23702
rect 15653 23762 15719 23765
rect 21541 23762 21607 23765
rect 23105 23762 23171 23765
rect 15653 23760 20776 23762
rect 15653 23704 15658 23760
rect 15714 23704 20776 23760
rect 15653 23702 20776 23704
rect 15653 23699 15719 23702
rect 0 23626 480 23656
rect 2589 23626 2655 23629
rect 0 23624 2655 23626
rect 0 23568 2594 23624
rect 2650 23568 2655 23624
rect 0 23566 2655 23568
rect 0 23536 480 23566
rect 2589 23563 2655 23566
rect 6545 23626 6611 23629
rect 11789 23626 11855 23629
rect 6545 23624 11855 23626
rect 6545 23568 6550 23624
rect 6606 23568 11794 23624
rect 11850 23568 11855 23624
rect 6545 23566 11855 23568
rect 6545 23563 6611 23566
rect 11789 23563 11855 23566
rect 11973 23626 12039 23629
rect 13445 23626 13511 23629
rect 17953 23626 18019 23629
rect 11973 23624 13511 23626
rect 11973 23568 11978 23624
rect 12034 23568 13450 23624
rect 13506 23568 13511 23624
rect 11973 23566 13511 23568
rect 11973 23563 12039 23566
rect 13445 23563 13511 23566
rect 13678 23624 18019 23626
rect 13678 23568 17958 23624
rect 18014 23568 18019 23624
rect 13678 23566 18019 23568
rect 4153 23490 4219 23493
rect 5022 23490 5028 23492
rect 4153 23488 5028 23490
rect 4153 23432 4158 23488
rect 4214 23432 5028 23488
rect 4153 23430 5028 23432
rect 4153 23427 4219 23430
rect 5022 23428 5028 23430
rect 5092 23428 5098 23492
rect 5441 23490 5507 23493
rect 9990 23490 9996 23492
rect 5441 23488 9996 23490
rect 5441 23432 5446 23488
rect 5502 23432 9996 23488
rect 5441 23430 9996 23432
rect 5441 23427 5507 23430
rect 9990 23428 9996 23430
rect 10060 23428 10066 23492
rect 12801 23490 12867 23493
rect 13678 23490 13738 23566
rect 17953 23563 18019 23566
rect 18597 23626 18663 23629
rect 20478 23626 20484 23628
rect 18597 23624 20484 23626
rect 18597 23568 18602 23624
rect 18658 23568 20484 23624
rect 18597 23566 20484 23568
rect 18597 23563 18663 23566
rect 20478 23564 20484 23566
rect 20548 23564 20554 23628
rect 12801 23488 13738 23490
rect 12801 23432 12806 23488
rect 12862 23432 13738 23488
rect 12801 23430 13738 23432
rect 16205 23490 16271 23493
rect 18597 23492 18663 23493
rect 20069 23492 20135 23493
rect 16614 23490 16620 23492
rect 16205 23488 16620 23490
rect 16205 23432 16210 23488
rect 16266 23432 16620 23488
rect 16205 23430 16620 23432
rect 12801 23427 12867 23430
rect 16205 23427 16271 23430
rect 16614 23428 16620 23430
rect 16684 23428 16690 23492
rect 18597 23490 18644 23492
rect 18552 23488 18644 23490
rect 18552 23432 18602 23488
rect 18552 23430 18644 23432
rect 18597 23428 18644 23430
rect 18708 23428 18714 23492
rect 20069 23488 20116 23492
rect 20180 23490 20186 23492
rect 20069 23432 20074 23488
rect 20069 23428 20116 23432
rect 20180 23430 20226 23490
rect 20180 23428 20186 23430
rect 18597 23427 18663 23428
rect 20069 23427 20135 23428
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 5625 23354 5691 23357
rect 6126 23354 6132 23356
rect 5625 23352 6132 23354
rect 5625 23296 5630 23352
rect 5686 23296 6132 23352
rect 5625 23294 6132 23296
rect 5625 23291 5691 23294
rect 6126 23292 6132 23294
rect 6196 23292 6202 23356
rect 8109 23354 8175 23357
rect 9857 23354 9923 23357
rect 8109 23352 9923 23354
rect 8109 23296 8114 23352
rect 8170 23296 9862 23352
rect 9918 23296 9923 23352
rect 8109 23294 9923 23296
rect 8109 23291 8175 23294
rect 9857 23291 9923 23294
rect 15377 23354 15443 23357
rect 19149 23354 19215 23357
rect 15377 23352 19215 23354
rect 15377 23296 15382 23352
rect 15438 23296 19154 23352
rect 19210 23296 19215 23352
rect 15377 23294 19215 23296
rect 15377 23291 15443 23294
rect 19149 23291 19215 23294
rect 2405 23218 2471 23221
rect 6821 23218 6887 23221
rect 8569 23218 8635 23221
rect 2405 23216 6700 23218
rect 2405 23160 2410 23216
rect 2466 23160 6700 23216
rect 2405 23158 6700 23160
rect 2405 23155 2471 23158
rect 3601 23082 3667 23085
rect 6453 23082 6519 23085
rect 3601 23080 6519 23082
rect 3601 23024 3606 23080
rect 3662 23024 6458 23080
rect 6514 23024 6519 23080
rect 3601 23022 6519 23024
rect 3601 23019 3667 23022
rect 6453 23019 6519 23022
rect 0 22946 480 22976
rect 2681 22946 2747 22949
rect 0 22944 2747 22946
rect 0 22888 2686 22944
rect 2742 22888 2747 22944
rect 0 22886 2747 22888
rect 6640 22946 6700 23158
rect 6821 23216 8635 23218
rect 6821 23160 6826 23216
rect 6882 23160 8574 23216
rect 8630 23160 8635 23216
rect 6821 23158 8635 23160
rect 6821 23155 6887 23158
rect 8569 23155 8635 23158
rect 8845 23218 8911 23221
rect 9070 23218 9076 23220
rect 8845 23216 9076 23218
rect 8845 23160 8850 23216
rect 8906 23160 9076 23216
rect 8845 23158 9076 23160
rect 8845 23155 8911 23158
rect 9070 23156 9076 23158
rect 9140 23156 9146 23220
rect 17585 23218 17651 23221
rect 19382 23218 19626 23252
rect 20716 23221 20776 23702
rect 21541 23760 23171 23762
rect 21541 23704 21546 23760
rect 21602 23704 23110 23760
rect 23166 23704 23171 23760
rect 21541 23702 23171 23704
rect 21541 23699 21607 23702
rect 23105 23699 23171 23702
rect 21357 23626 21423 23629
rect 24853 23626 24919 23629
rect 21357 23624 24919 23626
rect 21357 23568 21362 23624
rect 21418 23568 24858 23624
rect 24914 23568 24919 23624
rect 21357 23566 24919 23568
rect 21357 23563 21423 23566
rect 24853 23563 24919 23566
rect 22829 23490 22895 23493
rect 23749 23492 23815 23493
rect 23054 23490 23060 23492
rect 22829 23488 23060 23490
rect 22829 23432 22834 23488
rect 22890 23432 23060 23488
rect 22829 23430 23060 23432
rect 22829 23427 22895 23430
rect 23054 23428 23060 23430
rect 23124 23428 23130 23492
rect 23749 23488 23796 23492
rect 23860 23490 23866 23492
rect 23749 23432 23754 23488
rect 23749 23428 23796 23432
rect 23860 23430 23906 23490
rect 23860 23428 23866 23430
rect 24710 23428 24716 23492
rect 24780 23490 24786 23492
rect 24945 23490 25011 23493
rect 24780 23488 25011 23490
rect 24780 23432 24950 23488
rect 25006 23432 25011 23488
rect 24780 23430 25011 23432
rect 24780 23428 24786 23430
rect 23749 23427 23815 23428
rect 24945 23427 25011 23430
rect 21081 23354 21147 23357
rect 21582 23354 21588 23356
rect 21081 23352 21588 23354
rect 21081 23296 21086 23352
rect 21142 23296 21588 23352
rect 21081 23294 21588 23296
rect 21081 23291 21147 23294
rect 21582 23292 21588 23294
rect 21652 23292 21658 23356
rect 20253 23218 20319 23221
rect 17585 23216 20319 23218
rect 17585 23160 17590 23216
rect 17646 23192 20258 23216
rect 17646 23160 19442 23192
rect 17585 23158 19442 23160
rect 19566 23160 20258 23192
rect 20314 23160 20319 23216
rect 19566 23158 20319 23160
rect 17585 23155 17651 23158
rect 20253 23155 20319 23158
rect 20713 23216 20779 23221
rect 20713 23160 20718 23216
rect 20774 23160 20779 23216
rect 20713 23155 20779 23160
rect 21449 23218 21515 23221
rect 22829 23218 22895 23221
rect 21449 23216 22895 23218
rect 21449 23160 21454 23216
rect 21510 23160 22834 23216
rect 22890 23160 22895 23216
rect 21449 23158 22895 23160
rect 21449 23155 21515 23158
rect 22829 23155 22895 23158
rect 24761 23218 24827 23221
rect 27520 23218 28000 23248
rect 24761 23216 28000 23218
rect 24761 23160 24766 23216
rect 24822 23160 28000 23216
rect 24761 23158 28000 23160
rect 24761 23155 24827 23158
rect 27520 23128 28000 23158
rect 8017 23082 8083 23085
rect 11646 23082 11652 23084
rect 8017 23080 11652 23082
rect 8017 23024 8022 23080
rect 8078 23024 11652 23080
rect 8017 23022 11652 23024
rect 8017 23019 8083 23022
rect 11646 23020 11652 23022
rect 11716 23020 11722 23084
rect 15101 23082 15167 23085
rect 16849 23082 16915 23085
rect 15101 23080 16915 23082
rect 15101 23024 15106 23080
rect 15162 23024 16854 23080
rect 16910 23024 16915 23080
rect 15101 23022 16915 23024
rect 15101 23019 15167 23022
rect 16849 23019 16915 23022
rect 17677 23082 17743 23085
rect 19333 23082 19399 23085
rect 17677 23080 19399 23082
rect 17677 23024 17682 23080
rect 17738 23024 19338 23080
rect 19394 23024 19399 23080
rect 17677 23022 19399 23024
rect 17677 23019 17743 23022
rect 19333 23019 19399 23022
rect 20805 23082 20871 23085
rect 23974 23082 23980 23084
rect 20805 23080 23980 23082
rect 20805 23024 20810 23080
rect 20866 23024 23980 23080
rect 20805 23022 23980 23024
rect 20805 23019 20871 23022
rect 23974 23020 23980 23022
rect 24044 23020 24050 23084
rect 8109 22946 8175 22949
rect 6640 22944 8175 22946
rect 6640 22888 8114 22944
rect 8170 22888 8175 22944
rect 6640 22886 8175 22888
rect 0 22856 480 22886
rect 2681 22883 2747 22886
rect 8109 22883 8175 22886
rect 16757 22946 16823 22949
rect 19333 22946 19399 22949
rect 16757 22944 19399 22946
rect 16757 22888 16762 22944
rect 16818 22888 19338 22944
rect 19394 22888 19399 22944
rect 16757 22886 19399 22888
rect 16757 22883 16823 22886
rect 19333 22883 19399 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 8477 22810 8543 22813
rect 9438 22810 9444 22812
rect 8477 22808 9444 22810
rect 8477 22752 8482 22808
rect 8538 22752 9444 22808
rect 8477 22750 9444 22752
rect 8477 22747 8543 22750
rect 9438 22748 9444 22750
rect 9508 22748 9514 22812
rect 9576 22748 9582 22812
rect 9646 22810 9652 22812
rect 13813 22810 13879 22813
rect 21265 22810 21331 22813
rect 23381 22810 23447 22813
rect 9646 22808 13879 22810
rect 9646 22752 13818 22808
rect 13874 22752 13879 22808
rect 9646 22750 13879 22752
rect 9646 22748 9652 22750
rect 13813 22747 13879 22750
rect 17542 22808 23447 22810
rect 17542 22752 21270 22808
rect 21326 22752 23386 22808
rect 23442 22752 23447 22808
rect 17542 22750 23447 22752
rect 8201 22674 8267 22677
rect 8334 22674 8340 22676
rect 8201 22672 8340 22674
rect 8201 22616 8206 22672
rect 8262 22616 8340 22672
rect 8201 22614 8340 22616
rect 8201 22611 8267 22614
rect 8334 22612 8340 22614
rect 8404 22612 8410 22676
rect 17542 22674 17602 22750
rect 21265 22747 21331 22750
rect 23381 22747 23447 22750
rect 9078 22614 17602 22674
rect 18229 22674 18295 22677
rect 19333 22674 19399 22677
rect 18229 22672 19399 22674
rect 18229 22616 18234 22672
rect 18290 22616 19338 22672
rect 19394 22616 19399 22672
rect 18229 22614 19399 22616
rect 3049 22538 3115 22541
rect 3918 22538 3924 22540
rect 3049 22536 3924 22538
rect 3049 22480 3054 22536
rect 3110 22480 3924 22536
rect 3049 22478 3924 22480
rect 3049 22475 3115 22478
rect 3918 22476 3924 22478
rect 3988 22476 3994 22540
rect 5717 22402 5783 22405
rect 6545 22404 6611 22405
rect 6126 22402 6132 22404
rect 5717 22400 6132 22402
rect 5717 22344 5722 22400
rect 5778 22344 6132 22400
rect 5717 22342 6132 22344
rect 5717 22339 5783 22342
rect 6126 22340 6132 22342
rect 6196 22340 6202 22404
rect 6494 22340 6500 22404
rect 6564 22402 6611 22404
rect 7097 22402 7163 22405
rect 8661 22404 8727 22405
rect 7966 22402 7972 22404
rect 6564 22400 6656 22402
rect 6606 22344 6656 22400
rect 6564 22342 6656 22344
rect 7097 22400 7972 22402
rect 7097 22344 7102 22400
rect 7158 22344 7972 22400
rect 7097 22342 7972 22344
rect 6564 22340 6611 22342
rect 6545 22339 6611 22340
rect 7097 22339 7163 22342
rect 7966 22340 7972 22342
rect 8036 22340 8042 22404
rect 8661 22402 8708 22404
rect 8616 22400 8708 22402
rect 8616 22344 8666 22400
rect 8616 22342 8708 22344
rect 8661 22340 8708 22342
rect 8772 22340 8778 22404
rect 8661 22339 8727 22340
rect 0 22266 480 22296
rect 2405 22266 2471 22269
rect 0 22264 2471 22266
rect 0 22208 2410 22264
rect 2466 22208 2471 22264
rect 0 22206 2471 22208
rect 0 22176 480 22206
rect 2405 22203 2471 22206
rect 4838 22204 4844 22268
rect 4908 22266 4914 22268
rect 6361 22266 6427 22269
rect 9078 22266 9138 22614
rect 18229 22611 18295 22614
rect 19333 22611 19399 22614
rect 19701 22674 19767 22677
rect 22093 22674 22159 22677
rect 19701 22672 22159 22674
rect 19701 22616 19706 22672
rect 19762 22616 22098 22672
rect 22154 22616 22159 22672
rect 19701 22614 22159 22616
rect 19701 22611 19767 22614
rect 22093 22611 22159 22614
rect 25589 22674 25655 22677
rect 27520 22674 28000 22704
rect 25589 22672 28000 22674
rect 25589 22616 25594 22672
rect 25650 22616 28000 22672
rect 25589 22614 28000 22616
rect 25589 22611 25655 22614
rect 27520 22584 28000 22614
rect 9305 22538 9371 22541
rect 12157 22538 12223 22541
rect 9305 22536 12223 22538
rect 9305 22480 9310 22536
rect 9366 22480 12162 22536
rect 12218 22480 12223 22536
rect 9305 22478 12223 22480
rect 9305 22475 9371 22478
rect 12157 22475 12223 22478
rect 12525 22538 12591 22541
rect 19333 22538 19399 22541
rect 12525 22536 19399 22538
rect 12525 22480 12530 22536
rect 12586 22480 19338 22536
rect 19394 22480 19399 22536
rect 12525 22478 19399 22480
rect 12525 22475 12591 22478
rect 19333 22475 19399 22478
rect 20662 22340 20668 22404
rect 20732 22402 20738 22404
rect 21766 22402 21772 22404
rect 20732 22342 21772 22402
rect 20732 22340 20738 22342
rect 21766 22340 21772 22342
rect 21836 22340 21842 22404
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 4908 22264 6427 22266
rect 4908 22208 6366 22264
rect 6422 22208 6427 22264
rect 4908 22206 6427 22208
rect 4908 22204 4914 22206
rect 6361 22203 6427 22206
rect 6502 22206 9138 22266
rect 9213 22266 9279 22269
rect 11237 22266 11303 22269
rect 11697 22266 11763 22269
rect 9213 22264 9322 22266
rect 9213 22208 9218 22264
rect 9274 22208 9322 22264
rect 6502 22133 6562 22206
rect 9213 22203 9322 22208
rect 11237 22264 11763 22266
rect 11237 22208 11242 22264
rect 11298 22208 11702 22264
rect 11758 22208 11763 22264
rect 11237 22206 11763 22208
rect 11237 22203 11303 22206
rect 11697 22203 11763 22206
rect 13077 22266 13143 22269
rect 18505 22266 18571 22269
rect 13077 22264 18571 22266
rect 13077 22208 13082 22264
rect 13138 22208 18510 22264
rect 18566 22208 18571 22264
rect 13077 22206 18571 22208
rect 13077 22203 13143 22206
rect 18505 22203 18571 22206
rect 19149 22266 19215 22269
rect 21449 22266 21515 22269
rect 26325 22266 26391 22269
rect 19149 22264 19442 22266
rect 19149 22208 19154 22264
rect 19210 22208 19442 22264
rect 19149 22206 19442 22208
rect 19149 22203 19215 22206
rect 6453 22128 6562 22133
rect 6453 22072 6458 22128
rect 6514 22072 6562 22128
rect 6453 22070 6562 22072
rect 7833 22130 7899 22133
rect 8150 22130 8156 22132
rect 7833 22128 8156 22130
rect 7833 22072 7838 22128
rect 7894 22072 8156 22128
rect 7833 22070 8156 22072
rect 6453 22067 6519 22070
rect 7833 22067 7899 22070
rect 8150 22068 8156 22070
rect 8220 22068 8226 22132
rect 8702 22068 8708 22132
rect 8772 22130 8778 22132
rect 9262 22130 9322 22203
rect 8772 22070 9322 22130
rect 10961 22130 11027 22133
rect 12341 22130 12407 22133
rect 10961 22128 12407 22130
rect 10961 22072 10966 22128
rect 11022 22072 12346 22128
rect 12402 22072 12407 22128
rect 10961 22070 12407 22072
rect 8772 22068 8778 22070
rect 10961 22067 11027 22070
rect 12341 22067 12407 22070
rect 15285 22130 15351 22133
rect 15653 22130 15719 22133
rect 15285 22128 15719 22130
rect 15285 22072 15290 22128
rect 15346 22072 15658 22128
rect 15714 22072 15719 22128
rect 15285 22070 15719 22072
rect 19382 22130 19442 22206
rect 21449 22264 26391 22266
rect 21449 22208 21454 22264
rect 21510 22208 26330 22264
rect 26386 22208 26391 22264
rect 21449 22206 26391 22208
rect 21449 22203 21515 22206
rect 26325 22203 26391 22206
rect 19609 22130 19675 22133
rect 19382 22128 19675 22130
rect 19382 22072 19614 22128
rect 19670 22072 19675 22128
rect 19382 22070 19675 22072
rect 15285 22067 15351 22070
rect 15653 22067 15719 22070
rect 19609 22067 19675 22070
rect 20805 22132 20871 22133
rect 20805 22128 20852 22132
rect 20916 22130 20922 22132
rect 21265 22130 21331 22133
rect 22686 22130 22692 22132
rect 20805 22072 20810 22128
rect 20805 22068 20852 22072
rect 20916 22070 20962 22130
rect 21265 22128 22692 22130
rect 21265 22072 21270 22128
rect 21326 22072 22692 22128
rect 21265 22070 22692 22072
rect 20916 22068 20922 22070
rect 20805 22067 20871 22068
rect 21265 22067 21331 22070
rect 22686 22068 22692 22070
rect 22756 22068 22762 22132
rect 22921 22130 22987 22133
rect 25221 22130 25287 22133
rect 27520 22130 28000 22160
rect 22878 22128 22987 22130
rect 22878 22072 22926 22128
rect 22982 22072 22987 22128
rect 22878 22067 22987 22072
rect 23246 22128 25287 22130
rect 23246 22072 25226 22128
rect 25282 22072 25287 22128
rect 23246 22070 25287 22072
rect 4981 21994 5047 21997
rect 6637 21994 6703 21997
rect 6913 21994 6979 21997
rect 4981 21992 6979 21994
rect 4981 21936 4986 21992
rect 5042 21936 6642 21992
rect 6698 21936 6918 21992
rect 6974 21936 6979 21992
rect 4981 21934 6979 21936
rect 4981 21931 5047 21934
rect 6637 21931 6703 21934
rect 6913 21931 6979 21934
rect 8017 21994 8083 21997
rect 9857 21994 9923 21997
rect 8017 21992 9923 21994
rect 8017 21936 8022 21992
rect 8078 21936 9862 21992
rect 9918 21936 9923 21992
rect 8017 21934 9923 21936
rect 8017 21931 8083 21934
rect 9857 21931 9923 21934
rect 9990 21932 9996 21996
rect 10060 21994 10066 21996
rect 11145 21994 11211 21997
rect 10060 21992 11211 21994
rect 10060 21936 11150 21992
rect 11206 21936 11211 21992
rect 10060 21934 11211 21936
rect 10060 21932 10066 21934
rect 11145 21931 11211 21934
rect 15101 21994 15167 21997
rect 17033 21994 17099 21997
rect 15101 21992 17099 21994
rect 15101 21936 15106 21992
rect 15162 21936 17038 21992
rect 17094 21936 17099 21992
rect 15101 21934 17099 21936
rect 15101 21931 15167 21934
rect 17033 21931 17099 21934
rect 18086 21932 18092 21996
rect 18156 21994 18162 21996
rect 21265 21994 21331 21997
rect 22878 21994 22938 22067
rect 18156 21934 20914 21994
rect 18156 21932 18162 21934
rect 4705 21858 4771 21861
rect 5390 21858 5396 21860
rect 4705 21856 5396 21858
rect 4705 21800 4710 21856
rect 4766 21800 5396 21856
rect 4705 21798 5396 21800
rect 4705 21795 4771 21798
rect 5390 21796 5396 21798
rect 5460 21796 5466 21860
rect 9489 21858 9555 21861
rect 10041 21858 10107 21861
rect 11053 21858 11119 21861
rect 9489 21856 11119 21858
rect 9489 21800 9494 21856
rect 9550 21800 10046 21856
rect 10102 21800 11058 21856
rect 11114 21800 11119 21856
rect 9489 21798 11119 21800
rect 9489 21795 9555 21798
rect 10041 21795 10107 21798
rect 11053 21795 11119 21798
rect 16389 21858 16455 21861
rect 20713 21858 20779 21861
rect 16389 21856 20779 21858
rect 16389 21800 16394 21856
rect 16450 21800 20718 21856
rect 20774 21800 20779 21856
rect 16389 21798 20779 21800
rect 20854 21858 20914 21934
rect 21265 21992 22938 21994
rect 21265 21936 21270 21992
rect 21326 21936 22938 21992
rect 21265 21934 22938 21936
rect 21265 21931 21331 21934
rect 23246 21858 23306 22070
rect 25221 22067 25287 22070
rect 25408 22070 28000 22130
rect 25408 21997 25468 22070
rect 27520 22040 28000 22070
rect 25405 21992 25471 21997
rect 25405 21936 25410 21992
rect 25466 21936 25471 21992
rect 25405 21931 25471 21936
rect 20854 21798 23306 21858
rect 16389 21795 16455 21798
rect 20713 21795 20779 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 8293 21722 8359 21725
rect 3926 21662 4768 21722
rect 0 21586 480 21616
rect 1669 21586 1735 21589
rect 0 21584 1735 21586
rect 0 21528 1674 21584
rect 1730 21528 1735 21584
rect 0 21526 1735 21528
rect 0 21496 480 21526
rect 1669 21523 1735 21526
rect 2589 21178 2655 21181
rect 3926 21180 3986 21662
rect 4521 21588 4587 21589
rect 4470 21524 4476 21588
rect 4540 21586 4587 21588
rect 4708 21586 4768 21662
rect 8158 21720 8359 21722
rect 8158 21664 8298 21720
rect 8354 21664 8359 21720
rect 8158 21662 8359 21664
rect 8158 21586 8218 21662
rect 8293 21659 8359 21662
rect 8702 21660 8708 21724
rect 8772 21722 8778 21724
rect 8845 21722 8911 21725
rect 11053 21722 11119 21725
rect 8772 21720 8911 21722
rect 8772 21664 8850 21720
rect 8906 21664 8911 21720
rect 8772 21662 8911 21664
rect 8772 21660 8778 21662
rect 8845 21659 8911 21662
rect 9630 21720 11119 21722
rect 9630 21664 11058 21720
rect 11114 21664 11119 21720
rect 9630 21662 11119 21664
rect 9630 21620 9690 21662
rect 11053 21659 11119 21662
rect 15377 21722 15443 21725
rect 20662 21722 20668 21724
rect 15377 21720 20668 21722
rect 15377 21664 15382 21720
rect 15438 21664 20668 21720
rect 15377 21662 20668 21664
rect 15377 21659 15443 21662
rect 20662 21660 20668 21662
rect 20732 21660 20738 21724
rect 21030 21660 21036 21724
rect 21100 21722 21106 21724
rect 21633 21722 21699 21725
rect 21100 21720 21699 21722
rect 21100 21664 21638 21720
rect 21694 21664 21699 21720
rect 21100 21662 21699 21664
rect 21100 21660 21106 21662
rect 21633 21659 21699 21662
rect 22870 21660 22876 21724
rect 22940 21722 22946 21724
rect 23289 21722 23355 21725
rect 22940 21720 23355 21722
rect 22940 21664 23294 21720
rect 23350 21664 23355 21720
rect 22940 21662 23355 21664
rect 22940 21660 22946 21662
rect 23289 21659 23355 21662
rect 24761 21722 24827 21725
rect 25262 21722 25268 21724
rect 24761 21720 25268 21722
rect 24761 21664 24766 21720
rect 24822 21664 25268 21720
rect 24761 21662 25268 21664
rect 24761 21659 24827 21662
rect 25262 21660 25268 21662
rect 25332 21660 25338 21724
rect 9446 21589 9690 21620
rect 4540 21584 4632 21586
rect 4582 21528 4632 21584
rect 4540 21526 4632 21528
rect 4708 21526 8218 21586
rect 9397 21584 9690 21589
rect 9397 21528 9402 21584
rect 9458 21560 9690 21584
rect 9458 21528 9506 21560
rect 9397 21526 9506 21528
rect 9584 21526 9690 21560
rect 10685 21586 10751 21589
rect 13629 21586 13695 21589
rect 10685 21584 13695 21586
rect 10685 21528 10690 21584
rect 10746 21528 13634 21584
rect 13690 21528 13695 21584
rect 10685 21526 13695 21528
rect 4540 21524 4587 21526
rect 4521 21523 4587 21524
rect 9397 21523 9463 21526
rect 10685 21523 10751 21526
rect 13629 21523 13695 21526
rect 14641 21586 14707 21589
rect 21398 21586 21404 21588
rect 14641 21584 21404 21586
rect 14641 21528 14646 21584
rect 14702 21528 21404 21584
rect 14641 21526 21404 21528
rect 14641 21523 14707 21526
rect 21398 21524 21404 21526
rect 21468 21524 21474 21588
rect 25681 21586 25747 21589
rect 27520 21586 28000 21616
rect 25681 21584 28000 21586
rect 25681 21528 25686 21584
rect 25742 21528 28000 21584
rect 25681 21526 28000 21528
rect 25681 21523 25747 21526
rect 27520 21496 28000 21526
rect 4654 21388 4660 21452
rect 4724 21450 4730 21452
rect 5993 21450 6059 21453
rect 14549 21450 14615 21453
rect 4724 21448 6059 21450
rect 4724 21392 5998 21448
rect 6054 21392 6059 21448
rect 4724 21390 6059 21392
rect 4724 21388 4730 21390
rect 5993 21387 6059 21390
rect 10044 21448 14615 21450
rect 10044 21392 14554 21448
rect 14610 21392 14615 21448
rect 10044 21390 14615 21392
rect 4061 21314 4127 21317
rect 6678 21314 6684 21316
rect 4061 21312 6684 21314
rect 4061 21256 4066 21312
rect 4122 21256 6684 21312
rect 4061 21254 6684 21256
rect 4061 21251 4127 21254
rect 6678 21252 6684 21254
rect 6748 21252 6754 21316
rect 7005 21314 7071 21317
rect 7005 21312 9506 21314
rect 7005 21256 7010 21312
rect 7066 21256 9506 21312
rect 7005 21254 9506 21256
rect 7005 21251 7071 21254
rect 3918 21178 3924 21180
rect 2589 21176 3924 21178
rect 2589 21120 2594 21176
rect 2650 21120 3924 21176
rect 2589 21118 3924 21120
rect 2589 21115 2655 21118
rect 3918 21116 3924 21118
rect 3988 21116 3994 21180
rect 4153 21178 4219 21181
rect 7414 21178 7420 21180
rect 4153 21176 7420 21178
rect 4153 21120 4158 21176
rect 4214 21120 7420 21176
rect 4153 21118 7420 21120
rect 4153 21115 4219 21118
rect 7414 21116 7420 21118
rect 7484 21116 7490 21180
rect 9446 21178 9506 21254
rect 10044 21178 10104 21390
rect 14549 21387 14615 21390
rect 14825 21450 14891 21453
rect 16297 21450 16363 21453
rect 14825 21448 16363 21450
rect 14825 21392 14830 21448
rect 14886 21392 16302 21448
rect 16358 21392 16363 21448
rect 14825 21390 16363 21392
rect 14825 21387 14891 21390
rect 16297 21387 16363 21390
rect 21030 21388 21036 21452
rect 21100 21450 21106 21452
rect 22369 21450 22435 21453
rect 21100 21448 22435 21450
rect 21100 21392 22374 21448
rect 22430 21392 22435 21448
rect 21100 21390 22435 21392
rect 21100 21388 21106 21390
rect 22369 21387 22435 21390
rect 22553 21450 22619 21453
rect 25221 21450 25287 21453
rect 22553 21448 25287 21450
rect 22553 21392 22558 21448
rect 22614 21392 25226 21448
rect 25282 21392 25287 21448
rect 22553 21390 25287 21392
rect 22553 21387 22619 21390
rect 25221 21387 25287 21390
rect 16481 21314 16547 21317
rect 19425 21314 19491 21317
rect 16481 21312 19491 21314
rect 16481 21256 16486 21312
rect 16542 21256 19430 21312
rect 19486 21256 19491 21312
rect 16481 21254 19491 21256
rect 16481 21251 16547 21254
rect 19425 21251 19491 21254
rect 22093 21314 22159 21317
rect 22737 21314 22803 21317
rect 25957 21314 26023 21317
rect 22093 21312 26023 21314
rect 22093 21256 22098 21312
rect 22154 21256 22742 21312
rect 22798 21256 25962 21312
rect 26018 21256 26023 21312
rect 22093 21254 26023 21256
rect 22093 21251 22159 21254
rect 22737 21251 22803 21254
rect 25957 21251 26023 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 9446 21118 10104 21178
rect 15009 21178 15075 21181
rect 15377 21178 15443 21181
rect 16389 21178 16455 21181
rect 24853 21178 24919 21181
rect 15009 21176 16455 21178
rect 15009 21120 15014 21176
rect 15070 21120 15382 21176
rect 15438 21120 16394 21176
rect 16450 21120 16455 21176
rect 15009 21118 16455 21120
rect 15009 21115 15075 21118
rect 15377 21115 15443 21118
rect 16389 21115 16455 21118
rect 21176 21176 24919 21178
rect 21176 21120 24858 21176
rect 24914 21120 24919 21176
rect 21176 21118 24919 21120
rect 0 21042 480 21072
rect 7005 21042 7071 21045
rect 0 21040 7071 21042
rect 0 20984 7010 21040
rect 7066 20984 7071 21040
rect 0 20982 7071 20984
rect 0 20952 480 20982
rect 7005 20979 7071 20982
rect 7189 21042 7255 21045
rect 12709 21042 12775 21045
rect 7189 21040 12775 21042
rect 7189 20984 7194 21040
rect 7250 20984 12714 21040
rect 12770 20984 12775 21040
rect 7189 20982 12775 20984
rect 7189 20979 7255 20982
rect 12709 20979 12775 20982
rect 17033 21042 17099 21045
rect 20989 21042 21055 21045
rect 17033 21040 21055 21042
rect 17033 20984 17038 21040
rect 17094 20984 20994 21040
rect 21050 20984 21055 21040
rect 17033 20982 21055 20984
rect 17033 20979 17099 20982
rect 20989 20979 21055 20982
rect 3325 20906 3391 20909
rect 4429 20906 4495 20909
rect 3052 20904 3391 20906
rect 3052 20848 3330 20904
rect 3386 20848 3391 20904
rect 3052 20846 3391 20848
rect 3052 20637 3112 20846
rect 3325 20843 3391 20846
rect 3926 20904 4495 20906
rect 3926 20848 4434 20904
rect 4490 20848 4495 20904
rect 3926 20846 4495 20848
rect 3693 20772 3759 20773
rect 3693 20768 3740 20772
rect 3804 20770 3810 20772
rect 3693 20712 3698 20768
rect 3693 20708 3740 20712
rect 3804 20710 3850 20770
rect 3804 20708 3810 20710
rect 3693 20707 3759 20708
rect 2865 20634 2931 20637
rect 1718 20632 2931 20634
rect 1718 20576 2870 20632
rect 2926 20576 2931 20632
rect 1718 20574 2931 20576
rect 0 20362 480 20392
rect 1718 20365 1778 20574
rect 2865 20571 2931 20574
rect 3049 20632 3115 20637
rect 3049 20576 3054 20632
rect 3110 20576 3115 20632
rect 3049 20571 3115 20576
rect 3693 20634 3759 20637
rect 3926 20634 3986 20846
rect 4429 20843 4495 20846
rect 5625 20906 5691 20909
rect 7097 20906 7163 20909
rect 5625 20904 7163 20906
rect 5625 20848 5630 20904
rect 5686 20848 7102 20904
rect 7158 20848 7163 20904
rect 5625 20846 7163 20848
rect 5625 20843 5691 20846
rect 7097 20843 7163 20846
rect 8201 20906 8267 20909
rect 9673 20906 9739 20909
rect 8201 20904 9739 20906
rect 8201 20848 8206 20904
rect 8262 20848 9678 20904
rect 9734 20848 9739 20904
rect 8201 20846 9739 20848
rect 8201 20843 8267 20846
rect 9673 20843 9739 20846
rect 11697 20906 11763 20909
rect 15285 20906 15351 20909
rect 11697 20904 15351 20906
rect 11697 20848 11702 20904
rect 11758 20848 15290 20904
rect 15346 20848 15351 20904
rect 11697 20846 15351 20848
rect 11697 20843 11763 20846
rect 15285 20843 15351 20846
rect 19333 20906 19399 20909
rect 21176 20906 21236 21118
rect 24853 21115 24919 21118
rect 21398 20980 21404 21044
rect 21468 21042 21474 21044
rect 25497 21042 25563 21045
rect 27520 21042 28000 21072
rect 21468 21040 25563 21042
rect 21468 20984 25502 21040
rect 25558 20984 25563 21040
rect 21468 20982 25563 20984
rect 21468 20980 21474 20982
rect 25497 20979 25563 20982
rect 26006 20982 28000 21042
rect 19333 20904 21236 20906
rect 19333 20848 19338 20904
rect 19394 20848 21236 20904
rect 19333 20846 21236 20848
rect 21817 20906 21883 20909
rect 25773 20906 25839 20909
rect 21817 20904 25839 20906
rect 21817 20848 21822 20904
rect 21878 20848 25778 20904
rect 25834 20848 25839 20904
rect 21817 20846 25839 20848
rect 19333 20843 19399 20846
rect 21817 20843 21883 20846
rect 25773 20843 25839 20846
rect 9397 20770 9463 20773
rect 9765 20770 9831 20773
rect 12617 20770 12683 20773
rect 9397 20768 12683 20770
rect 9397 20712 9402 20768
rect 9458 20712 9770 20768
rect 9826 20712 12622 20768
rect 12678 20712 12683 20768
rect 9397 20710 12683 20712
rect 9397 20707 9463 20710
rect 9765 20707 9831 20710
rect 12617 20707 12683 20710
rect 15510 20708 15516 20772
rect 15580 20770 15586 20772
rect 18086 20770 18092 20772
rect 15580 20710 18092 20770
rect 15580 20708 15586 20710
rect 18086 20708 18092 20710
rect 18156 20708 18162 20772
rect 18505 20770 18571 20773
rect 23657 20770 23723 20773
rect 18505 20768 23723 20770
rect 18505 20712 18510 20768
rect 18566 20712 23662 20768
rect 23718 20712 23723 20768
rect 18505 20710 23723 20712
rect 18505 20707 18571 20710
rect 23657 20707 23723 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 3693 20632 3986 20634
rect 3693 20576 3698 20632
rect 3754 20576 3986 20632
rect 3693 20574 3986 20576
rect 9213 20634 9279 20637
rect 11237 20634 11303 20637
rect 9213 20632 11303 20634
rect 9213 20576 9218 20632
rect 9274 20576 11242 20632
rect 11298 20576 11303 20632
rect 9213 20574 11303 20576
rect 3693 20571 3759 20574
rect 9213 20571 9279 20574
rect 11237 20571 11303 20574
rect 11646 20572 11652 20636
rect 11716 20634 11722 20636
rect 14733 20634 14799 20637
rect 11716 20632 14799 20634
rect 11716 20576 14738 20632
rect 14794 20576 14799 20632
rect 11716 20574 14799 20576
rect 11716 20572 11722 20574
rect 14733 20571 14799 20574
rect 17861 20634 17927 20637
rect 18965 20634 19031 20637
rect 20713 20634 20779 20637
rect 23565 20634 23631 20637
rect 17861 20632 20779 20634
rect 17861 20576 17866 20632
rect 17922 20576 18970 20632
rect 19026 20576 20718 20632
rect 20774 20576 20779 20632
rect 17861 20574 20779 20576
rect 17861 20571 17927 20574
rect 18965 20571 19031 20574
rect 20713 20571 20779 20574
rect 21774 20632 23631 20634
rect 21774 20576 23570 20632
rect 23626 20576 23631 20632
rect 21774 20574 23631 20576
rect 21774 20501 21834 20574
rect 23565 20571 23631 20574
rect 25129 20634 25195 20637
rect 26006 20634 26066 20982
rect 27520 20952 28000 20982
rect 25129 20632 26066 20634
rect 25129 20576 25134 20632
rect 25190 20576 26066 20632
rect 25129 20574 26066 20576
rect 25129 20571 25195 20574
rect 1853 20498 1919 20501
rect 5625 20498 5691 20501
rect 8334 20498 8340 20500
rect 1853 20496 2928 20498
rect 1853 20440 1858 20496
rect 1914 20440 2928 20496
rect 1853 20438 2928 20440
rect 1853 20435 1919 20438
rect 1577 20362 1643 20365
rect 0 20360 1643 20362
rect 0 20304 1582 20360
rect 1638 20304 1643 20360
rect 0 20302 1643 20304
rect 1718 20360 1827 20365
rect 1718 20304 1766 20360
rect 1822 20304 1827 20360
rect 1718 20302 1827 20304
rect 0 20272 480 20302
rect 1577 20299 1643 20302
rect 1761 20299 1827 20302
rect 2405 20360 2471 20365
rect 2405 20304 2410 20360
rect 2466 20304 2471 20360
rect 2405 20299 2471 20304
rect 2868 20362 2928 20438
rect 5625 20496 8340 20498
rect 5625 20440 5630 20496
rect 5686 20440 8340 20496
rect 5625 20438 8340 20440
rect 5625 20435 5691 20438
rect 8334 20436 8340 20438
rect 8404 20436 8410 20500
rect 9489 20498 9555 20501
rect 14641 20498 14707 20501
rect 17309 20498 17375 20501
rect 9489 20496 14474 20498
rect 9489 20440 9494 20496
rect 9550 20440 14474 20496
rect 9489 20438 14474 20440
rect 9489 20435 9555 20438
rect 12617 20362 12683 20365
rect 2868 20360 12683 20362
rect 2868 20304 12622 20360
rect 12678 20304 12683 20360
rect 2868 20302 12683 20304
rect 12617 20299 12683 20302
rect 13169 20362 13235 20365
rect 13302 20362 13308 20364
rect 13169 20360 13308 20362
rect 13169 20304 13174 20360
rect 13230 20304 13308 20360
rect 13169 20302 13308 20304
rect 13169 20299 13235 20302
rect 13302 20300 13308 20302
rect 13372 20362 13378 20364
rect 13537 20362 13603 20365
rect 13372 20360 13603 20362
rect 13372 20304 13542 20360
rect 13598 20304 13603 20360
rect 13372 20302 13603 20304
rect 14414 20362 14474 20438
rect 14641 20496 17375 20498
rect 14641 20440 14646 20496
rect 14702 20440 17314 20496
rect 17370 20440 17375 20496
rect 14641 20438 17375 20440
rect 21774 20496 21883 20501
rect 21774 20440 21822 20496
rect 21878 20440 21883 20496
rect 21774 20438 21883 20440
rect 14641 20435 14707 20438
rect 17309 20435 17375 20438
rect 21817 20435 21883 20438
rect 22645 20498 22711 20501
rect 27520 20498 28000 20528
rect 22645 20496 28000 20498
rect 22645 20440 22650 20496
rect 22706 20440 28000 20496
rect 22645 20438 28000 20440
rect 22645 20435 22711 20438
rect 27520 20408 28000 20438
rect 15653 20362 15719 20365
rect 16389 20362 16455 20365
rect 20345 20362 20411 20365
rect 20897 20364 20963 20365
rect 20846 20362 20852 20364
rect 14414 20360 20411 20362
rect 14414 20304 15658 20360
rect 15714 20304 16394 20360
rect 16450 20304 20350 20360
rect 20406 20304 20411 20360
rect 14414 20302 20411 20304
rect 20806 20302 20852 20362
rect 20916 20360 20963 20364
rect 25221 20362 25287 20365
rect 20958 20304 20963 20360
rect 13372 20300 13378 20302
rect 13537 20299 13603 20302
rect 15653 20299 15719 20302
rect 16389 20299 16455 20302
rect 20345 20299 20411 20302
rect 20846 20300 20852 20302
rect 20916 20300 20963 20304
rect 20897 20299 20963 20300
rect 21084 20360 25287 20362
rect 21084 20304 25226 20360
rect 25282 20304 25287 20360
rect 21084 20302 25287 20304
rect 2408 20226 2468 20299
rect 9673 20228 9739 20229
rect 8150 20226 8156 20228
rect 2408 20166 8156 20226
rect 8150 20164 8156 20166
rect 8220 20164 8226 20228
rect 9622 20164 9628 20228
rect 9692 20226 9739 20228
rect 11329 20226 11395 20229
rect 11881 20226 11947 20229
rect 16205 20226 16271 20229
rect 21084 20226 21144 20302
rect 25221 20299 25287 20302
rect 9692 20224 9784 20226
rect 9734 20168 9784 20224
rect 9692 20166 9784 20168
rect 11329 20224 16271 20226
rect 11329 20168 11334 20224
rect 11390 20168 11886 20224
rect 11942 20168 16210 20224
rect 16266 20168 16271 20224
rect 11329 20166 16271 20168
rect 9692 20164 9739 20166
rect 9673 20163 9739 20164
rect 11329 20163 11395 20166
rect 11881 20163 11947 20166
rect 16205 20163 16271 20166
rect 20854 20166 21144 20226
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 2497 20090 2563 20093
rect 2630 20090 2636 20092
rect 2497 20088 2636 20090
rect 2497 20032 2502 20088
rect 2558 20032 2636 20088
rect 2497 20030 2636 20032
rect 2497 20027 2563 20030
rect 2630 20028 2636 20030
rect 2700 20028 2706 20092
rect 3182 20028 3188 20092
rect 3252 20090 3258 20092
rect 3969 20090 4035 20093
rect 7189 20090 7255 20093
rect 3252 20088 7255 20090
rect 3252 20032 3974 20088
rect 4030 20032 7194 20088
rect 7250 20032 7255 20088
rect 3252 20030 7255 20032
rect 3252 20028 3258 20030
rect 3969 20027 4035 20030
rect 7189 20027 7255 20030
rect 7373 20090 7439 20093
rect 9765 20090 9831 20093
rect 7373 20088 9831 20090
rect 7373 20032 7378 20088
rect 7434 20032 9770 20088
rect 9826 20032 9831 20088
rect 7373 20030 9831 20032
rect 7373 20027 7439 20030
rect 9765 20027 9831 20030
rect 9949 20092 10015 20093
rect 9949 20088 9996 20092
rect 10060 20090 10066 20092
rect 9949 20032 9954 20088
rect 9949 20028 9996 20032
rect 10060 20030 10106 20090
rect 10060 20028 10066 20030
rect 10910 20028 10916 20092
rect 10980 20090 10986 20092
rect 17166 20090 17172 20092
rect 10980 20030 17172 20090
rect 10980 20028 10986 20030
rect 17166 20028 17172 20030
rect 17236 20028 17242 20092
rect 9949 20027 10015 20028
rect 3233 19954 3299 19957
rect 14733 19954 14799 19957
rect 3233 19952 14799 19954
rect 3233 19896 3238 19952
rect 3294 19896 14738 19952
rect 14794 19896 14799 19952
rect 3233 19894 14799 19896
rect 3233 19891 3299 19894
rect 14733 19891 14799 19894
rect 15745 19954 15811 19957
rect 20854 19954 20914 20166
rect 21214 20164 21220 20228
rect 21284 20226 21290 20228
rect 21357 20226 21423 20229
rect 21284 20224 21423 20226
rect 21284 20168 21362 20224
rect 21418 20168 21423 20224
rect 21284 20166 21423 20168
rect 21284 20164 21290 20166
rect 21357 20163 21423 20166
rect 22093 20226 22159 20229
rect 24117 20226 24183 20229
rect 22093 20224 24183 20226
rect 22093 20168 22098 20224
rect 22154 20168 24122 20224
rect 24178 20168 24183 20224
rect 22093 20166 24183 20168
rect 22093 20163 22159 20166
rect 24117 20163 24183 20166
rect 20989 20090 21055 20093
rect 23473 20092 23539 20093
rect 20989 20088 23352 20090
rect 20989 20032 20994 20088
rect 21050 20032 23352 20088
rect 20989 20030 23352 20032
rect 20989 20027 21055 20030
rect 15745 19952 20914 19954
rect 15745 19896 15750 19952
rect 15806 19896 20914 19952
rect 15745 19894 20914 19896
rect 23292 19954 23352 20030
rect 23422 20028 23428 20092
rect 23492 20090 23539 20092
rect 23749 20090 23815 20093
rect 26325 20090 26391 20093
rect 23492 20088 23584 20090
rect 23534 20032 23584 20088
rect 23492 20030 23584 20032
rect 23749 20088 26391 20090
rect 23749 20032 23754 20088
rect 23810 20032 26330 20088
rect 26386 20032 26391 20088
rect 23749 20030 26391 20032
rect 23492 20028 23539 20030
rect 23473 20027 23539 20028
rect 23749 20027 23815 20030
rect 26325 20027 26391 20030
rect 24669 19954 24735 19957
rect 23292 19952 24735 19954
rect 23292 19896 24674 19952
rect 24730 19896 24735 19952
rect 23292 19894 24735 19896
rect 15745 19891 15811 19894
rect 24669 19891 24735 19894
rect 25497 19954 25563 19957
rect 27520 19954 28000 19984
rect 25497 19952 28000 19954
rect 25497 19896 25502 19952
rect 25558 19896 28000 19952
rect 25497 19894 28000 19896
rect 25497 19891 25563 19894
rect 27520 19864 28000 19894
rect 5390 19756 5396 19820
rect 5460 19818 5466 19820
rect 8385 19818 8451 19821
rect 5460 19816 8451 19818
rect 5460 19760 8390 19816
rect 8446 19760 8451 19816
rect 5460 19758 8451 19760
rect 5460 19756 5466 19758
rect 8385 19755 8451 19758
rect 9765 19818 9831 19821
rect 9990 19818 9996 19820
rect 9765 19816 9996 19818
rect 9765 19760 9770 19816
rect 9826 19760 9996 19816
rect 9765 19758 9996 19760
rect 9765 19755 9831 19758
rect 9990 19756 9996 19758
rect 10060 19818 10066 19820
rect 12341 19818 12407 19821
rect 23473 19818 23539 19821
rect 25221 19818 25287 19821
rect 25957 19820 26023 19821
rect 25957 19818 26004 19820
rect 10060 19758 12220 19818
rect 10060 19756 10066 19758
rect 0 19682 480 19712
rect 0 19622 5320 19682
rect 0 19592 480 19622
rect 5260 19410 5320 19622
rect 6310 19620 6316 19684
rect 6380 19682 6386 19684
rect 12014 19682 12020 19684
rect 6380 19622 12020 19682
rect 6380 19620 6386 19622
rect 12014 19620 12020 19622
rect 12084 19620 12090 19684
rect 12160 19682 12220 19758
rect 12341 19816 23539 19818
rect 12341 19760 12346 19816
rect 12402 19760 23478 19816
rect 23534 19760 23539 19816
rect 12341 19758 23539 19760
rect 12341 19755 12407 19758
rect 23473 19755 23539 19758
rect 23614 19816 25287 19818
rect 23614 19760 25226 19816
rect 25282 19760 25287 19816
rect 23614 19758 25287 19760
rect 25912 19816 26004 19818
rect 25912 19760 25962 19816
rect 25912 19758 26004 19760
rect 19333 19682 19399 19685
rect 23614 19682 23674 19758
rect 25221 19755 25287 19758
rect 25957 19756 26004 19758
rect 26068 19756 26074 19820
rect 25957 19755 26023 19756
rect 12160 19622 14842 19682
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 7189 19546 7255 19549
rect 10869 19546 10935 19549
rect 7189 19544 10935 19546
rect 7189 19488 7194 19544
rect 7250 19488 10874 19544
rect 10930 19488 10935 19544
rect 7189 19486 10935 19488
rect 7189 19483 7255 19486
rect 10869 19483 10935 19486
rect 11094 19484 11100 19548
rect 11164 19546 11170 19548
rect 11973 19546 12039 19549
rect 11164 19544 12039 19546
rect 11164 19488 11978 19544
rect 12034 19488 12039 19544
rect 11164 19486 12039 19488
rect 11164 19484 11170 19486
rect 11973 19483 12039 19486
rect 8293 19410 8359 19413
rect 5260 19408 8359 19410
rect 5260 19352 8298 19408
rect 8354 19352 8359 19408
rect 5260 19350 8359 19352
rect 8293 19347 8359 19350
rect 8845 19410 8911 19413
rect 14641 19410 14707 19413
rect 8845 19408 14707 19410
rect 8845 19352 8850 19408
rect 8906 19352 14646 19408
rect 14702 19352 14707 19408
rect 8845 19350 14707 19352
rect 14782 19410 14842 19622
rect 19333 19680 23674 19682
rect 19333 19624 19338 19680
rect 19394 19624 23674 19680
rect 19333 19622 23674 19624
rect 19333 19619 19399 19622
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 15377 19546 15443 19549
rect 21081 19546 21147 19549
rect 15377 19544 21147 19546
rect 15377 19488 15382 19544
rect 15438 19488 21086 19544
rect 21142 19488 21147 19544
rect 15377 19486 21147 19488
rect 15377 19483 15443 19486
rect 21081 19483 21147 19486
rect 22318 19484 22324 19548
rect 22388 19546 22394 19548
rect 24025 19546 24091 19549
rect 22388 19544 24091 19546
rect 22388 19488 24030 19544
rect 24086 19488 24091 19544
rect 22388 19486 24091 19488
rect 22388 19484 22394 19486
rect 24025 19483 24091 19486
rect 16113 19410 16179 19413
rect 14782 19408 16179 19410
rect 14782 19352 16118 19408
rect 16174 19352 16179 19408
rect 14782 19350 16179 19352
rect 8845 19347 8911 19350
rect 14641 19347 14707 19350
rect 16113 19347 16179 19350
rect 18873 19410 18939 19413
rect 24209 19410 24275 19413
rect 18873 19408 24275 19410
rect 18873 19352 18878 19408
rect 18934 19352 24214 19408
rect 24270 19352 24275 19408
rect 18873 19350 24275 19352
rect 18873 19347 18939 19350
rect 24209 19347 24275 19350
rect 24577 19410 24643 19413
rect 27520 19410 28000 19440
rect 24577 19408 28000 19410
rect 24577 19352 24582 19408
rect 24638 19352 28000 19408
rect 24577 19350 28000 19352
rect 24577 19347 24643 19350
rect 27520 19320 28000 19350
rect 2037 19274 2103 19277
rect 4153 19274 4219 19277
rect 4286 19274 4292 19276
rect 2037 19272 4292 19274
rect 2037 19216 2042 19272
rect 2098 19216 4158 19272
rect 4214 19216 4292 19272
rect 2037 19214 4292 19216
rect 2037 19211 2103 19214
rect 4153 19211 4219 19214
rect 4286 19212 4292 19214
rect 4356 19212 4362 19276
rect 5257 19274 5323 19277
rect 6821 19274 6887 19277
rect 5257 19272 6887 19274
rect 5257 19216 5262 19272
rect 5318 19216 6826 19272
rect 6882 19216 6887 19272
rect 5257 19214 6887 19216
rect 5257 19211 5323 19214
rect 6821 19211 6887 19214
rect 7005 19276 7071 19277
rect 7005 19272 7052 19276
rect 7116 19274 7122 19276
rect 7649 19274 7715 19277
rect 11237 19274 11303 19277
rect 15377 19274 15443 19277
rect 7005 19216 7010 19272
rect 7005 19212 7052 19216
rect 7116 19214 7162 19274
rect 7649 19272 11162 19274
rect 7649 19216 7654 19272
rect 7710 19216 11162 19272
rect 7649 19214 11162 19216
rect 7116 19212 7122 19214
rect 7005 19211 7071 19212
rect 7649 19211 7715 19214
rect 1945 19138 2011 19141
rect 2957 19138 3023 19141
rect 1945 19136 3023 19138
rect 1945 19080 1950 19136
rect 2006 19080 2962 19136
rect 3018 19080 3023 19136
rect 1945 19078 3023 19080
rect 1945 19075 2011 19078
rect 2957 19075 3023 19078
rect 5993 19138 6059 19141
rect 9765 19138 9831 19141
rect 5993 19136 9831 19138
rect 5993 19080 5998 19136
rect 6054 19080 9770 19136
rect 9826 19080 9831 19136
rect 5993 19078 9831 19080
rect 11102 19138 11162 19214
rect 11237 19272 15443 19274
rect 11237 19216 11242 19272
rect 11298 19216 15382 19272
rect 15438 19216 15443 19272
rect 11237 19214 15443 19216
rect 11237 19211 11303 19214
rect 15377 19211 15443 19214
rect 18045 19274 18111 19277
rect 20529 19274 20595 19277
rect 23013 19274 23079 19277
rect 18045 19272 23079 19274
rect 18045 19216 18050 19272
rect 18106 19216 20534 19272
rect 20590 19216 23018 19272
rect 23074 19216 23079 19272
rect 18045 19214 23079 19216
rect 18045 19211 18111 19214
rect 20529 19211 20595 19214
rect 23013 19211 23079 19214
rect 23422 19212 23428 19276
rect 23492 19274 23498 19276
rect 24669 19274 24735 19277
rect 23492 19272 24735 19274
rect 23492 19216 24674 19272
rect 24730 19216 24735 19272
rect 23492 19214 24735 19216
rect 23492 19212 23498 19214
rect 24669 19211 24735 19214
rect 11329 19138 11395 19141
rect 11102 19136 11395 19138
rect 11102 19080 11334 19136
rect 11390 19080 11395 19136
rect 11102 19078 11395 19080
rect 5993 19075 6059 19078
rect 9765 19075 9831 19078
rect 11329 19075 11395 19078
rect 11830 19076 11836 19140
rect 11900 19138 11906 19140
rect 12065 19138 12131 19141
rect 11900 19136 12131 19138
rect 11900 19080 12070 19136
rect 12126 19080 12131 19136
rect 11900 19078 12131 19080
rect 11900 19076 11906 19078
rect 12065 19075 12131 19078
rect 12198 19076 12204 19140
rect 12268 19138 12274 19140
rect 13629 19138 13695 19141
rect 12268 19136 13695 19138
rect 12268 19080 13634 19136
rect 13690 19080 13695 19136
rect 12268 19078 13695 19080
rect 12268 19076 12274 19078
rect 13629 19075 13695 19078
rect 14273 19138 14339 19141
rect 16941 19138 17007 19141
rect 14273 19136 17007 19138
rect 14273 19080 14278 19136
rect 14334 19080 16946 19136
rect 17002 19080 17007 19136
rect 14273 19078 17007 19080
rect 14273 19075 14339 19078
rect 16941 19075 17007 19078
rect 20989 19138 21055 19141
rect 24025 19138 24091 19141
rect 20989 19136 24091 19138
rect 20989 19080 20994 19136
rect 21050 19080 24030 19136
rect 24086 19080 24091 19136
rect 20989 19078 24091 19080
rect 20989 19075 21055 19078
rect 24025 19075 24091 19078
rect 24485 19138 24551 19141
rect 24894 19138 24900 19140
rect 24485 19136 24900 19138
rect 24485 19080 24490 19136
rect 24546 19080 24900 19136
rect 24485 19078 24900 19080
rect 24485 19075 24551 19078
rect 24894 19076 24900 19078
rect 24964 19076 24970 19140
rect 10277 19072 10597 19073
rect 0 19002 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 3417 19002 3483 19005
rect 0 19000 3483 19002
rect 0 18944 3422 19000
rect 3478 18944 3483 19000
rect 0 18942 3483 18944
rect 0 18912 480 18942
rect 3417 18939 3483 18942
rect 3785 19002 3851 19005
rect 5206 19002 5212 19004
rect 3785 19000 5212 19002
rect 3785 18944 3790 19000
rect 3846 18944 5212 19000
rect 3785 18942 5212 18944
rect 3785 18939 3851 18942
rect 5206 18940 5212 18942
rect 5276 18940 5282 19004
rect 7189 19002 7255 19005
rect 9489 19002 9555 19005
rect 7189 19000 9555 19002
rect 7189 18944 7194 19000
rect 7250 18944 9494 19000
rect 9550 18944 9555 19000
rect 7189 18942 9555 18944
rect 7189 18939 7255 18942
rect 9489 18939 9555 18942
rect 11646 18940 11652 19004
rect 11716 19002 11722 19004
rect 11973 19002 12039 19005
rect 11716 19000 12039 19002
rect 11716 18944 11978 19000
rect 12034 18944 12039 19000
rect 11716 18942 12039 18944
rect 11716 18940 11722 18942
rect 11973 18939 12039 18942
rect 12433 19002 12499 19005
rect 13261 19002 13327 19005
rect 18965 19002 19031 19005
rect 12433 19000 19031 19002
rect 12433 18944 12438 19000
rect 12494 18944 13266 19000
rect 13322 18944 18970 19000
rect 19026 18944 19031 19000
rect 12433 18942 19031 18944
rect 12433 18939 12499 18942
rect 13261 18939 13327 18942
rect 18965 18939 19031 18942
rect 20069 19000 20135 19005
rect 20069 18944 20074 19000
rect 20130 18944 20135 19000
rect 20069 18939 20135 18944
rect 20478 18940 20484 19004
rect 20548 19002 20554 19004
rect 21214 19002 21220 19004
rect 20548 18942 21220 19002
rect 20548 18940 20554 18942
rect 21214 18940 21220 18942
rect 21284 19002 21290 19004
rect 25221 19002 25287 19005
rect 21284 19000 25287 19002
rect 21284 18944 25226 19000
rect 25282 18944 25287 19000
rect 21284 18942 25287 18944
rect 21284 18940 21290 18942
rect 25221 18939 25287 18942
rect 1393 18866 1459 18869
rect 5993 18866 6059 18869
rect 1393 18864 6059 18866
rect 1393 18808 1398 18864
rect 1454 18808 5998 18864
rect 6054 18808 6059 18864
rect 1393 18806 6059 18808
rect 1393 18803 1459 18806
rect 5993 18803 6059 18806
rect 7005 18866 7071 18869
rect 7741 18866 7807 18869
rect 7005 18864 7807 18866
rect 7005 18808 7010 18864
rect 7066 18808 7746 18864
rect 7802 18808 7807 18864
rect 7005 18806 7807 18808
rect 7005 18803 7071 18806
rect 7741 18803 7807 18806
rect 8477 18866 8543 18869
rect 15101 18866 15167 18869
rect 18597 18866 18663 18869
rect 8477 18864 15026 18866
rect 8477 18808 8482 18864
rect 8538 18808 15026 18864
rect 8477 18806 15026 18808
rect 8477 18803 8543 18806
rect 2865 18730 2931 18733
rect 3785 18730 3851 18733
rect 12433 18730 12499 18733
rect 2865 18728 12499 18730
rect 2865 18672 2870 18728
rect 2926 18672 3790 18728
rect 3846 18672 12438 18728
rect 12494 18672 12499 18728
rect 2865 18670 12499 18672
rect 2865 18667 2931 18670
rect 3785 18667 3851 18670
rect 12433 18667 12499 18670
rect 12617 18730 12683 18733
rect 14825 18730 14891 18733
rect 12617 18728 14891 18730
rect 12617 18672 12622 18728
rect 12678 18672 14830 18728
rect 14886 18672 14891 18728
rect 12617 18670 14891 18672
rect 14966 18730 15026 18806
rect 15101 18864 18663 18866
rect 15101 18808 15106 18864
rect 15162 18808 18602 18864
rect 18658 18808 18663 18864
rect 15101 18806 18663 18808
rect 15101 18803 15167 18806
rect 18597 18803 18663 18806
rect 19609 18866 19675 18869
rect 20072 18866 20132 18939
rect 19609 18864 20132 18866
rect 19609 18808 19614 18864
rect 19670 18808 20132 18864
rect 19609 18806 20132 18808
rect 21449 18866 21515 18869
rect 25037 18866 25103 18869
rect 21449 18864 25103 18866
rect 21449 18808 21454 18864
rect 21510 18808 25042 18864
rect 25098 18808 25103 18864
rect 21449 18806 25103 18808
rect 19609 18803 19675 18806
rect 21449 18803 21515 18806
rect 25037 18803 25103 18806
rect 15837 18730 15903 18733
rect 17033 18730 17099 18733
rect 27520 18730 28000 18760
rect 14966 18728 16866 18730
rect 14966 18672 15842 18728
rect 15898 18672 16866 18728
rect 14966 18670 16866 18672
rect 12617 18667 12683 18670
rect 14825 18667 14891 18670
rect 15837 18667 15903 18670
rect 7373 18594 7439 18597
rect 12617 18594 12683 18597
rect 7373 18592 12683 18594
rect 7373 18536 7378 18592
rect 7434 18536 12622 18592
rect 12678 18536 12683 18592
rect 7373 18534 12683 18536
rect 16806 18594 16866 18670
rect 17033 18728 28000 18730
rect 17033 18672 17038 18728
rect 17094 18672 28000 18728
rect 17033 18670 28000 18672
rect 17033 18667 17099 18670
rect 27520 18640 28000 18670
rect 18505 18594 18571 18597
rect 16806 18592 18571 18594
rect 16806 18536 18510 18592
rect 18566 18536 18571 18592
rect 16806 18534 18571 18536
rect 7373 18531 7439 18534
rect 12617 18531 12683 18534
rect 18505 18531 18571 18534
rect 21357 18594 21423 18597
rect 23657 18594 23723 18597
rect 21357 18592 23723 18594
rect 21357 18536 21362 18592
rect 21418 18536 23662 18592
rect 23718 18536 23723 18592
rect 21357 18534 23723 18536
rect 21357 18531 21423 18534
rect 23657 18531 23723 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 11145 18458 11211 18461
rect 13261 18458 13327 18461
rect 11145 18456 13327 18458
rect 11145 18400 11150 18456
rect 11206 18400 13266 18456
rect 13322 18400 13327 18456
rect 11145 18398 13327 18400
rect 11145 18395 11211 18398
rect 13261 18395 13327 18398
rect 14590 18396 14596 18460
rect 14660 18458 14666 18460
rect 14733 18458 14799 18461
rect 14660 18456 14799 18458
rect 14660 18400 14738 18456
rect 14794 18400 14799 18456
rect 14660 18398 14799 18400
rect 14660 18396 14666 18398
rect 14733 18395 14799 18398
rect 15377 18458 15443 18461
rect 17125 18458 17191 18461
rect 21449 18458 21515 18461
rect 15377 18456 21515 18458
rect 15377 18400 15382 18456
rect 15438 18400 17130 18456
rect 17186 18400 21454 18456
rect 21510 18400 21515 18456
rect 15377 18398 21515 18400
rect 15377 18395 15443 18398
rect 17125 18395 17191 18398
rect 21449 18395 21515 18398
rect 0 18322 480 18352
rect 4061 18322 4127 18325
rect 0 18320 4127 18322
rect 0 18264 4066 18320
rect 4122 18264 4127 18320
rect 0 18262 4127 18264
rect 0 18232 480 18262
rect 4061 18259 4127 18262
rect 8937 18322 9003 18325
rect 11605 18322 11671 18325
rect 23473 18322 23539 18325
rect 8937 18320 10794 18322
rect 8937 18264 8942 18320
rect 8998 18264 10794 18320
rect 8937 18262 10794 18264
rect 8937 18259 9003 18262
rect 3233 18188 3299 18189
rect 3182 18124 3188 18188
rect 3252 18186 3299 18188
rect 3252 18184 3344 18186
rect 3294 18128 3344 18184
rect 3252 18126 3344 18128
rect 3252 18124 3299 18126
rect 3550 18124 3556 18188
rect 3620 18186 3626 18188
rect 6637 18186 6703 18189
rect 9806 18186 9812 18188
rect 3620 18184 6703 18186
rect 3620 18128 6642 18184
rect 6698 18128 6703 18184
rect 3620 18126 6703 18128
rect 3620 18124 3626 18126
rect 3233 18123 3299 18124
rect 6637 18123 6703 18126
rect 6870 18126 9812 18186
rect 2221 18052 2287 18053
rect 2773 18052 2839 18053
rect 2221 18048 2268 18052
rect 2332 18050 2338 18052
rect 2221 17992 2226 18048
rect 2221 17988 2268 17992
rect 2332 17990 2378 18050
rect 2773 18048 2820 18052
rect 2884 18050 2890 18052
rect 2773 17992 2778 18048
rect 2332 17988 2338 17990
rect 2773 17988 2820 17992
rect 2884 17990 2930 18050
rect 2884 17988 2890 17990
rect 5022 17988 5028 18052
rect 5092 18050 5098 18052
rect 6870 18050 6930 18126
rect 9806 18124 9812 18126
rect 9876 18124 9882 18188
rect 5092 17990 6930 18050
rect 5092 17988 5098 17990
rect 7046 17988 7052 18052
rect 7116 18050 7122 18052
rect 7833 18050 7899 18053
rect 7116 18048 7899 18050
rect 7116 17992 7838 18048
rect 7894 17992 7899 18048
rect 7116 17990 7899 17992
rect 7116 17988 7122 17990
rect 2221 17987 2287 17988
rect 2773 17987 2839 17988
rect 7833 17987 7899 17990
rect 8569 18050 8635 18053
rect 8937 18050 9003 18053
rect 8569 18048 9003 18050
rect 8569 17992 8574 18048
rect 8630 17992 8942 18048
rect 8998 17992 9003 18048
rect 8569 17990 9003 17992
rect 10734 18050 10794 18262
rect 11605 18320 23539 18322
rect 11605 18264 11610 18320
rect 11666 18264 23478 18320
rect 23534 18264 23539 18320
rect 11605 18262 23539 18264
rect 11605 18259 11671 18262
rect 23473 18259 23539 18262
rect 24117 18322 24183 18325
rect 26233 18322 26299 18325
rect 24117 18320 26299 18322
rect 24117 18264 24122 18320
rect 24178 18264 26238 18320
rect 26294 18264 26299 18320
rect 24117 18262 26299 18264
rect 24117 18259 24183 18262
rect 26233 18259 26299 18262
rect 11329 18186 11395 18189
rect 23657 18186 23723 18189
rect 27520 18186 28000 18216
rect 11329 18184 23723 18186
rect 11329 18128 11334 18184
rect 11390 18128 23662 18184
rect 23718 18128 23723 18184
rect 11329 18126 23723 18128
rect 11329 18123 11395 18126
rect 23657 18123 23723 18126
rect 25638 18126 28000 18186
rect 12525 18050 12591 18053
rect 16205 18052 16271 18053
rect 16205 18050 16252 18052
rect 10734 18048 12591 18050
rect 10734 17992 12530 18048
rect 12586 17992 12591 18048
rect 10734 17990 12591 17992
rect 16160 18048 16252 18050
rect 16160 17992 16210 18048
rect 16160 17990 16252 17992
rect 8569 17987 8635 17990
rect 8937 17987 9003 17990
rect 12525 17987 12591 17990
rect 16205 17988 16252 17990
rect 16316 17988 16322 18052
rect 21081 18050 21147 18053
rect 21398 18050 21404 18052
rect 21081 18048 21404 18050
rect 21081 17992 21086 18048
rect 21142 17992 21404 18048
rect 21081 17990 21404 17992
rect 16205 17987 16271 17988
rect 21081 17987 21147 17990
rect 21398 17988 21404 17990
rect 21468 17988 21474 18052
rect 21541 18050 21607 18053
rect 21766 18050 21772 18052
rect 21541 18048 21772 18050
rect 21541 17992 21546 18048
rect 21602 17992 21772 18048
rect 21541 17990 21772 17992
rect 21541 17987 21607 17990
rect 21766 17988 21772 17990
rect 21836 17988 21842 18052
rect 22134 17988 22140 18052
rect 22204 18050 22210 18052
rect 23657 18050 23723 18053
rect 22204 18048 23723 18050
rect 22204 17992 23662 18048
rect 23718 17992 23723 18048
rect 22204 17990 23723 17992
rect 22204 17988 22210 17990
rect 23657 17987 23723 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 25638 17917 25698 18126
rect 27520 18096 28000 18126
rect 2589 17916 2655 17917
rect 2589 17914 2636 17916
rect 2508 17912 2636 17914
rect 2700 17914 2706 17916
rect 3049 17914 3115 17917
rect 2700 17912 3115 17914
rect 2508 17856 2594 17912
rect 2700 17856 3054 17912
rect 3110 17856 3115 17912
rect 2508 17854 2636 17856
rect 2589 17852 2636 17854
rect 2700 17854 3115 17856
rect 2700 17852 2706 17854
rect 2589 17851 2655 17852
rect 3049 17851 3115 17854
rect 3509 17914 3575 17917
rect 6310 17914 6316 17916
rect 3509 17912 6316 17914
rect 3509 17856 3514 17912
rect 3570 17856 6316 17912
rect 3509 17854 6316 17856
rect 3509 17851 3575 17854
rect 6310 17852 6316 17854
rect 6380 17852 6386 17916
rect 7782 17852 7788 17916
rect 7852 17914 7858 17916
rect 8518 17914 8524 17916
rect 7852 17854 8524 17914
rect 7852 17852 7858 17854
rect 8518 17852 8524 17854
rect 8588 17852 8594 17916
rect 12801 17914 12867 17917
rect 13629 17914 13695 17917
rect 18689 17914 18755 17917
rect 12801 17912 13002 17914
rect 12801 17856 12806 17912
rect 12862 17856 13002 17912
rect 12801 17854 13002 17856
rect 12801 17851 12867 17854
rect 2497 17778 2563 17781
rect 4838 17778 4844 17780
rect 2497 17776 4844 17778
rect 2497 17720 2502 17776
rect 2558 17720 4844 17776
rect 2497 17718 4844 17720
rect 2497 17715 2563 17718
rect 4838 17716 4844 17718
rect 4908 17778 4914 17780
rect 6637 17778 6703 17781
rect 4908 17776 6703 17778
rect 4908 17720 6642 17776
rect 6698 17720 6703 17776
rect 4908 17718 6703 17720
rect 4908 17716 4914 17718
rect 6637 17715 6703 17718
rect 6821 17778 6887 17781
rect 10317 17778 10383 17781
rect 12525 17778 12591 17781
rect 6821 17776 10242 17778
rect 6821 17720 6826 17776
rect 6882 17720 10242 17776
rect 6821 17718 10242 17720
rect 6821 17715 6887 17718
rect 0 17642 480 17672
rect 9857 17642 9923 17645
rect 0 17640 9923 17642
rect 0 17584 9862 17640
rect 9918 17584 9923 17640
rect 0 17582 9923 17584
rect 0 17552 480 17582
rect 9857 17579 9923 17582
rect 10182 17506 10242 17718
rect 10317 17776 12591 17778
rect 10317 17720 10322 17776
rect 10378 17720 12530 17776
rect 12586 17720 12591 17776
rect 10317 17718 12591 17720
rect 10317 17715 10383 17718
rect 12525 17715 12591 17718
rect 12942 17642 13002 17854
rect 13629 17912 18755 17914
rect 13629 17856 13634 17912
rect 13690 17856 18694 17912
rect 18750 17856 18755 17912
rect 13629 17854 18755 17856
rect 13629 17851 13695 17854
rect 18689 17851 18755 17854
rect 20662 17852 20668 17916
rect 20732 17914 20738 17916
rect 24117 17914 24183 17917
rect 20732 17912 24183 17914
rect 20732 17856 24122 17912
rect 24178 17856 24183 17912
rect 20732 17854 24183 17856
rect 20732 17852 20738 17854
rect 24117 17851 24183 17854
rect 25589 17912 25698 17917
rect 25589 17856 25594 17912
rect 25650 17856 25698 17912
rect 25589 17854 25698 17856
rect 25589 17851 25655 17854
rect 13169 17778 13235 17781
rect 15837 17778 15903 17781
rect 13169 17776 15903 17778
rect 13169 17720 13174 17776
rect 13230 17720 15842 17776
rect 15898 17720 15903 17776
rect 13169 17718 15903 17720
rect 13169 17715 13235 17718
rect 13629 17642 13695 17645
rect 12942 17640 13695 17642
rect 12942 17584 13634 17640
rect 13690 17584 13695 17640
rect 12942 17582 13695 17584
rect 13629 17579 13695 17582
rect 14782 17509 14842 17718
rect 15837 17715 15903 17718
rect 18137 17778 18203 17781
rect 24393 17778 24459 17781
rect 18137 17776 24459 17778
rect 18137 17720 18142 17776
rect 18198 17720 24398 17776
rect 24454 17720 24459 17776
rect 18137 17718 24459 17720
rect 18137 17715 18203 17718
rect 24393 17715 24459 17718
rect 16614 17580 16620 17644
rect 16684 17642 16690 17644
rect 16941 17642 17007 17645
rect 16684 17640 17007 17642
rect 16684 17584 16946 17640
rect 17002 17584 17007 17640
rect 16684 17582 17007 17584
rect 16684 17580 16690 17582
rect 16941 17579 17007 17582
rect 18597 17642 18663 17645
rect 23749 17642 23815 17645
rect 18597 17640 23815 17642
rect 18597 17584 18602 17640
rect 18658 17584 23754 17640
rect 23810 17584 23815 17640
rect 18597 17582 23815 17584
rect 18597 17579 18663 17582
rect 23749 17579 23815 17582
rect 24025 17642 24091 17645
rect 27520 17642 28000 17672
rect 24025 17640 28000 17642
rect 24025 17584 24030 17640
rect 24086 17584 28000 17640
rect 24025 17582 28000 17584
rect 24025 17579 24091 17582
rect 27520 17552 28000 17582
rect 14038 17506 14044 17508
rect 10182 17446 14044 17506
rect 14038 17444 14044 17446
rect 14108 17444 14114 17508
rect 14733 17504 14842 17509
rect 18781 17506 18847 17509
rect 22553 17506 22619 17509
rect 14733 17448 14738 17504
rect 14794 17448 14842 17504
rect 14733 17446 14842 17448
rect 15334 17446 18706 17506
rect 14733 17443 14799 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 6637 17370 6703 17373
rect 10726 17370 10732 17372
rect 6637 17368 10732 17370
rect 6637 17312 6642 17368
rect 6698 17312 10732 17368
rect 6637 17310 10732 17312
rect 6637 17307 6703 17310
rect 10726 17308 10732 17310
rect 10796 17308 10802 17372
rect 11329 17370 11395 17373
rect 11462 17370 11468 17372
rect 11329 17368 11468 17370
rect 11329 17312 11334 17368
rect 11390 17312 11468 17368
rect 11329 17310 11468 17312
rect 11329 17307 11395 17310
rect 11462 17308 11468 17310
rect 11532 17308 11538 17372
rect 2037 17234 2103 17237
rect 12157 17234 12223 17237
rect 2037 17232 12223 17234
rect 2037 17176 2042 17232
rect 2098 17176 12162 17232
rect 12218 17176 12223 17232
rect 2037 17174 12223 17176
rect 2037 17171 2103 17174
rect 12157 17171 12223 17174
rect 14917 17234 14983 17237
rect 15334 17234 15394 17446
rect 16021 17370 16087 17373
rect 18229 17370 18295 17373
rect 16021 17368 18295 17370
rect 16021 17312 16026 17368
rect 16082 17312 18234 17368
rect 18290 17312 18295 17368
rect 16021 17310 18295 17312
rect 18646 17370 18706 17446
rect 18781 17504 22619 17506
rect 18781 17448 18786 17504
rect 18842 17448 22558 17504
rect 22614 17448 22619 17504
rect 18781 17446 22619 17448
rect 18781 17443 18847 17446
rect 22553 17443 22619 17446
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 19006 17370 19012 17372
rect 18646 17310 19012 17370
rect 16021 17307 16087 17310
rect 18229 17307 18295 17310
rect 19006 17308 19012 17310
rect 19076 17370 19082 17372
rect 19517 17370 19583 17373
rect 19076 17368 19583 17370
rect 19076 17312 19522 17368
rect 19578 17312 19583 17368
rect 19076 17310 19583 17312
rect 19076 17308 19082 17310
rect 19517 17307 19583 17310
rect 19885 17370 19951 17373
rect 23933 17370 23999 17373
rect 19885 17368 23999 17370
rect 19885 17312 19890 17368
rect 19946 17312 23938 17368
rect 23994 17312 23999 17368
rect 19885 17310 23999 17312
rect 19885 17307 19951 17310
rect 23933 17307 23999 17310
rect 14917 17232 15394 17234
rect 14917 17176 14922 17232
rect 14978 17176 15394 17232
rect 14917 17174 15394 17176
rect 15929 17234 15995 17237
rect 24669 17234 24735 17237
rect 15929 17232 24735 17234
rect 15929 17176 15934 17232
rect 15990 17176 24674 17232
rect 24730 17176 24735 17232
rect 15929 17174 24735 17176
rect 14917 17171 14983 17174
rect 15929 17171 15995 17174
rect 24669 17171 24735 17174
rect 3141 17098 3207 17101
rect 4797 17098 4863 17101
rect 3141 17096 4863 17098
rect 3141 17040 3146 17096
rect 3202 17040 4802 17096
rect 4858 17040 4863 17096
rect 3141 17038 4863 17040
rect 3141 17035 3207 17038
rect 4797 17035 4863 17038
rect 5625 17098 5691 17101
rect 12065 17098 12131 17101
rect 17585 17098 17651 17101
rect 5625 17096 12131 17098
rect 5625 17040 5630 17096
rect 5686 17040 12070 17096
rect 12126 17040 12131 17096
rect 5625 17038 12131 17040
rect 5625 17035 5691 17038
rect 12065 17035 12131 17038
rect 12206 17096 17651 17098
rect 12206 17040 17590 17096
rect 17646 17040 17651 17096
rect 12206 17038 17651 17040
rect 0 16962 480 16992
rect 3601 16962 3667 16965
rect 0 16960 3667 16962
rect 0 16904 3606 16960
rect 3662 16904 3667 16960
rect 0 16902 3667 16904
rect 0 16872 480 16902
rect 3601 16899 3667 16902
rect 8109 16962 8175 16965
rect 8845 16962 8911 16965
rect 8109 16960 8911 16962
rect 8109 16904 8114 16960
rect 8170 16904 8850 16960
rect 8906 16904 8911 16960
rect 8109 16902 8911 16904
rect 8109 16899 8175 16902
rect 8845 16899 8911 16902
rect 10726 16900 10732 16964
rect 10796 16962 10802 16964
rect 12206 16962 12266 17038
rect 17585 17035 17651 17038
rect 19374 17036 19380 17100
rect 19444 17098 19450 17100
rect 20294 17098 20300 17100
rect 19444 17038 20300 17098
rect 19444 17036 19450 17038
rect 20294 17036 20300 17038
rect 20364 17036 20370 17100
rect 20529 17098 20595 17101
rect 21449 17098 21515 17101
rect 20529 17096 21515 17098
rect 20529 17040 20534 17096
rect 20590 17040 21454 17096
rect 21510 17040 21515 17096
rect 20529 17038 21515 17040
rect 20529 17035 20595 17038
rect 21449 17035 21515 17038
rect 21766 17036 21772 17100
rect 21836 17098 21842 17100
rect 22093 17098 22159 17101
rect 21836 17096 22159 17098
rect 21836 17040 22098 17096
rect 22154 17040 22159 17096
rect 21836 17038 22159 17040
rect 21836 17036 21842 17038
rect 22093 17035 22159 17038
rect 23565 17100 23631 17101
rect 23565 17096 23612 17100
rect 23676 17098 23682 17100
rect 24209 17098 24275 17101
rect 24710 17098 24716 17100
rect 23565 17040 23570 17096
rect 23565 17036 23612 17040
rect 23676 17038 23722 17098
rect 24209 17096 24716 17098
rect 24209 17040 24214 17096
rect 24270 17040 24716 17096
rect 24209 17038 24716 17040
rect 23676 17036 23682 17038
rect 23565 17035 23631 17036
rect 24209 17035 24275 17038
rect 24710 17036 24716 17038
rect 24780 17036 24786 17100
rect 25865 17098 25931 17101
rect 27520 17098 28000 17128
rect 25865 17096 28000 17098
rect 25865 17040 25870 17096
rect 25926 17040 28000 17096
rect 25865 17038 28000 17040
rect 25865 17035 25931 17038
rect 27520 17008 28000 17038
rect 10796 16902 12266 16962
rect 12433 16962 12499 16965
rect 15009 16962 15075 16965
rect 12433 16960 15075 16962
rect 12433 16904 12438 16960
rect 12494 16904 15014 16960
rect 15070 16904 15075 16960
rect 12433 16902 15075 16904
rect 10796 16900 10802 16902
rect 12433 16899 12499 16902
rect 15009 16899 15075 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 1393 16826 1459 16829
rect 6913 16826 6979 16829
rect 1393 16824 6979 16826
rect 1393 16768 1398 16824
rect 1454 16768 6918 16824
rect 6974 16768 6979 16824
rect 1393 16766 6979 16768
rect 1393 16763 1459 16766
rect 6913 16763 6979 16766
rect 15469 16826 15535 16829
rect 26325 16826 26391 16829
rect 15469 16824 19488 16826
rect 15469 16768 15474 16824
rect 15530 16768 19488 16824
rect 15469 16766 19488 16768
rect 15469 16763 15535 16766
rect 1894 16628 1900 16692
rect 1964 16690 1970 16692
rect 2129 16690 2195 16693
rect 1964 16688 2195 16690
rect 1964 16632 2134 16688
rect 2190 16632 2195 16688
rect 1964 16630 2195 16632
rect 1964 16628 1970 16630
rect 2129 16627 2195 16630
rect 4061 16690 4127 16693
rect 6913 16690 6979 16693
rect 4061 16688 6979 16690
rect 4061 16632 4066 16688
rect 4122 16632 6918 16688
rect 6974 16632 6979 16688
rect 4061 16630 6979 16632
rect 4061 16627 4127 16630
rect 6913 16627 6979 16630
rect 9806 16628 9812 16692
rect 9876 16690 9882 16692
rect 10317 16690 10383 16693
rect 9876 16688 10383 16690
rect 9876 16632 10322 16688
rect 10378 16632 10383 16688
rect 9876 16630 10383 16632
rect 9876 16628 9882 16630
rect 10317 16627 10383 16630
rect 10869 16690 10935 16693
rect 11278 16690 11284 16692
rect 10869 16688 11284 16690
rect 10869 16632 10874 16688
rect 10930 16632 11284 16688
rect 10869 16630 11284 16632
rect 10869 16627 10935 16630
rect 11278 16628 11284 16630
rect 11348 16628 11354 16692
rect 11881 16690 11947 16693
rect 17033 16690 17099 16693
rect 11881 16688 17099 16690
rect 11881 16632 11886 16688
rect 11942 16632 17038 16688
rect 17094 16632 17099 16688
rect 11881 16630 17099 16632
rect 19428 16690 19488 16766
rect 20072 16824 26391 16826
rect 20072 16768 26330 16824
rect 26386 16768 26391 16824
rect 20072 16766 26391 16768
rect 20072 16724 20132 16766
rect 26325 16763 26391 16766
rect 19980 16690 20132 16724
rect 19428 16664 20132 16690
rect 22185 16690 22251 16693
rect 22318 16690 22324 16692
rect 22185 16688 22324 16690
rect 19428 16630 20040 16664
rect 22185 16632 22190 16688
rect 22246 16632 22324 16688
rect 22185 16630 22324 16632
rect 11881 16627 11947 16630
rect 17033 16627 17099 16630
rect 22185 16627 22251 16630
rect 22318 16628 22324 16630
rect 22388 16628 22394 16692
rect 23197 16690 23263 16693
rect 23197 16688 23490 16690
rect 23197 16632 23202 16688
rect 23258 16632 23490 16688
rect 23197 16630 23490 16632
rect 23197 16627 23263 16630
rect 2865 16554 2931 16557
rect 4470 16554 4476 16556
rect 2865 16552 4476 16554
rect 2865 16496 2870 16552
rect 2926 16496 4476 16552
rect 2865 16494 4476 16496
rect 2865 16491 2931 16494
rect 4470 16492 4476 16494
rect 4540 16492 4546 16556
rect 8293 16554 8359 16557
rect 12157 16554 12223 16557
rect 8293 16552 12223 16554
rect 8293 16496 8298 16552
rect 8354 16496 12162 16552
rect 12218 16496 12223 16552
rect 8293 16494 12223 16496
rect 8293 16491 8359 16494
rect 12157 16491 12223 16494
rect 16757 16554 16823 16557
rect 20989 16554 21055 16557
rect 16757 16552 21055 16554
rect 16757 16496 16762 16552
rect 16818 16496 20994 16552
rect 21050 16496 21055 16552
rect 16757 16494 21055 16496
rect 23430 16554 23490 16630
rect 23657 16554 23723 16557
rect 23430 16552 23723 16554
rect 23430 16496 23662 16552
rect 23718 16496 23723 16552
rect 23430 16494 23723 16496
rect 16757 16491 16823 16494
rect 20989 16491 21055 16494
rect 23657 16491 23723 16494
rect 25681 16554 25747 16557
rect 27520 16554 28000 16584
rect 25681 16552 28000 16554
rect 25681 16496 25686 16552
rect 25742 16496 28000 16552
rect 25681 16494 28000 16496
rect 25681 16491 25747 16494
rect 27520 16464 28000 16494
rect 6637 16418 6703 16421
rect 9305 16418 9371 16421
rect 10726 16418 10732 16420
rect 6637 16416 10732 16418
rect 6637 16360 6642 16416
rect 6698 16360 9310 16416
rect 9366 16360 10732 16416
rect 6637 16358 10732 16360
rect 6637 16355 6703 16358
rect 9305 16355 9371 16358
rect 10726 16356 10732 16358
rect 10796 16356 10802 16420
rect 10910 16356 10916 16420
rect 10980 16418 10986 16420
rect 14181 16418 14247 16421
rect 10980 16416 14247 16418
rect 10980 16360 14186 16416
rect 14242 16360 14247 16416
rect 10980 16358 14247 16360
rect 10980 16356 10986 16358
rect 14181 16355 14247 16358
rect 18781 16418 18847 16421
rect 19517 16418 19583 16421
rect 18781 16416 19583 16418
rect 18781 16360 18786 16416
rect 18842 16360 19522 16416
rect 19578 16360 19583 16416
rect 18781 16358 19583 16360
rect 18781 16355 18847 16358
rect 19517 16355 19583 16358
rect 5610 16352 5930 16353
rect 0 16282 480 16312
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16222 5458 16282
rect 0 16192 480 16222
rect 1393 16010 1459 16013
rect 4245 16010 4311 16013
rect 1393 16008 4311 16010
rect 1393 15952 1398 16008
rect 1454 15952 4250 16008
rect 4306 15952 4311 16008
rect 1393 15950 4311 15952
rect 5398 16010 5458 16222
rect 8150 16220 8156 16284
rect 8220 16282 8226 16284
rect 13629 16282 13695 16285
rect 8220 16280 13695 16282
rect 8220 16224 13634 16280
rect 13690 16224 13695 16280
rect 8220 16222 13695 16224
rect 8220 16220 8226 16222
rect 13629 16219 13695 16222
rect 15377 16282 15443 16285
rect 20069 16282 20135 16285
rect 23473 16282 23539 16285
rect 15377 16280 20135 16282
rect 15377 16224 15382 16280
rect 15438 16224 20074 16280
rect 20130 16224 20135 16280
rect 15377 16222 20135 16224
rect 15377 16219 15443 16222
rect 20069 16219 20135 16222
rect 20256 16280 23539 16282
rect 20256 16224 23478 16280
rect 23534 16224 23539 16280
rect 20256 16222 23539 16224
rect 9857 16146 9923 16149
rect 12525 16146 12591 16149
rect 9857 16144 12591 16146
rect 9857 16088 9862 16144
rect 9918 16088 12530 16144
rect 12586 16088 12591 16144
rect 9857 16086 12591 16088
rect 9857 16083 9923 16086
rect 12525 16083 12591 16086
rect 12709 16146 12775 16149
rect 15469 16146 15535 16149
rect 17861 16146 17927 16149
rect 12709 16144 17927 16146
rect 12709 16088 12714 16144
rect 12770 16088 15474 16144
rect 15530 16088 17866 16144
rect 17922 16088 17927 16144
rect 12709 16086 17927 16088
rect 12709 16083 12775 16086
rect 15469 16083 15535 16086
rect 17861 16083 17927 16086
rect 18137 16146 18203 16149
rect 19057 16146 19123 16149
rect 20256 16146 20316 16222
rect 23473 16219 23539 16222
rect 18137 16144 20316 16146
rect 18137 16088 18142 16144
rect 18198 16088 19062 16144
rect 19118 16088 20316 16144
rect 18137 16086 20316 16088
rect 18137 16083 18203 16086
rect 19057 16083 19123 16086
rect 20662 16084 20668 16148
rect 20732 16146 20738 16148
rect 24025 16146 24091 16149
rect 20732 16144 24091 16146
rect 20732 16088 24030 16144
rect 24086 16088 24091 16144
rect 20732 16086 24091 16088
rect 20732 16084 20738 16086
rect 24025 16083 24091 16086
rect 9765 16010 9831 16013
rect 16205 16010 16271 16013
rect 5398 16008 9831 16010
rect 5398 15952 9770 16008
rect 9826 15952 9831 16008
rect 5398 15950 9831 15952
rect 1393 15947 1459 15950
rect 4245 15947 4311 15950
rect 9765 15947 9831 15950
rect 9998 16008 16271 16010
rect 9998 15952 16210 16008
rect 16266 15952 16271 16008
rect 9998 15950 16271 15952
rect 7097 15874 7163 15877
rect 1166 15872 7163 15874
rect 1166 15816 7102 15872
rect 7158 15816 7163 15872
rect 1166 15814 7163 15816
rect 0 15602 480 15632
rect 1166 15602 1226 15814
rect 7097 15811 7163 15814
rect 7373 15874 7439 15877
rect 9998 15874 10058 15950
rect 16205 15947 16271 15950
rect 19333 16010 19399 16013
rect 24209 16010 24275 16013
rect 19333 16008 24275 16010
rect 19333 15952 19338 16008
rect 19394 15952 24214 16008
rect 24270 15952 24275 16008
rect 19333 15950 24275 15952
rect 19333 15947 19399 15950
rect 24209 15947 24275 15950
rect 25405 16010 25471 16013
rect 27520 16010 28000 16040
rect 25405 16008 28000 16010
rect 25405 15952 25410 16008
rect 25466 15952 28000 16008
rect 25405 15950 28000 15952
rect 25405 15947 25471 15950
rect 27520 15920 28000 15950
rect 7373 15872 10058 15874
rect 7373 15816 7378 15872
rect 7434 15816 10058 15872
rect 7373 15814 10058 15816
rect 7373 15811 7439 15814
rect 10726 15812 10732 15876
rect 10796 15874 10802 15876
rect 14365 15874 14431 15877
rect 10796 15872 14431 15874
rect 10796 15816 14370 15872
rect 14426 15816 14431 15872
rect 10796 15814 14431 15816
rect 10796 15812 10802 15814
rect 14365 15811 14431 15814
rect 14917 15874 14983 15877
rect 16757 15874 16823 15877
rect 24025 15876 24091 15877
rect 14917 15872 16823 15874
rect 14917 15816 14922 15872
rect 14978 15816 16762 15872
rect 16818 15816 16823 15872
rect 14917 15814 16823 15816
rect 14917 15811 14983 15814
rect 16757 15811 16823 15814
rect 21398 15812 21404 15876
rect 21468 15874 21474 15876
rect 21950 15874 21956 15876
rect 21468 15814 21956 15874
rect 21468 15812 21474 15814
rect 21950 15812 21956 15814
rect 22020 15812 22026 15876
rect 23974 15874 23980 15876
rect 23934 15814 23980 15874
rect 24044 15872 24091 15876
rect 24086 15816 24091 15872
rect 23974 15812 23980 15814
rect 24044 15812 24091 15816
rect 24025 15811 24091 15812
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 2497 15738 2563 15741
rect 4838 15738 4844 15740
rect 2497 15736 4844 15738
rect 2497 15680 2502 15736
rect 2558 15680 4844 15736
rect 2497 15678 4844 15680
rect 2497 15675 2563 15678
rect 4838 15676 4844 15678
rect 4908 15738 4914 15740
rect 5390 15738 5396 15740
rect 4908 15678 5396 15738
rect 4908 15676 4914 15678
rect 5390 15676 5396 15678
rect 5460 15676 5466 15740
rect 6729 15738 6795 15741
rect 9397 15738 9463 15741
rect 9581 15740 9647 15741
rect 9581 15738 9628 15740
rect 6729 15736 9463 15738
rect 6729 15680 6734 15736
rect 6790 15680 9402 15736
rect 9458 15680 9463 15736
rect 6729 15678 9463 15680
rect 9540 15736 9628 15738
rect 9540 15680 9586 15736
rect 9540 15678 9628 15680
rect 6729 15675 6795 15678
rect 9397 15675 9463 15678
rect 9581 15676 9628 15678
rect 9692 15676 9698 15740
rect 10869 15738 10935 15741
rect 13721 15738 13787 15741
rect 15653 15738 15719 15741
rect 10869 15736 12128 15738
rect 10869 15680 10874 15736
rect 10930 15680 12128 15736
rect 10869 15678 12128 15680
rect 9581 15675 9647 15676
rect 10869 15675 10935 15678
rect 0 15542 1226 15602
rect 1393 15602 1459 15605
rect 9949 15602 10015 15605
rect 1393 15600 10015 15602
rect 1393 15544 1398 15600
rect 1454 15544 9954 15600
rect 10010 15544 10015 15600
rect 1393 15542 10015 15544
rect 12068 15602 12128 15678
rect 13721 15736 15719 15738
rect 13721 15680 13726 15736
rect 13782 15680 15658 15736
rect 15714 15680 15719 15736
rect 13721 15678 15719 15680
rect 13721 15675 13787 15678
rect 15653 15675 15719 15678
rect 20069 15738 20135 15741
rect 24853 15738 24919 15741
rect 20069 15736 24919 15738
rect 20069 15680 20074 15736
rect 20130 15680 24858 15736
rect 24914 15680 24919 15736
rect 20069 15678 24919 15680
rect 20069 15675 20135 15678
rect 24853 15675 24919 15678
rect 19057 15602 19123 15605
rect 19425 15602 19491 15605
rect 12068 15600 19491 15602
rect 12068 15544 19062 15600
rect 19118 15544 19430 15600
rect 19486 15544 19491 15600
rect 12068 15542 19491 15544
rect 0 15512 480 15542
rect 1393 15539 1459 15542
rect 9949 15539 10015 15542
rect 19057 15539 19123 15542
rect 19425 15539 19491 15542
rect 22553 15602 22619 15605
rect 22870 15602 22876 15604
rect 22553 15600 22876 15602
rect 22553 15544 22558 15600
rect 22614 15544 22876 15600
rect 22553 15542 22876 15544
rect 22553 15539 22619 15542
rect 22870 15540 22876 15542
rect 22940 15540 22946 15604
rect 3417 15466 3483 15469
rect 7373 15466 7439 15469
rect 3417 15464 7439 15466
rect 3417 15408 3422 15464
rect 3478 15408 7378 15464
rect 7434 15408 7439 15464
rect 3417 15406 7439 15408
rect 3417 15403 3483 15406
rect 7373 15403 7439 15406
rect 9949 15466 10015 15469
rect 15837 15466 15903 15469
rect 9949 15464 15903 15466
rect 9949 15408 9954 15464
rect 10010 15408 15842 15464
rect 15898 15408 15903 15464
rect 9949 15406 15903 15408
rect 9949 15403 10015 15406
rect 15837 15403 15903 15406
rect 16849 15466 16915 15469
rect 18321 15466 18387 15469
rect 16849 15464 18387 15466
rect 16849 15408 16854 15464
rect 16910 15408 18326 15464
rect 18382 15408 18387 15464
rect 16849 15406 18387 15408
rect 16849 15403 16915 15406
rect 18321 15403 18387 15406
rect 20713 15466 20779 15469
rect 27520 15466 28000 15496
rect 20713 15464 28000 15466
rect 20713 15408 20718 15464
rect 20774 15408 28000 15464
rect 20713 15406 28000 15408
rect 20713 15403 20779 15406
rect 27520 15376 28000 15406
rect 6085 15330 6151 15333
rect 7557 15330 7623 15333
rect 14089 15330 14155 15333
rect 6085 15328 14155 15330
rect 6085 15272 6090 15328
rect 6146 15272 7562 15328
rect 7618 15272 14094 15328
rect 14150 15272 14155 15328
rect 6085 15270 14155 15272
rect 6085 15267 6151 15270
rect 7557 15267 7623 15270
rect 14089 15267 14155 15270
rect 15653 15330 15719 15333
rect 18137 15330 18203 15333
rect 15653 15328 18203 15330
rect 15653 15272 15658 15328
rect 15714 15272 18142 15328
rect 18198 15272 18203 15328
rect 15653 15270 18203 15272
rect 15653 15267 15719 15270
rect 18137 15267 18203 15270
rect 18965 15330 19031 15333
rect 23013 15330 23079 15333
rect 18965 15328 23079 15330
rect 18965 15272 18970 15328
rect 19026 15272 23018 15328
rect 23074 15272 23079 15328
rect 18965 15270 23079 15272
rect 18965 15267 19031 15270
rect 23013 15267 23079 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 6637 15194 6703 15197
rect 7833 15194 7899 15197
rect 9765 15194 9831 15197
rect 6637 15192 9831 15194
rect 6637 15136 6642 15192
rect 6698 15136 7838 15192
rect 7894 15136 9770 15192
rect 9826 15136 9831 15192
rect 6637 15134 9831 15136
rect 6637 15131 6703 15134
rect 7833 15131 7899 15134
rect 9765 15131 9831 15134
rect 12709 15194 12775 15197
rect 14641 15194 14707 15197
rect 23933 15194 23999 15197
rect 12709 15192 14707 15194
rect 12709 15136 12714 15192
rect 12770 15136 14646 15192
rect 14702 15136 14707 15192
rect 12709 15134 14707 15136
rect 12709 15131 12775 15134
rect 14641 15131 14707 15134
rect 15334 15192 23999 15194
rect 15334 15136 23938 15192
rect 23994 15136 23999 15192
rect 15334 15134 23999 15136
rect 3601 15058 3667 15061
rect 6913 15058 6979 15061
rect 3601 15056 6979 15058
rect 3601 15000 3606 15056
rect 3662 15000 6918 15056
rect 6974 15000 6979 15056
rect 3601 14998 6979 15000
rect 3601 14995 3667 14998
rect 6913 14995 6979 14998
rect 9489 15058 9555 15061
rect 15193 15058 15259 15061
rect 15334 15058 15394 15134
rect 23933 15131 23999 15134
rect 9489 15056 15394 15058
rect 9489 15000 9494 15056
rect 9550 15000 15198 15056
rect 15254 15000 15394 15056
rect 9489 14998 15394 15000
rect 19977 15058 20043 15061
rect 20662 15058 20668 15060
rect 19977 15056 20668 15058
rect 19977 15000 19982 15056
rect 20038 15000 20668 15056
rect 19977 14998 20668 15000
rect 9489 14995 9555 14998
rect 15193 14995 15259 14998
rect 19977 14995 20043 14998
rect 20662 14996 20668 14998
rect 20732 14996 20738 15060
rect 21081 15058 21147 15061
rect 21357 15058 21423 15061
rect 21081 15056 21423 15058
rect 21081 15000 21086 15056
rect 21142 15000 21362 15056
rect 21418 15000 21423 15056
rect 21081 14998 21423 15000
rect 21081 14995 21147 14998
rect 21357 14995 21423 14998
rect 21633 15058 21699 15061
rect 26141 15058 26207 15061
rect 21633 15056 26207 15058
rect 21633 15000 21638 15056
rect 21694 15000 26146 15056
rect 26202 15000 26207 15056
rect 21633 14998 26207 15000
rect 21633 14995 21699 14998
rect 26141 14995 26207 14998
rect 0 14922 480 14952
rect 6310 14922 6316 14924
rect 0 14862 6316 14922
rect 0 14832 480 14862
rect 6310 14860 6316 14862
rect 6380 14860 6386 14924
rect 6494 14860 6500 14924
rect 6564 14922 6570 14924
rect 6862 14922 6868 14924
rect 6564 14862 6868 14922
rect 6564 14860 6570 14862
rect 6862 14860 6868 14862
rect 6932 14860 6938 14924
rect 8385 14922 8451 14925
rect 12709 14922 12775 14925
rect 16941 14922 17007 14925
rect 22318 14922 22324 14924
rect 8385 14920 12775 14922
rect 8385 14864 8390 14920
rect 8446 14864 12714 14920
rect 12770 14864 12775 14920
rect 8385 14862 12775 14864
rect 8385 14859 8451 14862
rect 12709 14859 12775 14862
rect 12942 14862 15578 14922
rect 4470 14724 4476 14788
rect 4540 14786 4546 14788
rect 5165 14786 5231 14789
rect 4540 14784 5231 14786
rect 4540 14728 5170 14784
rect 5226 14728 5231 14784
rect 4540 14726 5231 14728
rect 4540 14724 4546 14726
rect 5165 14723 5231 14726
rect 6177 14786 6243 14789
rect 6729 14786 6795 14789
rect 8845 14786 8911 14789
rect 6177 14784 6562 14786
rect 6177 14728 6182 14784
rect 6238 14728 6562 14784
rect 6177 14726 6562 14728
rect 6177 14723 6243 14726
rect 4337 14652 4403 14653
rect 4286 14588 4292 14652
rect 4356 14650 4403 14652
rect 4356 14648 4448 14650
rect 4398 14592 4448 14648
rect 4356 14590 4448 14592
rect 4356 14588 4403 14590
rect 5206 14588 5212 14652
rect 5276 14650 5282 14652
rect 6361 14650 6427 14653
rect 5276 14648 6427 14650
rect 5276 14592 6366 14648
rect 6422 14592 6427 14648
rect 5276 14590 6427 14592
rect 6502 14650 6562 14726
rect 6729 14784 8911 14786
rect 6729 14728 6734 14784
rect 6790 14728 8850 14784
rect 8906 14728 8911 14784
rect 6729 14726 8911 14728
rect 6729 14723 6795 14726
rect 8845 14723 8911 14726
rect 11053 14786 11119 14789
rect 12942 14786 13002 14862
rect 11053 14784 13002 14786
rect 11053 14728 11058 14784
rect 11114 14728 13002 14784
rect 11053 14726 13002 14728
rect 13169 14786 13235 14789
rect 15377 14786 15443 14789
rect 13169 14784 15443 14786
rect 13169 14728 13174 14784
rect 13230 14728 15382 14784
rect 15438 14728 15443 14784
rect 13169 14726 15443 14728
rect 15518 14786 15578 14862
rect 16941 14920 22324 14922
rect 16941 14864 16946 14920
rect 17002 14864 22324 14920
rect 16941 14862 22324 14864
rect 16941 14859 17007 14862
rect 22318 14860 22324 14862
rect 22388 14922 22394 14924
rect 22645 14922 22711 14925
rect 22388 14920 22711 14922
rect 22388 14864 22650 14920
rect 22706 14864 22711 14920
rect 22388 14862 22711 14864
rect 22388 14860 22394 14862
rect 22645 14859 22711 14862
rect 24853 14922 24919 14925
rect 27520 14922 28000 14952
rect 24853 14920 28000 14922
rect 24853 14864 24858 14920
rect 24914 14864 28000 14920
rect 24853 14862 28000 14864
rect 24853 14859 24919 14862
rect 27520 14832 28000 14862
rect 17493 14786 17559 14789
rect 17861 14786 17927 14789
rect 15518 14784 17927 14786
rect 15518 14728 17498 14784
rect 17554 14728 17866 14784
rect 17922 14728 17927 14784
rect 15518 14726 17927 14728
rect 11053 14723 11119 14726
rect 13169 14723 13235 14726
rect 15377 14723 15443 14726
rect 17493 14723 17559 14726
rect 17861 14723 17927 14726
rect 20989 14786 21055 14789
rect 24025 14786 24091 14789
rect 20989 14784 24091 14786
rect 20989 14728 20994 14784
rect 21050 14728 24030 14784
rect 24086 14728 24091 14784
rect 20989 14726 24091 14728
rect 20989 14723 21055 14726
rect 24025 14723 24091 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 10041 14650 10107 14653
rect 22134 14650 22140 14652
rect 6502 14648 10107 14650
rect 6502 14592 10046 14648
rect 10102 14592 10107 14648
rect 6502 14590 10107 14592
rect 5276 14588 5282 14590
rect 4337 14587 4403 14588
rect 6361 14587 6427 14590
rect 10041 14587 10107 14590
rect 20532 14590 22140 14650
rect 8569 14516 8635 14517
rect 8518 14514 8524 14516
rect 8442 14454 8524 14514
rect 8588 14514 8635 14516
rect 16614 14514 16620 14516
rect 8588 14512 16620 14514
rect 8630 14456 16620 14512
rect 8518 14452 8524 14454
rect 8588 14454 16620 14456
rect 8588 14452 8635 14454
rect 16614 14452 16620 14454
rect 16684 14452 16690 14516
rect 17033 14514 17099 14517
rect 19425 14514 19491 14517
rect 20532 14514 20592 14590
rect 22134 14588 22140 14590
rect 22204 14588 22210 14652
rect 23473 14650 23539 14653
rect 23606 14650 23612 14652
rect 23473 14648 23612 14650
rect 23473 14592 23478 14648
rect 23534 14592 23612 14648
rect 23473 14590 23612 14592
rect 23473 14587 23539 14590
rect 23606 14588 23612 14590
rect 23676 14588 23682 14652
rect 17033 14512 19491 14514
rect 17033 14456 17038 14512
rect 17094 14456 19430 14512
rect 19486 14456 19491 14512
rect 17033 14454 19491 14456
rect 8569 14451 8635 14452
rect 17033 14451 17099 14454
rect 19425 14451 19491 14454
rect 19980 14454 20592 14514
rect 20713 14514 20779 14517
rect 20713 14512 24962 14514
rect 20713 14456 20718 14512
rect 20774 14456 24962 14512
rect 20713 14454 24962 14456
rect 0 14378 480 14408
rect 19980 14381 20040 14454
rect 20713 14451 20779 14454
rect 6729 14378 6795 14381
rect 0 14376 6795 14378
rect 0 14320 6734 14376
rect 6790 14320 6795 14376
rect 0 14318 6795 14320
rect 0 14288 480 14318
rect 6729 14315 6795 14318
rect 9857 14378 9923 14381
rect 13445 14378 13511 14381
rect 9857 14376 13511 14378
rect 9857 14320 9862 14376
rect 9918 14320 13450 14376
rect 13506 14320 13511 14376
rect 9857 14318 13511 14320
rect 9857 14315 9923 14318
rect 13445 14315 13511 14318
rect 13997 14378 14063 14381
rect 16757 14378 16823 14381
rect 13997 14376 16823 14378
rect 13997 14320 14002 14376
rect 14058 14320 16762 14376
rect 16818 14320 16823 14376
rect 13997 14318 16823 14320
rect 13997 14315 14063 14318
rect 16757 14315 16823 14318
rect 16941 14378 17007 14381
rect 19977 14378 20043 14381
rect 16941 14376 20043 14378
rect 16941 14320 16946 14376
rect 17002 14320 19982 14376
rect 20038 14320 20043 14376
rect 16941 14318 20043 14320
rect 16941 14315 17007 14318
rect 19977 14315 20043 14318
rect 20294 14316 20300 14380
rect 20364 14378 20370 14380
rect 24902 14378 24962 14454
rect 27520 14378 28000 14408
rect 20364 14318 24778 14378
rect 24902 14318 28000 14378
rect 20364 14316 20370 14318
rect 7189 14242 7255 14245
rect 13077 14242 13143 14245
rect 13353 14242 13419 14245
rect 7189 14240 13419 14242
rect 7189 14184 7194 14240
rect 7250 14184 13082 14240
rect 13138 14184 13358 14240
rect 13414 14184 13419 14240
rect 7189 14182 13419 14184
rect 7189 14179 7255 14182
rect 13077 14179 13143 14182
rect 13353 14179 13419 14182
rect 18229 14242 18295 14245
rect 20713 14242 20779 14245
rect 18229 14240 20779 14242
rect 18229 14184 18234 14240
rect 18290 14184 20718 14240
rect 20774 14184 20779 14240
rect 18229 14182 20779 14184
rect 18229 14179 18295 14182
rect 20713 14179 20779 14182
rect 22134 14180 22140 14244
rect 22204 14242 22210 14244
rect 22829 14242 22895 14245
rect 22204 14240 22895 14242
rect 22204 14184 22834 14240
rect 22890 14184 22895 14240
rect 22204 14182 22895 14184
rect 24718 14242 24778 14318
rect 27520 14288 28000 14318
rect 25078 14242 25084 14244
rect 24718 14182 25084 14242
rect 22204 14180 22210 14182
rect 22829 14179 22895 14182
rect 25078 14180 25084 14182
rect 25148 14180 25154 14244
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 6637 14106 6703 14109
rect 9489 14106 9555 14109
rect 6637 14104 9555 14106
rect 6637 14048 6642 14104
rect 6698 14048 9494 14104
rect 9550 14048 9555 14104
rect 6637 14046 9555 14048
rect 6637 14043 6703 14046
rect 9489 14043 9555 14046
rect 10041 14106 10107 14109
rect 14641 14106 14707 14109
rect 10041 14104 14707 14106
rect 10041 14048 10046 14104
rect 10102 14048 14646 14104
rect 14702 14048 14707 14104
rect 10041 14046 14707 14048
rect 10041 14043 10107 14046
rect 14641 14043 14707 14046
rect 16849 14106 16915 14109
rect 20161 14106 20227 14109
rect 16849 14104 20227 14106
rect 16849 14048 16854 14104
rect 16910 14048 20166 14104
rect 20222 14048 20227 14104
rect 16849 14046 20227 14048
rect 16849 14043 16915 14046
rect 20161 14043 20227 14046
rect 20345 14106 20411 14109
rect 23013 14106 23079 14109
rect 20345 14104 23079 14106
rect 20345 14048 20350 14104
rect 20406 14048 23018 14104
rect 23074 14048 23079 14104
rect 20345 14046 23079 14048
rect 20345 14043 20411 14046
rect 23013 14043 23079 14046
rect 3785 13970 3851 13973
rect 9673 13970 9739 13973
rect 11053 13970 11119 13973
rect 3785 13968 7252 13970
rect 3785 13912 3790 13968
rect 3846 13912 7252 13968
rect 3785 13910 7252 13912
rect 3785 13907 3851 13910
rect 4153 13834 4219 13837
rect 6637 13834 6703 13837
rect 4153 13832 6703 13834
rect 4153 13776 4158 13832
rect 4214 13776 6642 13832
rect 6698 13776 6703 13832
rect 4153 13774 6703 13776
rect 4153 13771 4219 13774
rect 6637 13771 6703 13774
rect 0 13698 480 13728
rect 4245 13698 4311 13701
rect 7046 13698 7052 13700
rect 0 13696 4311 13698
rect 0 13640 4250 13696
rect 4306 13640 4311 13696
rect 0 13638 4311 13640
rect 0 13608 480 13638
rect 4245 13635 4311 13638
rect 4478 13638 7052 13698
rect 2773 13562 2839 13565
rect 4478 13562 4538 13638
rect 7046 13636 7052 13638
rect 7116 13636 7122 13700
rect 7192 13698 7252 13910
rect 9673 13968 11119 13970
rect 9673 13912 9678 13968
rect 9734 13912 11058 13968
rect 11114 13912 11119 13968
rect 9673 13910 11119 13912
rect 9673 13907 9739 13910
rect 11053 13907 11119 13910
rect 11697 13970 11763 13973
rect 16297 13970 16363 13973
rect 11697 13968 16363 13970
rect 11697 13912 11702 13968
rect 11758 13912 16302 13968
rect 16358 13912 16363 13968
rect 11697 13910 16363 13912
rect 11697 13907 11763 13910
rect 16297 13907 16363 13910
rect 16614 13908 16620 13972
rect 16684 13970 16690 13972
rect 20294 13970 20300 13972
rect 16684 13910 20300 13970
rect 16684 13908 16690 13910
rect 20294 13908 20300 13910
rect 20364 13908 20370 13972
rect 20846 13908 20852 13972
rect 20916 13970 20922 13972
rect 21357 13970 21423 13973
rect 20916 13968 21423 13970
rect 20916 13912 21362 13968
rect 21418 13912 21423 13968
rect 20916 13910 21423 13912
rect 20916 13908 20922 13910
rect 21357 13907 21423 13910
rect 24853 13970 24919 13973
rect 25405 13970 25471 13973
rect 24853 13968 25471 13970
rect 24853 13912 24858 13968
rect 24914 13912 25410 13968
rect 25466 13912 25471 13968
rect 24853 13910 25471 13912
rect 24853 13907 24919 13910
rect 25405 13907 25471 13910
rect 9765 13834 9831 13837
rect 14733 13834 14799 13837
rect 19701 13834 19767 13837
rect 9765 13832 14799 13834
rect 9765 13776 9770 13832
rect 9826 13776 14738 13832
rect 14794 13776 14799 13832
rect 9765 13774 14799 13776
rect 9765 13771 9831 13774
rect 14733 13771 14799 13774
rect 19382 13832 19767 13834
rect 19382 13776 19706 13832
rect 19762 13776 19767 13832
rect 19382 13774 19767 13776
rect 9673 13698 9739 13701
rect 7192 13696 9739 13698
rect 7192 13640 9678 13696
rect 9734 13640 9739 13696
rect 7192 13638 9739 13640
rect 9673 13635 9739 13638
rect 19057 13698 19123 13701
rect 19382 13698 19442 13774
rect 19701 13771 19767 13774
rect 20161 13834 20227 13837
rect 21173 13834 21239 13837
rect 20161 13832 21239 13834
rect 20161 13776 20166 13832
rect 20222 13776 21178 13832
rect 21234 13776 21239 13832
rect 20161 13774 21239 13776
rect 20161 13771 20227 13774
rect 21173 13771 21239 13774
rect 19057 13696 19442 13698
rect 19057 13640 19062 13696
rect 19118 13640 19442 13696
rect 19057 13638 19442 13640
rect 19057 13635 19123 13638
rect 20110 13636 20116 13700
rect 20180 13698 20186 13700
rect 20662 13698 20668 13700
rect 20180 13638 20668 13698
rect 20180 13636 20186 13638
rect 20662 13636 20668 13638
rect 20732 13636 20738 13700
rect 21030 13636 21036 13700
rect 21100 13698 21106 13700
rect 25221 13698 25287 13701
rect 27520 13698 28000 13728
rect 21100 13638 25146 13698
rect 21100 13636 21106 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 2773 13560 4538 13562
rect 2773 13504 2778 13560
rect 2834 13504 4538 13560
rect 2773 13502 4538 13504
rect 4613 13562 4679 13565
rect 4838 13562 4844 13564
rect 4613 13560 4844 13562
rect 4613 13504 4618 13560
rect 4674 13504 4844 13560
rect 4613 13502 4844 13504
rect 2773 13499 2839 13502
rect 4613 13499 4679 13502
rect 4838 13500 4844 13502
rect 4908 13500 4914 13564
rect 5390 13500 5396 13564
rect 5460 13562 5466 13564
rect 6085 13562 6151 13565
rect 5460 13560 6151 13562
rect 5460 13504 6090 13560
rect 6146 13504 6151 13560
rect 5460 13502 6151 13504
rect 5460 13500 5466 13502
rect 6085 13499 6151 13502
rect 6310 13500 6316 13564
rect 6380 13562 6386 13564
rect 10041 13562 10107 13565
rect 6380 13560 10107 13562
rect 6380 13504 10046 13560
rect 10102 13504 10107 13560
rect 6380 13502 10107 13504
rect 6380 13500 6386 13502
rect 10041 13499 10107 13502
rect 11053 13562 11119 13565
rect 16757 13562 16823 13565
rect 11053 13560 16823 13562
rect 11053 13504 11058 13560
rect 11114 13504 16762 13560
rect 16818 13504 16823 13560
rect 11053 13502 16823 13504
rect 11053 13499 11119 13502
rect 16757 13499 16823 13502
rect 19241 13562 19307 13565
rect 19374 13562 19380 13564
rect 19241 13560 19380 13562
rect 19241 13504 19246 13560
rect 19302 13504 19380 13560
rect 19241 13502 19380 13504
rect 19241 13499 19307 13502
rect 19374 13500 19380 13502
rect 19444 13500 19450 13564
rect 20069 13562 20135 13565
rect 22277 13562 22343 13565
rect 22553 13564 22619 13565
rect 22502 13562 22508 13564
rect 20069 13560 22343 13562
rect 20069 13504 20074 13560
rect 20130 13504 22282 13560
rect 22338 13504 22343 13560
rect 20069 13502 22343 13504
rect 22462 13502 22508 13562
rect 22572 13560 22619 13564
rect 22614 13504 22619 13560
rect 20069 13499 20135 13502
rect 22277 13499 22343 13502
rect 22502 13500 22508 13502
rect 22572 13500 22619 13504
rect 23422 13500 23428 13564
rect 23492 13562 23498 13564
rect 23933 13562 23999 13565
rect 23492 13560 23999 13562
rect 23492 13504 23938 13560
rect 23994 13504 23999 13560
rect 23492 13502 23999 13504
rect 23492 13500 23498 13502
rect 22553 13499 22619 13500
rect 23933 13499 23999 13502
rect 24117 13562 24183 13565
rect 24710 13562 24716 13564
rect 24117 13560 24716 13562
rect 24117 13504 24122 13560
rect 24178 13504 24716 13560
rect 24117 13502 24716 13504
rect 24117 13499 24183 13502
rect 24710 13500 24716 13502
rect 24780 13500 24786 13564
rect 3141 13426 3207 13429
rect 4797 13426 4863 13429
rect 3141 13424 4863 13426
rect 3141 13368 3146 13424
rect 3202 13368 4802 13424
rect 4858 13368 4863 13424
rect 3141 13366 4863 13368
rect 3141 13363 3207 13366
rect 4797 13363 4863 13366
rect 5441 13426 5507 13429
rect 7925 13426 7991 13429
rect 5441 13424 7991 13426
rect 5441 13368 5446 13424
rect 5502 13368 7930 13424
rect 7986 13368 7991 13424
rect 5441 13366 7991 13368
rect 5441 13363 5507 13366
rect 7925 13363 7991 13366
rect 13721 13426 13787 13429
rect 15929 13426 15995 13429
rect 22737 13426 22803 13429
rect 13721 13424 22803 13426
rect 13721 13368 13726 13424
rect 13782 13368 15934 13424
rect 15990 13368 22742 13424
rect 22798 13368 22803 13424
rect 13721 13366 22803 13368
rect 13721 13363 13787 13366
rect 15929 13363 15995 13366
rect 22737 13363 22803 13366
rect 23289 13426 23355 13429
rect 24025 13426 24091 13429
rect 23289 13424 24091 13426
rect 23289 13368 23294 13424
rect 23350 13368 24030 13424
rect 24086 13368 24091 13424
rect 23289 13366 24091 13368
rect 23289 13363 23355 13366
rect 24025 13363 24091 13366
rect 4337 13290 4403 13293
rect 10685 13290 10751 13293
rect 16481 13290 16547 13293
rect 24945 13290 25011 13293
rect 4337 13288 10751 13290
rect 4337 13232 4342 13288
rect 4398 13232 10690 13288
rect 10746 13232 10751 13288
rect 4337 13230 10751 13232
rect 4337 13227 4403 13230
rect 10685 13227 10751 13230
rect 13724 13230 15394 13290
rect 3918 13092 3924 13156
rect 3988 13154 3994 13156
rect 4061 13154 4127 13157
rect 5022 13154 5028 13156
rect 3988 13152 5028 13154
rect 3988 13096 4066 13152
rect 4122 13096 5028 13152
rect 3988 13094 5028 13096
rect 3988 13092 3994 13094
rect 4061 13091 4127 13094
rect 5022 13092 5028 13094
rect 5092 13092 5098 13156
rect 6678 13092 6684 13156
rect 6748 13154 6754 13156
rect 7598 13154 7604 13156
rect 6748 13094 7604 13154
rect 6748 13092 6754 13094
rect 7598 13092 7604 13094
rect 7668 13092 7674 13156
rect 7925 13154 7991 13157
rect 13724 13154 13784 13230
rect 7925 13152 13784 13154
rect 7925 13096 7930 13152
rect 7986 13096 13784 13152
rect 7925 13094 13784 13096
rect 13905 13154 13971 13157
rect 14038 13154 14044 13156
rect 13905 13152 14044 13154
rect 13905 13096 13910 13152
rect 13966 13096 14044 13152
rect 13905 13094 14044 13096
rect 7925 13091 7991 13094
rect 13905 13091 13971 13094
rect 14038 13092 14044 13094
rect 14108 13092 14114 13156
rect 5610 13088 5930 13089
rect 0 13018 480 13048
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 2865 13018 2931 13021
rect 0 13016 2931 13018
rect 0 12960 2870 13016
rect 2926 12960 2931 13016
rect 0 12958 2931 12960
rect 0 12928 480 12958
rect 2865 12955 2931 12958
rect 3233 13018 3299 13021
rect 5993 13018 6059 13021
rect 7046 13018 7052 13020
rect 3233 13016 5458 13018
rect 3233 12960 3238 13016
rect 3294 12960 5458 13016
rect 3233 12958 5458 12960
rect 3233 12955 3299 12958
rect 1393 12882 1459 12885
rect 5257 12882 5323 12885
rect 1393 12880 5323 12882
rect 1393 12824 1398 12880
rect 1454 12824 5262 12880
rect 5318 12824 5323 12880
rect 1393 12822 5323 12824
rect 5398 12882 5458 12958
rect 5993 13016 7052 13018
rect 5993 12960 5998 13016
rect 6054 12960 7052 13016
rect 5993 12958 7052 12960
rect 5993 12955 6059 12958
rect 7046 12956 7052 12958
rect 7116 12956 7122 13020
rect 7966 12956 7972 13020
rect 8036 13018 8042 13020
rect 9029 13018 9095 13021
rect 8036 13016 9095 13018
rect 8036 12960 9034 13016
rect 9090 12960 9095 13016
rect 8036 12958 9095 12960
rect 8036 12956 8042 12958
rect 9029 12955 9095 12958
rect 9673 13018 9739 13021
rect 15334 13018 15394 13230
rect 16481 13288 25011 13290
rect 16481 13232 16486 13288
rect 16542 13232 24950 13288
rect 25006 13232 25011 13288
rect 16481 13230 25011 13232
rect 16481 13227 16547 13230
rect 24945 13227 25011 13230
rect 16757 13154 16823 13157
rect 24117 13154 24183 13157
rect 16757 13152 24183 13154
rect 16757 13096 16762 13152
rect 16818 13096 24122 13152
rect 24178 13096 24183 13152
rect 16757 13094 24183 13096
rect 25086 13154 25146 13638
rect 25221 13696 28000 13698
rect 25221 13640 25226 13696
rect 25282 13640 28000 13696
rect 25221 13638 28000 13640
rect 25221 13635 25287 13638
rect 27520 13608 28000 13638
rect 25957 13564 26023 13565
rect 25957 13560 26004 13564
rect 26068 13562 26074 13564
rect 25957 13504 25962 13560
rect 25957 13500 26004 13504
rect 26068 13502 26114 13562
rect 26068 13500 26074 13502
rect 25957 13499 26023 13500
rect 27520 13154 28000 13184
rect 25086 13094 28000 13154
rect 16757 13091 16823 13094
rect 24117 13091 24183 13094
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 9673 13016 14658 13018
rect 9673 12960 9678 13016
rect 9734 12960 14658 13016
rect 9673 12958 14658 12960
rect 15334 12958 24042 13018
rect 9673 12955 9739 12958
rect 14365 12882 14431 12885
rect 5398 12880 14431 12882
rect 5398 12824 14370 12880
rect 14426 12824 14431 12880
rect 5398 12822 14431 12824
rect 1393 12819 1459 12822
rect 5257 12819 5323 12822
rect 14365 12819 14431 12822
rect 1393 12746 1459 12749
rect 10593 12746 10659 12749
rect 1393 12744 10659 12746
rect 1393 12688 1398 12744
rect 1454 12688 10598 12744
rect 10654 12688 10659 12744
rect 1393 12686 10659 12688
rect 14598 12746 14658 12958
rect 14733 12882 14799 12885
rect 19149 12882 19215 12885
rect 14733 12880 19215 12882
rect 14733 12824 14738 12880
rect 14794 12824 19154 12880
rect 19210 12824 19215 12880
rect 14733 12822 19215 12824
rect 14733 12819 14799 12822
rect 19149 12819 19215 12822
rect 19333 12884 19399 12885
rect 19333 12880 19380 12884
rect 19444 12882 19450 12884
rect 19793 12882 19859 12885
rect 23473 12882 23539 12885
rect 19333 12824 19338 12880
rect 19333 12820 19380 12824
rect 19444 12822 19490 12882
rect 19793 12880 23539 12882
rect 19793 12824 19798 12880
rect 19854 12824 23478 12880
rect 23534 12824 23539 12880
rect 19793 12822 23539 12824
rect 23982 12882 24042 12958
rect 25221 12882 25287 12885
rect 23982 12880 25287 12882
rect 23982 12824 25226 12880
rect 25282 12824 25287 12880
rect 23982 12822 25287 12824
rect 19444 12820 19450 12822
rect 19333 12819 19399 12820
rect 19793 12819 19859 12822
rect 23473 12819 23539 12822
rect 25221 12819 25287 12822
rect 18873 12746 18939 12749
rect 22461 12746 22527 12749
rect 24025 12746 24091 12749
rect 14598 12744 22018 12746
rect 14598 12688 18878 12744
rect 18934 12688 22018 12744
rect 14598 12686 22018 12688
rect 1393 12683 1459 12686
rect 10593 12683 10659 12686
rect 18873 12683 18939 12686
rect 2865 12610 2931 12613
rect 3325 12612 3391 12613
rect 3325 12610 3372 12612
rect 2865 12608 3112 12610
rect 2865 12552 2870 12608
rect 2926 12552 3112 12608
rect 2865 12550 3112 12552
rect 3244 12608 3372 12610
rect 3436 12610 3442 12612
rect 3877 12610 3943 12613
rect 3436 12608 3943 12610
rect 3244 12552 3330 12608
rect 3436 12552 3882 12608
rect 3938 12552 3943 12608
rect 3244 12550 3372 12552
rect 2865 12547 2931 12550
rect 3052 12474 3112 12550
rect 3325 12548 3372 12550
rect 3436 12550 3943 12552
rect 3436 12548 3442 12550
rect 3325 12547 3391 12548
rect 3877 12547 3943 12550
rect 4429 12610 4495 12613
rect 4797 12610 4863 12613
rect 4429 12608 4863 12610
rect 4429 12552 4434 12608
rect 4490 12552 4802 12608
rect 4858 12552 4863 12608
rect 4429 12550 4863 12552
rect 4429 12547 4495 12550
rect 4797 12547 4863 12550
rect 11094 12548 11100 12612
rect 11164 12610 11170 12612
rect 11237 12610 11303 12613
rect 15101 12610 15167 12613
rect 11164 12608 15167 12610
rect 11164 12552 11242 12608
rect 11298 12552 15106 12608
rect 15162 12552 15167 12608
rect 11164 12550 15167 12552
rect 11164 12548 11170 12550
rect 11237 12547 11303 12550
rect 15101 12547 15167 12550
rect 20529 12610 20595 12613
rect 21633 12610 21699 12613
rect 21958 12610 22018 12686
rect 22461 12744 24091 12746
rect 22461 12688 22466 12744
rect 22522 12688 24030 12744
rect 24086 12688 24091 12744
rect 22461 12686 24091 12688
rect 22461 12683 22527 12686
rect 24025 12683 24091 12686
rect 22461 12610 22527 12613
rect 20529 12608 21834 12610
rect 20529 12552 20534 12608
rect 20590 12552 21638 12608
rect 21694 12552 21834 12608
rect 20529 12550 21834 12552
rect 21958 12608 22527 12610
rect 21958 12552 22466 12608
rect 22522 12552 22527 12608
rect 21958 12550 22527 12552
rect 20529 12547 20595 12550
rect 21633 12547 21699 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 7966 12474 7972 12476
rect 3052 12414 7972 12474
rect 7966 12412 7972 12414
rect 8036 12412 8042 12476
rect 8109 12474 8175 12477
rect 8886 12474 8892 12476
rect 8109 12472 8892 12474
rect 8109 12416 8114 12472
rect 8170 12416 8892 12472
rect 8109 12414 8892 12416
rect 8109 12411 8175 12414
rect 8886 12412 8892 12414
rect 8956 12412 8962 12476
rect 9673 12474 9739 12477
rect 9857 12474 9923 12477
rect 9673 12472 9923 12474
rect 9673 12416 9678 12472
rect 9734 12416 9862 12472
rect 9918 12416 9923 12472
rect 9673 12414 9923 12416
rect 9673 12411 9739 12414
rect 9857 12411 9923 12414
rect 14590 12412 14596 12476
rect 14660 12474 14666 12476
rect 19333 12474 19399 12477
rect 14660 12472 19399 12474
rect 14660 12416 19338 12472
rect 19394 12416 19399 12472
rect 14660 12414 19399 12416
rect 21774 12474 21834 12550
rect 22461 12547 22527 12550
rect 23422 12548 23428 12612
rect 23492 12610 23498 12612
rect 27520 12610 28000 12640
rect 23492 12550 28000 12610
rect 23492 12548 23498 12550
rect 27520 12520 28000 12550
rect 25037 12474 25103 12477
rect 21774 12472 25103 12474
rect 21774 12416 25042 12472
rect 25098 12416 25103 12472
rect 21774 12414 25103 12416
rect 14660 12412 14666 12414
rect 19333 12411 19399 12414
rect 25037 12411 25103 12414
rect 0 12338 480 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 480 12278
rect 1485 12275 1551 12278
rect 2497 12338 2563 12341
rect 3550 12338 3556 12340
rect 2497 12336 3556 12338
rect 2497 12280 2502 12336
rect 2558 12280 3556 12336
rect 2497 12278 3556 12280
rect 2497 12275 2563 12278
rect 3550 12276 3556 12278
rect 3620 12276 3626 12340
rect 4061 12338 4127 12341
rect 8150 12338 8156 12340
rect 4061 12336 8156 12338
rect 4061 12280 4066 12336
rect 4122 12280 8156 12336
rect 4061 12278 8156 12280
rect 4061 12275 4127 12278
rect 8150 12276 8156 12278
rect 8220 12276 8226 12340
rect 9029 12338 9095 12341
rect 9438 12338 9444 12340
rect 9029 12336 9444 12338
rect 9029 12280 9034 12336
rect 9090 12280 9444 12336
rect 9029 12278 9444 12280
rect 9029 12275 9095 12278
rect 9438 12276 9444 12278
rect 9508 12276 9514 12340
rect 9673 12338 9739 12341
rect 12382 12338 12388 12340
rect 9673 12336 12388 12338
rect 9673 12280 9678 12336
rect 9734 12280 12388 12336
rect 9673 12278 12388 12280
rect 9673 12275 9739 12278
rect 12382 12276 12388 12278
rect 12452 12276 12458 12340
rect 12525 12338 12591 12341
rect 20253 12338 20319 12341
rect 12525 12336 20319 12338
rect 12525 12280 12530 12336
rect 12586 12280 20258 12336
rect 20314 12280 20319 12336
rect 12525 12278 20319 12280
rect 12525 12275 12591 12278
rect 20253 12275 20319 12278
rect 21030 12276 21036 12340
rect 21100 12338 21106 12340
rect 21100 12278 24732 12338
rect 21100 12276 21106 12278
rect 2957 12202 3023 12205
rect 8201 12202 8267 12205
rect 8753 12202 8819 12205
rect 14917 12202 14983 12205
rect 2957 12200 7666 12202
rect 2957 12144 2962 12200
rect 3018 12144 7666 12200
rect 2957 12142 7666 12144
rect 2957 12139 3023 12142
rect 7606 12066 7666 12142
rect 8201 12200 14983 12202
rect 8201 12144 8206 12200
rect 8262 12144 8758 12200
rect 8814 12144 14922 12200
rect 14978 12144 14983 12200
rect 8201 12142 14983 12144
rect 8201 12139 8267 12142
rect 8753 12139 8819 12142
rect 14917 12139 14983 12142
rect 15101 12202 15167 12205
rect 15653 12202 15719 12205
rect 18965 12202 19031 12205
rect 15101 12200 15394 12202
rect 15101 12144 15106 12200
rect 15162 12144 15394 12200
rect 15101 12142 15394 12144
rect 15101 12139 15167 12142
rect 12525 12066 12591 12069
rect 7606 12064 12591 12066
rect 7606 12008 12530 12064
rect 12586 12008 12591 12064
rect 7606 12006 12591 12008
rect 15334 12066 15394 12142
rect 15653 12200 19031 12202
rect 15653 12144 15658 12200
rect 15714 12144 18970 12200
rect 19026 12144 19031 12200
rect 15653 12142 19031 12144
rect 15653 12139 15719 12142
rect 18965 12139 19031 12142
rect 19149 12202 19215 12205
rect 24301 12202 24367 12205
rect 19149 12200 24367 12202
rect 19149 12144 19154 12200
rect 19210 12144 24306 12200
rect 24362 12144 24367 12200
rect 19149 12142 24367 12144
rect 19149 12139 19215 12142
rect 24301 12139 24367 12142
rect 23841 12066 23907 12069
rect 15334 12064 23907 12066
rect 15334 12008 23846 12064
rect 23902 12008 23907 12064
rect 15334 12006 23907 12008
rect 24672 12066 24732 12278
rect 27520 12066 28000 12096
rect 24672 12006 28000 12066
rect 12525 12003 12591 12006
rect 23841 12003 23907 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 27520 11976 28000 12006
rect 24277 11935 24597 11936
rect 3141 11930 3207 11933
rect 4797 11930 4863 11933
rect 5022 11930 5028 11932
rect 3141 11928 5028 11930
rect 3141 11872 3146 11928
rect 3202 11872 4802 11928
rect 4858 11872 5028 11928
rect 3141 11870 5028 11872
rect 3141 11867 3207 11870
rect 4797 11867 4863 11870
rect 5022 11868 5028 11870
rect 5092 11868 5098 11932
rect 6126 11868 6132 11932
rect 6196 11930 6202 11932
rect 6494 11930 6500 11932
rect 6196 11870 6500 11930
rect 6196 11868 6202 11870
rect 6494 11868 6500 11870
rect 6564 11868 6570 11932
rect 8477 11930 8543 11933
rect 18597 11930 18663 11933
rect 20253 11930 20319 11933
rect 21265 11932 21331 11933
rect 8477 11928 14060 11930
rect 8477 11872 8482 11928
rect 8538 11872 14060 11928
rect 8477 11870 14060 11872
rect 8477 11867 8543 11870
rect 3509 11794 3575 11797
rect 4654 11794 4660 11796
rect 3509 11792 4660 11794
rect 3509 11736 3514 11792
rect 3570 11736 4660 11792
rect 3509 11734 4660 11736
rect 3509 11731 3575 11734
rect 4654 11732 4660 11734
rect 4724 11732 4730 11796
rect 6126 11732 6132 11796
rect 6196 11794 6202 11796
rect 6637 11794 6703 11797
rect 6196 11792 6703 11794
rect 6196 11736 6642 11792
rect 6698 11736 6703 11792
rect 6196 11734 6703 11736
rect 6196 11732 6202 11734
rect 6637 11731 6703 11734
rect 8109 11794 8175 11797
rect 10685 11794 10751 11797
rect 8109 11792 10751 11794
rect 8109 11736 8114 11792
rect 8170 11736 10690 11792
rect 10746 11736 10751 11792
rect 8109 11734 10751 11736
rect 14000 11794 14060 11870
rect 18597 11928 20319 11930
rect 18597 11872 18602 11928
rect 18658 11872 20258 11928
rect 20314 11872 20319 11928
rect 18597 11870 20319 11872
rect 18597 11867 18663 11870
rect 20253 11867 20319 11870
rect 21214 11868 21220 11932
rect 21284 11930 21331 11932
rect 24853 11932 24919 11933
rect 24853 11930 24900 11932
rect 21284 11928 21376 11930
rect 21326 11872 21376 11928
rect 21284 11870 21376 11872
rect 24808 11928 24900 11930
rect 24808 11872 24858 11928
rect 24808 11870 24900 11872
rect 21284 11868 21331 11870
rect 21265 11867 21331 11868
rect 24853 11868 24900 11870
rect 24964 11868 24970 11932
rect 24853 11867 24919 11868
rect 18321 11794 18387 11797
rect 14000 11792 18387 11794
rect 14000 11736 18326 11792
rect 18382 11736 18387 11792
rect 14000 11734 18387 11736
rect 8109 11731 8175 11734
rect 10685 11731 10751 11734
rect 18321 11731 18387 11734
rect 18505 11794 18571 11797
rect 21030 11794 21036 11796
rect 18505 11792 21036 11794
rect 18505 11736 18510 11792
rect 18566 11736 21036 11792
rect 18505 11734 21036 11736
rect 18505 11731 18571 11734
rect 21030 11732 21036 11734
rect 21100 11732 21106 11796
rect 22553 11794 22619 11797
rect 25037 11794 25103 11797
rect 22553 11792 25103 11794
rect 22553 11736 22558 11792
rect 22614 11736 25042 11792
rect 25098 11736 25103 11792
rect 22553 11734 25103 11736
rect 22553 11731 22619 11734
rect 25037 11731 25103 11734
rect 0 11658 480 11688
rect 4613 11658 4679 11661
rect 0 11656 4679 11658
rect 0 11600 4618 11656
rect 4674 11600 4679 11656
rect 0 11598 4679 11600
rect 0 11568 480 11598
rect 4613 11595 4679 11598
rect 5165 11658 5231 11661
rect 7833 11658 7899 11661
rect 5165 11656 7899 11658
rect 5165 11600 5170 11656
rect 5226 11600 7838 11656
rect 7894 11600 7899 11656
rect 5165 11598 7899 11600
rect 5165 11595 5231 11598
rect 7833 11595 7899 11598
rect 8937 11658 9003 11661
rect 12341 11658 12407 11661
rect 8937 11656 12407 11658
rect 8937 11600 8942 11656
rect 8998 11600 12346 11656
rect 12402 11600 12407 11656
rect 8937 11598 12407 11600
rect 8937 11595 9003 11598
rect 12341 11595 12407 11598
rect 14181 11658 14247 11661
rect 15653 11658 15719 11661
rect 14181 11656 15719 11658
rect 14181 11600 14186 11656
rect 14242 11600 15658 11656
rect 15714 11600 15719 11656
rect 14181 11598 15719 11600
rect 14181 11595 14247 11598
rect 15653 11595 15719 11598
rect 16389 11658 16455 11661
rect 18873 11658 18939 11661
rect 25589 11658 25655 11661
rect 16389 11656 25655 11658
rect 16389 11600 16394 11656
rect 16450 11600 18878 11656
rect 18934 11600 25594 11656
rect 25650 11600 25655 11656
rect 16389 11598 25655 11600
rect 16389 11595 16455 11598
rect 18873 11595 18939 11598
rect 25589 11595 25655 11598
rect 4705 11522 4771 11525
rect 8293 11522 8359 11525
rect 8845 11524 8911 11525
rect 10777 11524 10843 11525
rect 8845 11522 8892 11524
rect 4705 11520 8359 11522
rect 4705 11464 4710 11520
rect 4766 11464 8298 11520
rect 8354 11464 8359 11520
rect 4705 11462 8359 11464
rect 8800 11520 8892 11522
rect 8800 11464 8850 11520
rect 8800 11462 8892 11464
rect 4705 11459 4771 11462
rect 8293 11459 8359 11462
rect 8845 11460 8892 11462
rect 8956 11460 8962 11524
rect 10726 11460 10732 11524
rect 10796 11522 10843 11524
rect 14825 11522 14891 11525
rect 19333 11522 19399 11525
rect 23473 11522 23539 11525
rect 27520 11522 28000 11552
rect 10796 11520 10888 11522
rect 10838 11464 10888 11520
rect 10796 11462 10888 11464
rect 14825 11520 19399 11522
rect 14825 11464 14830 11520
rect 14886 11464 19338 11520
rect 19394 11464 19399 11520
rect 14825 11462 19399 11464
rect 10796 11460 10843 11462
rect 8845 11459 8911 11460
rect 10777 11459 10843 11460
rect 14825 11459 14891 11462
rect 19333 11459 19399 11462
rect 20118 11462 23306 11522
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 1393 11386 1459 11389
rect 5901 11386 5967 11389
rect 1393 11384 5967 11386
rect 1393 11328 1398 11384
rect 1454 11328 5906 11384
rect 5962 11328 5967 11384
rect 1393 11326 5967 11328
rect 1393 11323 1459 11326
rect 5901 11323 5967 11326
rect 6637 11386 6703 11389
rect 9765 11386 9831 11389
rect 6637 11384 9831 11386
rect 6637 11328 6642 11384
rect 6698 11328 9770 11384
rect 9826 11328 9831 11384
rect 6637 11326 9831 11328
rect 6637 11323 6703 11326
rect 9765 11323 9831 11326
rect 12382 11324 12388 11388
rect 12452 11386 12458 11388
rect 12452 11326 18522 11386
rect 12452 11324 12458 11326
rect 2129 11250 2195 11253
rect 2957 11250 3023 11253
rect 17769 11250 17835 11253
rect 2129 11248 17835 11250
rect 2129 11192 2134 11248
rect 2190 11192 2962 11248
rect 3018 11192 17774 11248
rect 17830 11192 17835 11248
rect 2129 11190 17835 11192
rect 2129 11187 2195 11190
rect 2957 11187 3023 11190
rect 17769 11187 17835 11190
rect 1577 11114 1643 11117
rect 8017 11114 8083 11117
rect 10317 11114 10383 11117
rect 15469 11114 15535 11117
rect 1577 11112 6700 11114
rect 1577 11056 1582 11112
rect 1638 11056 6700 11112
rect 1577 11054 6700 11056
rect 1577 11051 1643 11054
rect 0 10978 480 11008
rect 6640 10981 6700 11054
rect 8017 11112 15535 11114
rect 8017 11056 8022 11112
rect 8078 11056 10322 11112
rect 10378 11056 15474 11112
rect 15530 11056 15535 11112
rect 8017 11054 15535 11056
rect 18462 11114 18522 11326
rect 18965 11250 19031 11253
rect 20118 11250 20178 11462
rect 20294 11324 20300 11388
rect 20364 11386 20370 11388
rect 22829 11386 22895 11389
rect 20364 11384 22895 11386
rect 20364 11328 22834 11384
rect 22890 11328 22895 11384
rect 20364 11326 22895 11328
rect 20364 11324 20370 11326
rect 22829 11323 22895 11326
rect 18965 11248 20178 11250
rect 18965 11192 18970 11248
rect 19026 11192 20178 11248
rect 18965 11190 20178 11192
rect 20253 11250 20319 11253
rect 23013 11250 23079 11253
rect 20253 11248 23079 11250
rect 20253 11192 20258 11248
rect 20314 11192 23018 11248
rect 23074 11192 23079 11248
rect 20253 11190 23079 11192
rect 23246 11250 23306 11462
rect 23473 11520 28000 11522
rect 23473 11464 23478 11520
rect 23534 11464 28000 11520
rect 23473 11462 28000 11464
rect 23473 11459 23539 11462
rect 27520 11432 28000 11462
rect 24209 11386 24275 11389
rect 24894 11386 24900 11388
rect 24209 11384 24900 11386
rect 24209 11328 24214 11384
rect 24270 11328 24900 11384
rect 24209 11326 24900 11328
rect 24209 11323 24275 11326
rect 24894 11324 24900 11326
rect 24964 11324 24970 11388
rect 25957 11250 26023 11253
rect 23246 11248 26023 11250
rect 23246 11192 25962 11248
rect 26018 11192 26023 11248
rect 23246 11190 26023 11192
rect 18965 11187 19031 11190
rect 20253 11187 20319 11190
rect 23013 11187 23079 11190
rect 25957 11187 26023 11190
rect 20069 11114 20135 11117
rect 18462 11112 20135 11114
rect 18462 11056 20074 11112
rect 20130 11056 20135 11112
rect 18462 11054 20135 11056
rect 8017 11051 8083 11054
rect 10317 11051 10383 11054
rect 15469 11051 15535 11054
rect 20069 11051 20135 11054
rect 3049 10978 3115 10981
rect 5257 10978 5323 10981
rect 0 10918 2146 10978
rect 0 10888 480 10918
rect 2086 10842 2146 10918
rect 3049 10976 5323 10978
rect 3049 10920 3054 10976
rect 3110 10920 5262 10976
rect 5318 10920 5323 10976
rect 3049 10918 5323 10920
rect 3049 10915 3115 10918
rect 5257 10915 5323 10918
rect 6637 10978 6703 10981
rect 15469 10980 15535 10981
rect 7046 10978 7052 10980
rect 6637 10976 7052 10978
rect 6637 10920 6642 10976
rect 6698 10920 7052 10976
rect 6637 10918 7052 10920
rect 6637 10915 6703 10918
rect 7046 10916 7052 10918
rect 7116 10916 7122 10980
rect 15469 10976 15516 10980
rect 15580 10978 15586 10980
rect 25589 10978 25655 10981
rect 27520 10978 28000 11008
rect 15469 10920 15474 10976
rect 15469 10916 15516 10920
rect 15580 10918 15626 10978
rect 25589 10976 28000 10978
rect 25589 10920 25594 10976
rect 25650 10920 28000 10976
rect 25589 10918 28000 10920
rect 15580 10916 15586 10918
rect 15469 10915 15535 10916
rect 25589 10915 25655 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 27520 10888 28000 10918
rect 24277 10847 24597 10848
rect 4981 10842 5047 10845
rect 2086 10840 5047 10842
rect 2086 10784 4986 10840
rect 5042 10784 5047 10840
rect 2086 10782 5047 10784
rect 4981 10779 5047 10782
rect 6269 10842 6335 10845
rect 14641 10844 14707 10845
rect 8518 10842 8524 10844
rect 6269 10840 8524 10842
rect 6269 10784 6274 10840
rect 6330 10784 8524 10840
rect 6269 10782 8524 10784
rect 6269 10779 6335 10782
rect 8518 10780 8524 10782
rect 8588 10780 8594 10844
rect 14590 10780 14596 10844
rect 14660 10842 14707 10844
rect 14660 10840 14752 10842
rect 14702 10784 14752 10840
rect 14660 10782 14752 10784
rect 14660 10780 14707 10782
rect 22318 10780 22324 10844
rect 22388 10842 22394 10844
rect 23565 10842 23631 10845
rect 22388 10840 23631 10842
rect 22388 10784 23570 10840
rect 23626 10784 23631 10840
rect 22388 10782 23631 10784
rect 22388 10780 22394 10782
rect 14641 10779 14707 10780
rect 23565 10779 23631 10782
rect 23974 10780 23980 10844
rect 24044 10842 24050 10844
rect 24117 10842 24183 10845
rect 24044 10840 24183 10842
rect 24044 10784 24122 10840
rect 24178 10784 24183 10840
rect 24044 10782 24183 10784
rect 24044 10780 24050 10782
rect 24117 10779 24183 10782
rect 2630 10644 2636 10708
rect 2700 10706 2706 10708
rect 3233 10706 3299 10709
rect 2700 10704 3299 10706
rect 2700 10648 3238 10704
rect 3294 10648 3299 10704
rect 2700 10646 3299 10648
rect 2700 10644 2706 10646
rect 3233 10643 3299 10646
rect 5165 10706 5231 10709
rect 17125 10706 17191 10709
rect 19333 10706 19399 10709
rect 5165 10704 17191 10706
rect 5165 10648 5170 10704
rect 5226 10648 17130 10704
rect 17186 10648 17191 10704
rect 5165 10646 17191 10648
rect 5165 10643 5231 10646
rect 17125 10643 17191 10646
rect 17910 10704 19399 10706
rect 17910 10648 19338 10704
rect 19394 10648 19399 10704
rect 17910 10646 19399 10648
rect 5257 10570 5323 10573
rect 7005 10570 7071 10573
rect 17769 10570 17835 10573
rect 5257 10568 17835 10570
rect 5257 10512 5262 10568
rect 5318 10512 7010 10568
rect 7066 10512 17774 10568
rect 17830 10512 17835 10568
rect 5257 10510 17835 10512
rect 5257 10507 5323 10510
rect 7005 10507 7071 10510
rect 17769 10507 17835 10510
rect 4889 10434 4955 10437
rect 9765 10434 9831 10437
rect 11329 10436 11395 10437
rect 11278 10434 11284 10436
rect 4889 10432 9831 10434
rect 4889 10376 4894 10432
rect 4950 10376 9770 10432
rect 9826 10376 9831 10432
rect 4889 10374 9831 10376
rect 11202 10374 11284 10434
rect 11348 10434 11395 10436
rect 17910 10434 17970 10646
rect 19333 10643 19399 10646
rect 20110 10644 20116 10708
rect 20180 10706 20186 10708
rect 20478 10706 20484 10708
rect 20180 10646 20484 10706
rect 20180 10644 20186 10646
rect 20478 10644 20484 10646
rect 20548 10644 20554 10708
rect 18597 10570 18663 10573
rect 25221 10570 25287 10573
rect 18597 10568 25287 10570
rect 18597 10512 18602 10568
rect 18658 10512 25226 10568
rect 25282 10512 25287 10568
rect 18597 10510 25287 10512
rect 18597 10507 18663 10510
rect 25221 10507 25287 10510
rect 11348 10432 17970 10434
rect 11390 10376 17970 10432
rect 4889 10371 4955 10374
rect 9765 10371 9831 10374
rect 11278 10372 11284 10374
rect 11348 10374 17970 10376
rect 21449 10434 21515 10437
rect 23933 10434 23999 10437
rect 21449 10432 23999 10434
rect 21449 10376 21454 10432
rect 21510 10376 23938 10432
rect 23994 10376 23999 10432
rect 21449 10374 23999 10376
rect 11348 10372 11395 10374
rect 11329 10371 11395 10372
rect 21449 10371 21515 10374
rect 23933 10371 23999 10374
rect 24117 10434 24183 10437
rect 24945 10434 25011 10437
rect 24117 10432 25011 10434
rect 24117 10376 24122 10432
rect 24178 10376 24950 10432
rect 25006 10376 25011 10432
rect 24117 10374 25011 10376
rect 24117 10371 24183 10374
rect 24945 10371 25011 10374
rect 26417 10434 26483 10437
rect 27520 10434 28000 10464
rect 26417 10432 28000 10434
rect 26417 10376 26422 10432
rect 26478 10376 28000 10432
rect 26417 10374 28000 10376
rect 26417 10371 26483 10374
rect 10277 10368 10597 10369
rect 0 10298 480 10328
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 27520 10344 28000 10374
rect 19610 10303 19930 10304
rect 3049 10298 3115 10301
rect 0 10296 3115 10298
rect 0 10240 3054 10296
rect 3110 10240 3115 10296
rect 0 10238 3115 10240
rect 0 10208 480 10238
rect 3049 10235 3115 10238
rect 5390 10236 5396 10300
rect 5460 10298 5466 10300
rect 5533 10298 5599 10301
rect 5460 10296 5599 10298
rect 5460 10240 5538 10296
rect 5594 10240 5599 10296
rect 5460 10238 5599 10240
rect 5460 10236 5466 10238
rect 5533 10235 5599 10238
rect 7097 10298 7163 10301
rect 7097 10296 8540 10298
rect 7097 10240 7102 10296
rect 7158 10240 8540 10296
rect 7097 10238 8540 10240
rect 7097 10235 7163 10238
rect 2865 10162 2931 10165
rect 8293 10162 8359 10165
rect 2865 10160 8359 10162
rect 2865 10104 2870 10160
rect 2926 10104 8298 10160
rect 8354 10104 8359 10160
rect 2865 10102 8359 10104
rect 8480 10162 8540 10238
rect 9990 10236 9996 10300
rect 10060 10298 10066 10300
rect 10133 10298 10199 10301
rect 10060 10296 10199 10298
rect 10060 10240 10138 10296
rect 10194 10240 10199 10296
rect 10060 10238 10199 10240
rect 10060 10236 10066 10238
rect 10133 10235 10199 10238
rect 12065 10298 12131 10301
rect 16389 10298 16455 10301
rect 22093 10300 22159 10301
rect 22369 10300 22435 10301
rect 22093 10298 22140 10300
rect 12065 10296 16455 10298
rect 12065 10240 12070 10296
rect 12126 10240 16394 10296
rect 16450 10240 16455 10296
rect 12065 10238 16455 10240
rect 22048 10296 22140 10298
rect 22048 10240 22098 10296
rect 22048 10238 22140 10240
rect 12065 10235 12131 10238
rect 16389 10235 16455 10238
rect 22093 10236 22140 10238
rect 22204 10236 22210 10300
rect 22318 10298 22324 10300
rect 22278 10238 22324 10298
rect 22388 10296 22435 10300
rect 22430 10240 22435 10296
rect 22318 10236 22324 10238
rect 22388 10236 22435 10240
rect 22093 10235 22159 10236
rect 22369 10235 22435 10236
rect 22737 10298 22803 10301
rect 25405 10298 25471 10301
rect 22737 10296 25471 10298
rect 22737 10240 22742 10296
rect 22798 10240 25410 10296
rect 25466 10240 25471 10296
rect 22737 10238 25471 10240
rect 22737 10235 22803 10238
rect 25405 10235 25471 10238
rect 17953 10162 18019 10165
rect 8480 10160 18019 10162
rect 8480 10104 17958 10160
rect 18014 10104 18019 10160
rect 8480 10102 18019 10104
rect 2865 10099 2931 10102
rect 8293 10099 8359 10102
rect 17953 10099 18019 10102
rect 19057 10162 19123 10165
rect 23473 10162 23539 10165
rect 19057 10160 23539 10162
rect 19057 10104 19062 10160
rect 19118 10104 23478 10160
rect 23534 10104 23539 10160
rect 19057 10102 23539 10104
rect 19057 10099 19123 10102
rect 23473 10099 23539 10102
rect 23657 10162 23723 10165
rect 24853 10162 24919 10165
rect 23657 10160 24919 10162
rect 23657 10104 23662 10160
rect 23718 10104 24858 10160
rect 24914 10104 24919 10160
rect 23657 10102 24919 10104
rect 23657 10099 23723 10102
rect 24853 10099 24919 10102
rect 2405 10026 2471 10029
rect 5717 10026 5783 10029
rect 2405 10024 5783 10026
rect 2405 9968 2410 10024
rect 2466 9968 5722 10024
rect 5778 9968 5783 10024
rect 2405 9966 5783 9968
rect 2405 9963 2471 9966
rect 5717 9963 5783 9966
rect 9397 10026 9463 10029
rect 20253 10026 20319 10029
rect 9397 10024 20319 10026
rect 9397 9968 9402 10024
rect 9458 9968 20258 10024
rect 20314 9968 20319 10024
rect 9397 9966 20319 9968
rect 9397 9963 9463 9966
rect 20253 9963 20319 9966
rect 22461 10026 22527 10029
rect 24853 10026 24919 10029
rect 22461 10024 24919 10026
rect 22461 9968 22466 10024
rect 22522 9968 24858 10024
rect 24914 9968 24919 10024
rect 22461 9966 24919 9968
rect 22461 9963 22527 9966
rect 24853 9963 24919 9966
rect 7373 9890 7439 9893
rect 9213 9890 9279 9893
rect 7373 9888 9279 9890
rect 7373 9832 7378 9888
rect 7434 9832 9218 9888
rect 9274 9832 9279 9888
rect 7373 9830 9279 9832
rect 7373 9827 7439 9830
rect 9213 9827 9279 9830
rect 9489 9890 9555 9893
rect 10685 9890 10751 9893
rect 9489 9888 10751 9890
rect 9489 9832 9494 9888
rect 9550 9832 10690 9888
rect 10746 9832 10751 9888
rect 9489 9830 10751 9832
rect 9489 9827 9555 9830
rect 10685 9827 10751 9830
rect 15561 9890 15627 9893
rect 17217 9890 17283 9893
rect 15561 9888 17283 9890
rect 15561 9832 15566 9888
rect 15622 9832 17222 9888
rect 17278 9832 17283 9888
rect 15561 9830 17283 9832
rect 15561 9827 15627 9830
rect 17217 9827 17283 9830
rect 17401 9890 17467 9893
rect 20989 9890 21055 9893
rect 17401 9888 21055 9890
rect 17401 9832 17406 9888
rect 17462 9832 20994 9888
rect 21050 9832 21055 9888
rect 17401 9830 21055 9832
rect 17401 9827 17467 9830
rect 20989 9827 21055 9830
rect 21398 9828 21404 9892
rect 21468 9890 21474 9892
rect 21541 9890 21607 9893
rect 21468 9888 21607 9890
rect 21468 9832 21546 9888
rect 21602 9832 21607 9888
rect 21468 9830 21607 9832
rect 21468 9828 21474 9830
rect 21541 9827 21607 9830
rect 22318 9828 22324 9892
rect 22388 9890 22394 9892
rect 22388 9830 22524 9890
rect 22388 9828 22394 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 22464 9757 22524 9830
rect 23054 9828 23060 9892
rect 23124 9890 23130 9892
rect 23197 9890 23263 9893
rect 23124 9888 23263 9890
rect 23124 9832 23202 9888
rect 23258 9832 23263 9888
rect 23124 9830 23263 9832
rect 23124 9828 23130 9830
rect 23197 9827 23263 9830
rect 24945 9890 25011 9893
rect 27520 9890 28000 9920
rect 24945 9888 28000 9890
rect 24945 9832 24950 9888
rect 25006 9832 28000 9888
rect 24945 9830 28000 9832
rect 24945 9827 25011 9830
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9830
rect 24277 9759 24597 9760
rect 1945 9754 2011 9757
rect 3785 9754 3851 9757
rect 1945 9752 3851 9754
rect 1945 9696 1950 9752
rect 2006 9696 3790 9752
rect 3846 9696 3851 9752
rect 1945 9694 3851 9696
rect 1945 9691 2011 9694
rect 3785 9691 3851 9694
rect 11421 9754 11487 9757
rect 14089 9754 14155 9757
rect 11421 9752 14155 9754
rect 11421 9696 11426 9752
rect 11482 9696 14094 9752
rect 14150 9696 14155 9752
rect 11421 9694 14155 9696
rect 11421 9691 11487 9694
rect 14089 9691 14155 9694
rect 17033 9754 17099 9757
rect 21357 9754 21423 9757
rect 17033 9752 21423 9754
rect 17033 9696 17038 9752
rect 17094 9696 21362 9752
rect 21418 9696 21423 9752
rect 17033 9694 21423 9696
rect 17033 9691 17099 9694
rect 21357 9691 21423 9694
rect 22461 9752 22527 9757
rect 22461 9696 22466 9752
rect 22522 9696 22527 9752
rect 22461 9691 22527 9696
rect 24669 9754 24735 9757
rect 25497 9754 25563 9757
rect 24669 9752 25563 9754
rect 24669 9696 24674 9752
rect 24730 9696 25502 9752
rect 25558 9696 25563 9752
rect 24669 9694 25563 9696
rect 24669 9691 24735 9694
rect 25497 9691 25563 9694
rect 0 9618 480 9648
rect 5257 9618 5323 9621
rect 8661 9618 8727 9621
rect 0 9558 2514 9618
rect 0 9528 480 9558
rect 2454 9482 2514 9558
rect 5257 9616 8727 9618
rect 5257 9560 5262 9616
rect 5318 9560 8666 9616
rect 8722 9560 8727 9616
rect 5257 9558 8727 9560
rect 5257 9555 5323 9558
rect 8661 9555 8727 9558
rect 10869 9618 10935 9621
rect 17493 9618 17559 9621
rect 25957 9618 26023 9621
rect 10869 9616 26023 9618
rect 10869 9560 10874 9616
rect 10930 9560 17498 9616
rect 17554 9560 25962 9616
rect 26018 9560 26023 9616
rect 10869 9558 26023 9560
rect 10869 9555 10935 9558
rect 17493 9555 17559 9558
rect 25957 9555 26023 9558
rect 2957 9482 3023 9485
rect 3509 9482 3575 9485
rect 2454 9480 3575 9482
rect 2454 9424 2962 9480
rect 3018 9424 3514 9480
rect 3570 9424 3575 9480
rect 2454 9422 3575 9424
rect 2957 9419 3023 9422
rect 3509 9419 3575 9422
rect 3785 9482 3851 9485
rect 6361 9482 6427 9485
rect 3785 9480 6427 9482
rect 3785 9424 3790 9480
rect 3846 9424 6366 9480
rect 6422 9424 6427 9480
rect 3785 9422 6427 9424
rect 3785 9419 3851 9422
rect 6361 9419 6427 9422
rect 7649 9482 7715 9485
rect 11053 9482 11119 9485
rect 7649 9480 11119 9482
rect 7649 9424 7654 9480
rect 7710 9424 11058 9480
rect 11114 9424 11119 9480
rect 7649 9422 11119 9424
rect 7649 9419 7715 9422
rect 11053 9419 11119 9422
rect 18781 9482 18847 9485
rect 20253 9482 20319 9485
rect 22277 9482 22343 9485
rect 18781 9480 20178 9482
rect 18781 9424 18786 9480
rect 18842 9424 20178 9480
rect 18781 9422 20178 9424
rect 18781 9419 18847 9422
rect 2773 9346 2839 9349
rect 6545 9346 6611 9349
rect 2773 9344 6611 9346
rect 2773 9288 2778 9344
rect 2834 9288 6550 9344
rect 6606 9288 6611 9344
rect 2773 9286 6611 9288
rect 2773 9283 2839 9286
rect 6545 9283 6611 9286
rect 9990 9284 9996 9348
rect 10060 9346 10066 9348
rect 10133 9346 10199 9349
rect 10060 9344 10199 9346
rect 10060 9288 10138 9344
rect 10194 9288 10199 9344
rect 10060 9286 10199 9288
rect 10060 9284 10066 9286
rect 10133 9283 10199 9286
rect 13813 9346 13879 9349
rect 14273 9346 14339 9349
rect 17309 9346 17375 9349
rect 13813 9344 17375 9346
rect 13813 9288 13818 9344
rect 13874 9288 14278 9344
rect 14334 9288 17314 9344
rect 17370 9288 17375 9344
rect 13813 9286 17375 9288
rect 20118 9346 20178 9422
rect 20253 9480 22343 9482
rect 20253 9424 20258 9480
rect 20314 9424 22282 9480
rect 22338 9424 22343 9480
rect 20253 9422 22343 9424
rect 20253 9419 20319 9422
rect 22277 9419 22343 9422
rect 23974 9420 23980 9484
rect 24044 9482 24050 9484
rect 24710 9482 24716 9484
rect 24044 9422 24716 9482
rect 24044 9420 24050 9422
rect 24710 9420 24716 9422
rect 24780 9420 24786 9484
rect 24669 9346 24735 9349
rect 20118 9344 24735 9346
rect 20118 9288 24674 9344
rect 24730 9288 24735 9344
rect 20118 9286 24735 9288
rect 13813 9283 13879 9286
rect 14273 9283 14339 9286
rect 17309 9283 17375 9286
rect 24669 9283 24735 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 1393 9210 1459 9213
rect 4429 9210 4495 9213
rect 1393 9208 4495 9210
rect 1393 9152 1398 9208
rect 1454 9152 4434 9208
rect 4490 9152 4495 9208
rect 1393 9150 4495 9152
rect 1393 9147 1459 9150
rect 4429 9147 4495 9150
rect 4613 9210 4679 9213
rect 8293 9210 8359 9213
rect 22001 9210 22067 9213
rect 4613 9208 8359 9210
rect 4613 9152 4618 9208
rect 4674 9152 8298 9208
rect 8354 9152 8359 9208
rect 4613 9150 8359 9152
rect 4613 9147 4679 9150
rect 8293 9147 8359 9150
rect 20164 9208 22067 9210
rect 20164 9152 22006 9208
rect 22062 9152 22067 9208
rect 20164 9150 22067 9152
rect 2681 9074 2747 9077
rect 2998 9074 3004 9076
rect 2681 9072 3004 9074
rect 2681 9016 2686 9072
rect 2742 9016 3004 9072
rect 2681 9014 3004 9016
rect 2681 9011 2747 9014
rect 2998 9012 3004 9014
rect 3068 9012 3074 9076
rect 3325 9074 3391 9077
rect 4102 9074 4108 9076
rect 3325 9072 4108 9074
rect 3325 9016 3330 9072
rect 3386 9016 4108 9072
rect 3325 9014 4108 9016
rect 3325 9011 3391 9014
rect 4102 9012 4108 9014
rect 4172 9012 4178 9076
rect 5257 9074 5323 9077
rect 6678 9074 6684 9076
rect 5257 9072 6684 9074
rect 5257 9016 5262 9072
rect 5318 9016 6684 9072
rect 5257 9014 6684 9016
rect 5257 9011 5323 9014
rect 6678 9012 6684 9014
rect 6748 9012 6754 9076
rect 7925 9074 7991 9077
rect 9857 9074 9923 9077
rect 17033 9074 17099 9077
rect 7925 9072 8954 9074
rect 7925 9016 7930 9072
rect 7986 9016 8954 9072
rect 7925 9014 8954 9016
rect 7925 9011 7991 9014
rect 0 8938 480 8968
rect 5390 8938 5396 8940
rect 0 8878 5396 8938
rect 0 8848 480 8878
rect 5390 8876 5396 8878
rect 5460 8876 5466 8940
rect 7649 8938 7715 8941
rect 8753 8938 8819 8941
rect 7649 8936 8819 8938
rect 7649 8880 7654 8936
rect 7710 8880 8758 8936
rect 8814 8880 8819 8936
rect 7649 8878 8819 8880
rect 8894 8938 8954 9014
rect 9857 9072 17099 9074
rect 9857 9016 9862 9072
rect 9918 9016 17038 9072
rect 17094 9016 17099 9072
rect 9857 9014 17099 9016
rect 9857 9011 9923 9014
rect 17033 9011 17099 9014
rect 17309 9074 17375 9077
rect 20164 9074 20224 9150
rect 22001 9147 22067 9150
rect 25129 9210 25195 9213
rect 27520 9210 28000 9240
rect 25129 9208 28000 9210
rect 25129 9152 25134 9208
rect 25190 9152 28000 9208
rect 25129 9150 28000 9152
rect 25129 9147 25195 9150
rect 27520 9120 28000 9150
rect 17309 9072 20224 9074
rect 17309 9016 17314 9072
rect 17370 9016 20224 9072
rect 17309 9014 20224 9016
rect 20989 9074 21055 9077
rect 25681 9074 25747 9077
rect 20989 9072 25747 9074
rect 20989 9016 20994 9072
rect 21050 9016 25686 9072
rect 25742 9016 25747 9072
rect 20989 9014 25747 9016
rect 17309 9011 17375 9014
rect 20989 9011 21055 9014
rect 25681 9011 25747 9014
rect 13169 8938 13235 8941
rect 13905 8940 13971 8941
rect 13854 8938 13860 8940
rect 8894 8936 13235 8938
rect 8894 8880 13174 8936
rect 13230 8880 13235 8936
rect 8894 8878 13235 8880
rect 13814 8878 13860 8938
rect 13924 8936 13971 8940
rect 15745 8938 15811 8941
rect 26325 8938 26391 8941
rect 13966 8880 13971 8936
rect 7649 8875 7715 8878
rect 8753 8875 8819 8878
rect 13169 8875 13235 8878
rect 13854 8876 13860 8878
rect 13924 8876 13971 8880
rect 13905 8875 13971 8876
rect 14598 8878 15394 8938
rect 14598 8805 14658 8878
rect 6821 8802 6887 8805
rect 7046 8802 7052 8804
rect 6821 8800 7052 8802
rect 6821 8744 6826 8800
rect 6882 8744 7052 8800
rect 6821 8742 7052 8744
rect 6821 8739 6887 8742
rect 7046 8740 7052 8742
rect 7116 8740 7122 8804
rect 7557 8802 7623 8805
rect 14365 8802 14431 8805
rect 7557 8800 14431 8802
rect 7557 8744 7562 8800
rect 7618 8744 14370 8800
rect 14426 8744 14431 8800
rect 7557 8742 14431 8744
rect 7557 8739 7623 8742
rect 14365 8739 14431 8742
rect 14549 8800 14658 8805
rect 14549 8744 14554 8800
rect 14610 8744 14658 8800
rect 14549 8742 14658 8744
rect 15334 8802 15394 8878
rect 15745 8936 26391 8938
rect 15745 8880 15750 8936
rect 15806 8880 26330 8936
rect 26386 8880 26391 8936
rect 15745 8878 26391 8880
rect 15745 8875 15811 8878
rect 26325 8875 26391 8878
rect 22001 8802 22067 8805
rect 15334 8800 22067 8802
rect 15334 8744 22006 8800
rect 22062 8744 22067 8800
rect 15334 8742 22067 8744
rect 14549 8739 14615 8742
rect 22001 8739 22067 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 6913 8666 6979 8669
rect 14641 8666 14707 8669
rect 6913 8664 14707 8666
rect 6913 8608 6918 8664
rect 6974 8608 14646 8664
rect 14702 8608 14707 8664
rect 6913 8606 14707 8608
rect 6913 8603 6979 8606
rect 14641 8603 14707 8606
rect 16205 8666 16271 8669
rect 22553 8666 22619 8669
rect 16205 8664 22619 8666
rect 16205 8608 16210 8664
rect 16266 8608 22558 8664
rect 22614 8608 22619 8664
rect 16205 8606 22619 8608
rect 16205 8603 16271 8606
rect 22553 8603 22619 8606
rect 25078 8604 25084 8668
rect 25148 8666 25154 8668
rect 27520 8666 28000 8696
rect 25148 8606 28000 8666
rect 25148 8604 25154 8606
rect 27520 8576 28000 8606
rect 1669 8530 1735 8533
rect 5441 8530 5507 8533
rect 16665 8530 16731 8533
rect 1669 8528 16731 8530
rect 1669 8472 1674 8528
rect 1730 8472 5446 8528
rect 5502 8472 16670 8528
rect 16726 8472 16731 8528
rect 1669 8470 16731 8472
rect 1669 8467 1735 8470
rect 5441 8467 5507 8470
rect 16665 8467 16731 8470
rect 16798 8468 16804 8532
rect 16868 8530 16874 8532
rect 17401 8530 17467 8533
rect 16868 8528 17467 8530
rect 16868 8472 17406 8528
rect 17462 8472 17467 8528
rect 16868 8470 17467 8472
rect 16868 8468 16874 8470
rect 17401 8467 17467 8470
rect 18781 8530 18847 8533
rect 20161 8530 20227 8533
rect 25037 8530 25103 8533
rect 18781 8528 25103 8530
rect 18781 8472 18786 8528
rect 18842 8472 20166 8528
rect 20222 8472 25042 8528
rect 25098 8472 25103 8528
rect 18781 8470 25103 8472
rect 18781 8467 18847 8470
rect 20161 8467 20227 8470
rect 25037 8467 25103 8470
rect 3141 8394 3207 8397
rect 8201 8394 8267 8397
rect 13077 8394 13143 8397
rect 16389 8394 16455 8397
rect 3141 8392 8770 8394
rect 3141 8336 3146 8392
rect 3202 8336 8206 8392
rect 8262 8336 8770 8392
rect 3141 8334 8770 8336
rect 3141 8331 3207 8334
rect 8201 8331 8267 8334
rect 0 8258 480 8288
rect 3918 8258 3924 8260
rect 0 8198 3924 8258
rect 0 8168 480 8198
rect 3918 8196 3924 8198
rect 3988 8196 3994 8260
rect 6729 8258 6795 8261
rect 8477 8258 8543 8261
rect 6729 8256 8543 8258
rect 6729 8200 6734 8256
rect 6790 8200 8482 8256
rect 8538 8200 8543 8256
rect 6729 8198 8543 8200
rect 8710 8258 8770 8334
rect 9998 8334 10748 8394
rect 9998 8258 10058 8334
rect 8710 8198 10058 8258
rect 6729 8195 6795 8198
rect 8477 8195 8543 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 2865 8122 2931 8125
rect 4061 8122 4127 8125
rect 6637 8122 6703 8125
rect 8477 8122 8543 8125
rect 2865 8120 5826 8122
rect 2865 8064 2870 8120
rect 2926 8064 4066 8120
rect 4122 8064 5826 8120
rect 2865 8062 5826 8064
rect 2865 8059 2931 8062
rect 4061 8059 4127 8062
rect 2313 7986 2379 7989
rect 5533 7986 5599 7989
rect 2313 7984 5599 7986
rect 2313 7928 2318 7984
rect 2374 7928 5538 7984
rect 5594 7928 5599 7984
rect 2313 7926 5599 7928
rect 5766 7986 5826 8062
rect 6637 8120 8543 8122
rect 6637 8064 6642 8120
rect 6698 8064 8482 8120
rect 8538 8064 8543 8120
rect 6637 8062 8543 8064
rect 10688 8122 10748 8334
rect 13077 8392 16455 8394
rect 13077 8336 13082 8392
rect 13138 8336 16394 8392
rect 16450 8336 16455 8392
rect 13077 8334 16455 8336
rect 13077 8331 13143 8334
rect 16389 8331 16455 8334
rect 19006 8332 19012 8396
rect 19076 8394 19082 8396
rect 19241 8394 19307 8397
rect 20621 8394 20687 8397
rect 21214 8394 21220 8396
rect 19076 8392 19307 8394
rect 19076 8336 19246 8392
rect 19302 8336 19307 8392
rect 19076 8334 19307 8336
rect 19076 8332 19082 8334
rect 19241 8331 19307 8334
rect 19382 8334 20178 8394
rect 11145 8292 11211 8295
rect 11102 8290 11211 8292
rect 11102 8260 11150 8290
rect 11094 8258 11100 8260
rect 11088 8198 11100 8258
rect 11206 8234 11211 8290
rect 11094 8196 11100 8198
rect 11164 8229 11211 8234
rect 12433 8258 12499 8261
rect 19382 8258 19442 8334
rect 12433 8256 19442 8258
rect 11164 8196 11170 8229
rect 12433 8200 12438 8256
rect 12494 8200 19442 8256
rect 12433 8198 19442 8200
rect 20118 8258 20178 8334
rect 20621 8392 21220 8394
rect 20621 8336 20626 8392
rect 20682 8336 21220 8392
rect 20621 8334 21220 8336
rect 20621 8331 20687 8334
rect 21214 8332 21220 8334
rect 21284 8332 21290 8396
rect 22093 8394 22159 8397
rect 22502 8394 22508 8396
rect 22093 8392 22508 8394
rect 22093 8336 22098 8392
rect 22154 8336 22508 8392
rect 22093 8334 22508 8336
rect 22093 8331 22159 8334
rect 22502 8332 22508 8334
rect 22572 8332 22578 8396
rect 21265 8258 21331 8261
rect 20118 8256 21331 8258
rect 20118 8200 21270 8256
rect 21326 8200 21331 8256
rect 20118 8198 21331 8200
rect 12433 8195 12499 8198
rect 21265 8195 21331 8198
rect 21582 8196 21588 8260
rect 21652 8258 21658 8260
rect 21725 8258 21791 8261
rect 21652 8256 21791 8258
rect 21652 8200 21730 8256
rect 21786 8200 21791 8256
rect 21652 8198 21791 8200
rect 21652 8196 21658 8198
rect 21725 8195 21791 8198
rect 23606 8196 23612 8260
rect 23676 8258 23682 8260
rect 24710 8258 24716 8260
rect 23676 8198 24716 8258
rect 23676 8196 23682 8198
rect 24710 8196 24716 8198
rect 24780 8258 24786 8260
rect 25681 8258 25747 8261
rect 24780 8256 25747 8258
rect 24780 8200 25686 8256
rect 25742 8200 25747 8256
rect 24780 8198 25747 8200
rect 24780 8196 24786 8198
rect 25681 8195 25747 8198
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 19241 8122 19307 8125
rect 10688 8120 19307 8122
rect 10688 8064 19246 8120
rect 19302 8064 19307 8120
rect 10688 8062 19307 8064
rect 6637 8059 6703 8062
rect 8477 8059 8543 8062
rect 19241 8059 19307 8062
rect 22553 8122 22619 8125
rect 23013 8122 23079 8125
rect 27520 8122 28000 8152
rect 22553 8120 23079 8122
rect 22553 8064 22558 8120
rect 22614 8064 23018 8120
rect 23074 8064 23079 8120
rect 22553 8062 23079 8064
rect 22553 8059 22619 8062
rect 23013 8059 23079 8062
rect 25638 8062 28000 8122
rect 11053 7986 11119 7989
rect 5766 7984 11119 7986
rect 5766 7928 11058 7984
rect 11114 7928 11119 7984
rect 5766 7926 11119 7928
rect 2313 7923 2379 7926
rect 5533 7923 5599 7926
rect 11053 7923 11119 7926
rect 13537 7986 13603 7989
rect 16021 7986 16087 7989
rect 25405 7986 25471 7989
rect 13537 7984 25471 7986
rect 13537 7928 13542 7984
rect 13598 7928 16026 7984
rect 16082 7928 25410 7984
rect 25466 7928 25471 7984
rect 13537 7926 25471 7928
rect 13537 7923 13603 7926
rect 16021 7923 16087 7926
rect 25405 7923 25471 7926
rect 4889 7850 4955 7853
rect 8293 7850 8359 7853
rect 10777 7852 10843 7853
rect 4889 7848 8359 7850
rect 4889 7792 4894 7848
rect 4950 7792 8298 7848
rect 8354 7792 8359 7848
rect 4889 7790 8359 7792
rect 4889 7787 4955 7790
rect 8293 7787 8359 7790
rect 10726 7788 10732 7852
rect 10796 7850 10843 7852
rect 14917 7850 14983 7853
rect 22277 7850 22343 7853
rect 23565 7850 23631 7853
rect 10796 7848 10888 7850
rect 10838 7792 10888 7848
rect 10796 7790 10888 7792
rect 14917 7848 23631 7850
rect 14917 7792 14922 7848
rect 14978 7792 22282 7848
rect 22338 7792 23570 7848
rect 23626 7792 23631 7848
rect 14917 7790 23631 7792
rect 10796 7788 10843 7790
rect 10777 7787 10843 7788
rect 14917 7787 14983 7790
rect 22277 7787 22343 7790
rect 23565 7787 23631 7790
rect 23974 7788 23980 7852
rect 24044 7850 24050 7852
rect 25638 7850 25698 8062
rect 27520 8032 28000 8062
rect 24044 7790 25698 7850
rect 24044 7788 24050 7790
rect 3509 7714 3575 7717
rect 5441 7714 5507 7717
rect 3509 7712 5507 7714
rect 3509 7656 3514 7712
rect 3570 7656 5446 7712
rect 5502 7656 5507 7712
rect 3509 7654 5507 7656
rect 3509 7651 3575 7654
rect 5441 7651 5507 7654
rect 6637 7714 6703 7717
rect 11881 7714 11947 7717
rect 6637 7712 11947 7714
rect 6637 7656 6642 7712
rect 6698 7656 11886 7712
rect 11942 7656 11947 7712
rect 6637 7654 11947 7656
rect 6637 7651 6703 7654
rect 11881 7651 11947 7654
rect 13169 7714 13235 7717
rect 14222 7714 14228 7716
rect 13169 7712 14228 7714
rect 13169 7656 13174 7712
rect 13230 7656 14228 7712
rect 13169 7654 14228 7656
rect 13169 7651 13235 7654
rect 14222 7652 14228 7654
rect 14292 7652 14298 7716
rect 16113 7714 16179 7717
rect 18597 7714 18663 7717
rect 16113 7712 18663 7714
rect 16113 7656 16118 7712
rect 16174 7656 18602 7712
rect 18658 7656 18663 7712
rect 16113 7654 18663 7656
rect 16113 7651 16179 7654
rect 18597 7651 18663 7654
rect 19333 7714 19399 7717
rect 20345 7714 20411 7717
rect 19333 7712 20411 7714
rect 19333 7656 19338 7712
rect 19394 7656 20350 7712
rect 20406 7656 20411 7712
rect 19333 7654 20411 7656
rect 19333 7651 19399 7654
rect 20345 7651 20411 7654
rect 20478 7652 20484 7716
rect 20548 7714 20554 7716
rect 21817 7714 21883 7717
rect 22737 7714 22803 7717
rect 20548 7654 21420 7714
rect 20548 7652 20554 7654
rect 5610 7648 5930 7649
rect 0 7578 480 7608
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 2129 7578 2195 7581
rect 0 7576 2195 7578
rect 0 7520 2134 7576
rect 2190 7520 2195 7576
rect 0 7518 2195 7520
rect 0 7488 480 7518
rect 2129 7515 2195 7518
rect 6126 7516 6132 7580
rect 6196 7578 6202 7580
rect 6821 7578 6887 7581
rect 6196 7576 6887 7578
rect 6196 7520 6826 7576
rect 6882 7520 6887 7576
rect 6196 7518 6887 7520
rect 6196 7516 6202 7518
rect 6821 7515 6887 7518
rect 9581 7578 9647 7581
rect 10409 7578 10475 7581
rect 9581 7576 10475 7578
rect 9581 7520 9586 7576
rect 9642 7520 10414 7576
rect 10470 7520 10475 7576
rect 9581 7518 10475 7520
rect 9581 7515 9647 7518
rect 10409 7515 10475 7518
rect 18229 7578 18295 7581
rect 20713 7578 20779 7581
rect 18229 7576 20779 7578
rect 18229 7520 18234 7576
rect 18290 7520 20718 7576
rect 20774 7520 20779 7576
rect 18229 7518 20779 7520
rect 18229 7515 18295 7518
rect 20713 7515 20779 7518
rect 4797 7442 4863 7445
rect 9213 7442 9279 7445
rect 4797 7440 9279 7442
rect 4797 7384 4802 7440
rect 4858 7384 9218 7440
rect 9274 7384 9279 7440
rect 4797 7382 9279 7384
rect 4797 7379 4863 7382
rect 9213 7379 9279 7382
rect 9765 7442 9831 7445
rect 17401 7442 17467 7445
rect 9765 7440 17467 7442
rect 9765 7384 9770 7440
rect 9826 7384 17406 7440
rect 17462 7384 17467 7440
rect 9765 7382 17467 7384
rect 9765 7379 9831 7382
rect 17401 7379 17467 7382
rect 18597 7442 18663 7445
rect 21360 7442 21420 7654
rect 21817 7712 22803 7714
rect 21817 7656 21822 7712
rect 21878 7656 22742 7712
rect 22798 7656 22803 7712
rect 21817 7654 22803 7656
rect 21817 7651 21883 7654
rect 22737 7651 22803 7654
rect 23197 7714 23263 7717
rect 23473 7714 23539 7717
rect 23197 7712 23539 7714
rect 23197 7656 23202 7712
rect 23258 7656 23478 7712
rect 23534 7656 23539 7712
rect 23197 7654 23539 7656
rect 23197 7651 23263 7654
rect 23473 7651 23539 7654
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 21817 7578 21883 7581
rect 23473 7578 23539 7581
rect 27520 7578 28000 7608
rect 21817 7576 23539 7578
rect 21817 7520 21822 7576
rect 21878 7520 23478 7576
rect 23534 7520 23539 7576
rect 21817 7518 23539 7520
rect 21817 7515 21883 7518
rect 23473 7515 23539 7518
rect 24718 7518 28000 7578
rect 22185 7442 22251 7445
rect 23197 7442 23263 7445
rect 18597 7440 21282 7442
rect 18597 7384 18602 7440
rect 18658 7384 21282 7440
rect 18597 7382 21282 7384
rect 21360 7440 22251 7442
rect 21360 7384 22190 7440
rect 22246 7384 22251 7440
rect 21360 7382 22251 7384
rect 18597 7379 18663 7382
rect 12249 7306 12315 7309
rect 16941 7306 17007 7309
rect 4846 7246 12128 7306
rect 0 7034 480 7064
rect 4846 7034 4906 7246
rect 4981 7170 5047 7173
rect 8661 7170 8727 7173
rect 4981 7168 8727 7170
rect 4981 7112 4986 7168
rect 5042 7112 8666 7168
rect 8722 7112 8727 7168
rect 4981 7110 8727 7112
rect 12068 7170 12128 7246
rect 12249 7304 17007 7306
rect 12249 7248 12254 7304
rect 12310 7248 16946 7304
rect 17002 7248 17007 7304
rect 12249 7246 17007 7248
rect 12249 7243 12315 7246
rect 16941 7243 17007 7246
rect 18413 7306 18479 7309
rect 20989 7306 21055 7309
rect 18413 7304 21055 7306
rect 18413 7248 18418 7304
rect 18474 7248 20994 7304
rect 21050 7248 21055 7304
rect 18413 7246 21055 7248
rect 18413 7243 18479 7246
rect 20989 7243 21055 7246
rect 15377 7170 15443 7173
rect 12068 7168 15443 7170
rect 12068 7112 15382 7168
rect 15438 7112 15443 7168
rect 12068 7110 15443 7112
rect 4981 7107 5047 7110
rect 8661 7107 8727 7110
rect 15377 7107 15443 7110
rect 15745 7170 15811 7173
rect 19241 7170 19307 7173
rect 15745 7168 19307 7170
rect 15745 7112 15750 7168
rect 15806 7112 19246 7168
rect 19302 7112 19307 7168
rect 15745 7110 19307 7112
rect 21222 7170 21282 7382
rect 22185 7379 22251 7382
rect 23062 7440 23263 7442
rect 23062 7384 23202 7440
rect 23258 7384 23263 7440
rect 23062 7382 23263 7384
rect 21449 7306 21515 7309
rect 23062 7306 23122 7382
rect 23197 7379 23263 7382
rect 23422 7380 23428 7444
rect 23492 7442 23498 7444
rect 24718 7442 24778 7518
rect 27520 7488 28000 7518
rect 23492 7382 24778 7442
rect 23492 7380 23498 7382
rect 21449 7304 23122 7306
rect 21449 7248 21454 7304
rect 21510 7248 23122 7304
rect 21449 7246 23122 7248
rect 23289 7306 23355 7309
rect 24945 7306 25011 7309
rect 23289 7304 25011 7306
rect 23289 7248 23294 7304
rect 23350 7248 24950 7304
rect 25006 7248 25011 7304
rect 23289 7246 25011 7248
rect 21449 7243 21515 7246
rect 23289 7243 23355 7246
rect 24945 7243 25011 7246
rect 23473 7170 23539 7173
rect 21222 7168 23539 7170
rect 21222 7112 23478 7168
rect 23534 7112 23539 7168
rect 21222 7110 23539 7112
rect 15745 7107 15811 7110
rect 19241 7107 19307 7110
rect 23473 7107 23539 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 0 6974 4906 7034
rect 5165 7034 5231 7037
rect 7925 7034 7991 7037
rect 5165 7032 7991 7034
rect 5165 6976 5170 7032
rect 5226 6976 7930 7032
rect 7986 6976 7991 7032
rect 5165 6974 7991 6976
rect 0 6944 480 6974
rect 5165 6971 5231 6974
rect 7925 6971 7991 6974
rect 14917 7034 14983 7037
rect 14917 7032 19396 7034
rect 14917 6976 14922 7032
rect 14978 6976 19396 7032
rect 14917 6974 19396 6976
rect 14917 6971 14983 6974
rect 2497 6898 2563 6901
rect 5073 6898 5139 6901
rect 8753 6898 8819 6901
rect 2497 6896 5139 6898
rect 2497 6840 2502 6896
rect 2558 6840 5078 6896
rect 5134 6840 5139 6896
rect 2497 6838 5139 6840
rect 2497 6835 2563 6838
rect 5073 6835 5139 6838
rect 5214 6896 8819 6898
rect 5214 6840 8758 6896
rect 8814 6840 8819 6896
rect 5214 6838 8819 6840
rect 1761 6762 1827 6765
rect 5214 6762 5274 6838
rect 8753 6835 8819 6838
rect 10726 6836 10732 6900
rect 10796 6898 10802 6900
rect 14365 6898 14431 6901
rect 10796 6896 14431 6898
rect 10796 6840 14370 6896
rect 14426 6840 14431 6896
rect 10796 6838 14431 6840
rect 19336 6898 19396 6974
rect 20110 6972 20116 7036
rect 20180 7034 20186 7036
rect 20345 7034 20411 7037
rect 20180 7032 20411 7034
rect 20180 6976 20350 7032
rect 20406 6976 20411 7032
rect 20180 6974 20411 6976
rect 20180 6972 20186 6974
rect 20345 6971 20411 6974
rect 21541 7034 21607 7037
rect 24577 7034 24643 7037
rect 21541 7032 24643 7034
rect 21541 6976 21546 7032
rect 21602 6976 24582 7032
rect 24638 6976 24643 7032
rect 21541 6974 24643 6976
rect 21541 6971 21607 6974
rect 24577 6971 24643 6974
rect 25129 7034 25195 7037
rect 27520 7034 28000 7064
rect 25129 7032 28000 7034
rect 25129 6976 25134 7032
rect 25190 6976 28000 7032
rect 25129 6974 28000 6976
rect 25129 6971 25195 6974
rect 27520 6944 28000 6974
rect 20805 6898 20871 6901
rect 19336 6896 20871 6898
rect 19336 6840 20810 6896
rect 20866 6840 20871 6896
rect 19336 6838 20871 6840
rect 10796 6836 10802 6838
rect 14365 6835 14431 6838
rect 20805 6835 20871 6838
rect 20989 6898 21055 6901
rect 25405 6898 25471 6901
rect 20989 6896 25471 6898
rect 20989 6840 20994 6896
rect 21050 6840 25410 6896
rect 25466 6840 25471 6896
rect 20989 6838 25471 6840
rect 20989 6835 21055 6838
rect 25405 6835 25471 6838
rect 1761 6760 5274 6762
rect 1761 6704 1766 6760
rect 1822 6704 5274 6760
rect 1761 6702 5274 6704
rect 5441 6762 5507 6765
rect 7373 6762 7439 6765
rect 8150 6762 8156 6764
rect 5441 6760 6194 6762
rect 5441 6704 5446 6760
rect 5502 6704 6194 6760
rect 5441 6702 6194 6704
rect 1761 6699 1827 6702
rect 5441 6699 5507 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 6134 6490 6194 6702
rect 7373 6760 8156 6762
rect 7373 6704 7378 6760
rect 7434 6704 8156 6760
rect 7373 6702 8156 6704
rect 7373 6699 7439 6702
rect 8150 6700 8156 6702
rect 8220 6700 8226 6764
rect 8661 6762 8727 6765
rect 8937 6762 9003 6765
rect 8661 6760 9003 6762
rect 8661 6704 8666 6760
rect 8722 6704 8942 6760
rect 8998 6704 9003 6760
rect 8661 6702 9003 6704
rect 8661 6699 8727 6702
rect 8937 6699 9003 6702
rect 12198 6700 12204 6764
rect 12268 6762 12274 6764
rect 12433 6762 12499 6765
rect 12268 6760 12499 6762
rect 12268 6704 12438 6760
rect 12494 6704 12499 6760
rect 12268 6702 12499 6704
rect 12268 6700 12274 6702
rect 12433 6699 12499 6702
rect 16481 6762 16547 6765
rect 19793 6762 19859 6765
rect 16481 6760 19859 6762
rect 16481 6704 16486 6760
rect 16542 6704 19798 6760
rect 19854 6704 19859 6760
rect 16481 6702 19859 6704
rect 16481 6699 16547 6702
rect 19793 6699 19859 6702
rect 19977 6762 20043 6765
rect 25773 6762 25839 6765
rect 19977 6760 25839 6762
rect 19977 6704 19982 6760
rect 20038 6704 25778 6760
rect 25834 6704 25839 6760
rect 19977 6702 25839 6704
rect 19977 6699 20043 6702
rect 25773 6699 25839 6702
rect 7925 6626 7991 6629
rect 11053 6626 11119 6629
rect 7925 6624 11119 6626
rect 7925 6568 7930 6624
rect 7986 6568 11058 6624
rect 11114 6568 11119 6624
rect 7925 6566 11119 6568
rect 7925 6563 7991 6566
rect 11053 6563 11119 6566
rect 17585 6626 17651 6629
rect 20253 6626 20319 6629
rect 17585 6624 20319 6626
rect 17585 6568 17590 6624
rect 17646 6568 20258 6624
rect 20314 6568 20319 6624
rect 17585 6566 20319 6568
rect 17585 6563 17651 6566
rect 20253 6563 20319 6566
rect 21541 6626 21607 6629
rect 23197 6626 23263 6629
rect 21541 6624 23263 6626
rect 21541 6568 21546 6624
rect 21602 6568 23202 6624
rect 23258 6568 23263 6624
rect 21541 6566 23263 6568
rect 21541 6563 21607 6566
rect 23197 6563 23263 6566
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 6913 6490 6979 6493
rect 11789 6490 11855 6493
rect 6134 6488 11855 6490
rect 6134 6432 6918 6488
rect 6974 6432 11794 6488
rect 11850 6432 11855 6488
rect 6134 6430 11855 6432
rect 6913 6427 6979 6430
rect 11789 6427 11855 6430
rect 18505 6490 18571 6493
rect 21541 6490 21607 6493
rect 27520 6490 28000 6520
rect 18505 6488 21607 6490
rect 18505 6432 18510 6488
rect 18566 6432 21546 6488
rect 21602 6432 21607 6488
rect 18505 6430 21607 6432
rect 18505 6427 18571 6430
rect 21541 6427 21607 6430
rect 26190 6430 28000 6490
rect 0 6354 480 6384
rect 3141 6354 3207 6357
rect 0 6352 3207 6354
rect 0 6296 3146 6352
rect 3202 6296 3207 6352
rect 0 6294 3207 6296
rect 0 6264 480 6294
rect 3141 6291 3207 6294
rect 5073 6354 5139 6357
rect 11329 6354 11395 6357
rect 5073 6352 11395 6354
rect 5073 6296 5078 6352
rect 5134 6296 11334 6352
rect 11390 6296 11395 6352
rect 5073 6294 11395 6296
rect 5073 6291 5139 6294
rect 11329 6291 11395 6294
rect 15469 6354 15535 6357
rect 19977 6354 20043 6357
rect 15469 6352 20043 6354
rect 15469 6296 15474 6352
rect 15530 6296 19982 6352
rect 20038 6296 20043 6352
rect 15469 6294 20043 6296
rect 15469 6291 15535 6294
rect 19977 6291 20043 6294
rect 21265 6354 21331 6357
rect 25957 6354 26023 6357
rect 21265 6352 26023 6354
rect 21265 6296 21270 6352
rect 21326 6296 25962 6352
rect 26018 6296 26023 6352
rect 21265 6294 26023 6296
rect 21265 6291 21331 6294
rect 25957 6291 26023 6294
rect 4797 6218 4863 6221
rect 8569 6218 8635 6221
rect 4797 6216 8635 6218
rect 4797 6160 4802 6216
rect 4858 6160 8574 6216
rect 8630 6160 8635 6216
rect 4797 6158 8635 6160
rect 4797 6155 4863 6158
rect 8569 6155 8635 6158
rect 9765 6218 9831 6221
rect 16297 6218 16363 6221
rect 9765 6216 16363 6218
rect 9765 6160 9770 6216
rect 9826 6160 16302 6216
rect 16358 6160 16363 6216
rect 9765 6158 16363 6160
rect 9765 6155 9831 6158
rect 16297 6155 16363 6158
rect 19701 6218 19767 6221
rect 19701 6216 23904 6218
rect 19701 6160 19706 6216
rect 19762 6160 23904 6216
rect 19701 6158 23904 6160
rect 19701 6155 19767 6158
rect 23844 6082 23904 6158
rect 23974 6156 23980 6220
rect 24044 6218 24050 6220
rect 26190 6218 26250 6430
rect 27520 6400 28000 6430
rect 24044 6158 26250 6218
rect 24044 6156 24050 6158
rect 25865 6082 25931 6085
rect 23844 6080 25931 6082
rect 23844 6024 25870 6080
rect 25926 6024 25931 6080
rect 23844 6022 25931 6024
rect 25865 6019 25931 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 4153 5946 4219 5949
rect 8661 5946 8727 5949
rect 4153 5944 8727 5946
rect 4153 5888 4158 5944
rect 4214 5888 8666 5944
rect 8722 5888 8727 5944
rect 4153 5886 8727 5888
rect 4153 5883 4219 5886
rect 8661 5883 8727 5886
rect 12433 5946 12499 5949
rect 17217 5946 17283 5949
rect 12433 5944 17283 5946
rect 12433 5888 12438 5944
rect 12494 5888 17222 5944
rect 17278 5888 17283 5944
rect 12433 5886 17283 5888
rect 12433 5883 12499 5886
rect 17217 5883 17283 5886
rect 22829 5946 22895 5949
rect 27520 5946 28000 5976
rect 22829 5944 28000 5946
rect 22829 5888 22834 5944
rect 22890 5888 28000 5944
rect 22829 5886 28000 5888
rect 22829 5883 22895 5886
rect 27520 5856 28000 5886
rect 1485 5810 1551 5813
rect 5165 5810 5231 5813
rect 1485 5808 5231 5810
rect 1485 5752 1490 5808
rect 1546 5752 5170 5808
rect 5226 5752 5231 5808
rect 1485 5750 5231 5752
rect 1485 5747 1551 5750
rect 5165 5747 5231 5750
rect 5390 5748 5396 5812
rect 5460 5810 5466 5812
rect 5901 5810 5967 5813
rect 5460 5808 5967 5810
rect 5460 5752 5906 5808
rect 5962 5752 5967 5808
rect 5460 5750 5967 5752
rect 5460 5748 5466 5750
rect 5901 5747 5967 5750
rect 6913 5810 6979 5813
rect 11605 5810 11671 5813
rect 18045 5810 18111 5813
rect 6913 5808 10794 5810
rect 6913 5752 6918 5808
rect 6974 5752 10794 5808
rect 6913 5750 10794 5752
rect 6913 5747 6979 5750
rect 0 5674 480 5704
rect 2773 5674 2839 5677
rect 0 5672 2839 5674
rect 0 5616 2778 5672
rect 2834 5616 2839 5672
rect 0 5614 2839 5616
rect 0 5584 480 5614
rect 2773 5611 2839 5614
rect 2957 5674 3023 5677
rect 3182 5674 3188 5676
rect 2957 5672 3188 5674
rect 2957 5616 2962 5672
rect 3018 5616 3188 5672
rect 2957 5614 3188 5616
rect 2957 5611 3023 5614
rect 3182 5612 3188 5614
rect 3252 5612 3258 5676
rect 10734 5674 10794 5750
rect 11605 5808 18111 5810
rect 11605 5752 11610 5808
rect 11666 5752 18050 5808
rect 18106 5752 18111 5808
rect 11605 5750 18111 5752
rect 11605 5747 11671 5750
rect 18045 5747 18111 5750
rect 18597 5810 18663 5813
rect 26325 5810 26391 5813
rect 18597 5808 26391 5810
rect 18597 5752 18602 5808
rect 18658 5752 26330 5808
rect 26386 5752 26391 5808
rect 18597 5750 26391 5752
rect 18597 5747 18663 5750
rect 26325 5747 26391 5750
rect 10910 5674 10916 5676
rect 10734 5614 10916 5674
rect 10910 5612 10916 5614
rect 10980 5674 10986 5676
rect 11605 5674 11671 5677
rect 11789 5674 11855 5677
rect 10980 5672 11855 5674
rect 10980 5616 11610 5672
rect 11666 5616 11794 5672
rect 11850 5616 11855 5672
rect 10980 5614 11855 5616
rect 10980 5612 10986 5614
rect 11605 5611 11671 5614
rect 11789 5611 11855 5614
rect 16481 5674 16547 5677
rect 18413 5674 18479 5677
rect 16481 5672 18479 5674
rect 16481 5616 16486 5672
rect 16542 5616 18418 5672
rect 18474 5616 18479 5672
rect 16481 5614 18479 5616
rect 16481 5611 16547 5614
rect 18413 5611 18479 5614
rect 18597 5674 18663 5677
rect 25129 5674 25195 5677
rect 18597 5672 25195 5674
rect 18597 5616 18602 5672
rect 18658 5616 25134 5672
rect 25190 5616 25195 5672
rect 18597 5614 25195 5616
rect 18597 5611 18663 5614
rect 25129 5611 25195 5614
rect 9438 5476 9444 5540
rect 9508 5538 9514 5540
rect 9673 5538 9739 5541
rect 9508 5536 9739 5538
rect 9508 5480 9678 5536
rect 9734 5480 9739 5536
rect 9508 5478 9739 5480
rect 9508 5476 9514 5478
rect 9673 5475 9739 5478
rect 9990 5476 9996 5540
rect 10060 5538 10066 5540
rect 12801 5538 12867 5541
rect 17585 5538 17651 5541
rect 10060 5536 12867 5538
rect 10060 5480 12806 5536
rect 12862 5480 12867 5536
rect 10060 5478 12867 5480
rect 10060 5476 10066 5478
rect 12801 5475 12867 5478
rect 15334 5536 17651 5538
rect 15334 5480 17590 5536
rect 17646 5480 17651 5536
rect 15334 5478 17651 5480
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 12985 5402 13051 5405
rect 13118 5402 13124 5404
rect 12985 5400 13124 5402
rect 12985 5344 12990 5400
rect 13046 5344 13124 5400
rect 12985 5342 13124 5344
rect 12985 5339 13051 5342
rect 13118 5340 13124 5342
rect 13188 5340 13194 5404
rect 3877 5266 3943 5269
rect 6361 5266 6427 5269
rect 3877 5264 6427 5266
rect 3877 5208 3882 5264
rect 3938 5208 6366 5264
rect 6422 5208 6427 5264
rect 3877 5206 6427 5208
rect 3877 5203 3943 5206
rect 6361 5203 6427 5206
rect 11697 5266 11763 5269
rect 15334 5266 15394 5478
rect 17585 5475 17651 5478
rect 17769 5538 17835 5541
rect 18321 5538 18387 5541
rect 17769 5536 18387 5538
rect 17769 5480 17774 5536
rect 17830 5480 18326 5536
rect 18382 5480 18387 5536
rect 17769 5478 18387 5480
rect 17769 5475 17835 5478
rect 18321 5475 18387 5478
rect 18505 5538 18571 5541
rect 18505 5536 24088 5538
rect 18505 5480 18510 5536
rect 18566 5480 24088 5536
rect 18505 5478 24088 5480
rect 18505 5475 18571 5478
rect 22829 5402 22895 5405
rect 11697 5264 15394 5266
rect 11697 5208 11702 5264
rect 11758 5208 15394 5264
rect 11697 5206 15394 5208
rect 17174 5400 22895 5402
rect 17174 5344 22834 5400
rect 22890 5344 22895 5400
rect 17174 5342 22895 5344
rect 11697 5203 11763 5206
rect 4613 5130 4679 5133
rect 8753 5130 8819 5133
rect 17174 5130 17234 5342
rect 22829 5339 22895 5342
rect 19333 5266 19399 5269
rect 24028 5266 24088 5478
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 24894 5340 24900 5404
rect 24964 5402 24970 5404
rect 25773 5402 25839 5405
rect 27520 5402 28000 5432
rect 24964 5400 28000 5402
rect 24964 5344 25778 5400
rect 25834 5344 28000 5400
rect 24964 5342 28000 5344
rect 24964 5340 24970 5342
rect 25773 5339 25839 5342
rect 27520 5312 28000 5342
rect 26233 5266 26299 5269
rect 19333 5264 23904 5266
rect 19333 5208 19338 5264
rect 19394 5208 23904 5264
rect 19333 5206 23904 5208
rect 24028 5264 26299 5266
rect 24028 5208 26238 5264
rect 26294 5208 26299 5264
rect 24028 5206 26299 5208
rect 19333 5203 19399 5206
rect 4613 5128 17234 5130
rect 4613 5072 4618 5128
rect 4674 5072 8758 5128
rect 8814 5072 17234 5128
rect 4613 5070 17234 5072
rect 17309 5130 17375 5133
rect 18597 5130 18663 5133
rect 17309 5128 20178 5130
rect 17309 5072 17314 5128
rect 17370 5072 18602 5128
rect 18658 5072 20178 5128
rect 17309 5070 20178 5072
rect 4613 5067 4679 5070
rect 8753 5067 8819 5070
rect 17309 5067 17375 5070
rect 18597 5067 18663 5070
rect 0 4994 480 5024
rect 3969 4994 4035 4997
rect 0 4992 4035 4994
rect 0 4936 3974 4992
rect 4030 4936 4035 4992
rect 0 4934 4035 4936
rect 0 4904 480 4934
rect 3969 4931 4035 4934
rect 12433 4994 12499 4997
rect 13997 4994 14063 4997
rect 15653 4994 15719 4997
rect 12433 4992 15719 4994
rect 12433 4936 12438 4992
rect 12494 4936 14002 4992
rect 14058 4936 15658 4992
rect 15714 4936 15719 4992
rect 12433 4934 15719 4936
rect 20118 4994 20178 5070
rect 20846 5068 20852 5132
rect 20916 5130 20922 5132
rect 21398 5130 21404 5132
rect 20916 5070 21404 5130
rect 20916 5068 20922 5070
rect 21398 5068 21404 5070
rect 21468 5130 21474 5132
rect 21909 5130 21975 5133
rect 21468 5128 21975 5130
rect 21468 5072 21914 5128
rect 21970 5072 21975 5128
rect 21468 5070 21975 5072
rect 21468 5068 21474 5070
rect 21909 5067 21975 5070
rect 22134 5068 22140 5132
rect 22204 5130 22210 5132
rect 22277 5130 22343 5133
rect 22204 5128 22343 5130
rect 22204 5072 22282 5128
rect 22338 5072 22343 5128
rect 22204 5070 22343 5072
rect 23844 5130 23904 5206
rect 26233 5203 26299 5206
rect 25221 5130 25287 5133
rect 23844 5128 25287 5130
rect 23844 5072 25226 5128
rect 25282 5072 25287 5128
rect 23844 5070 25287 5072
rect 22204 5068 22210 5070
rect 22277 5067 22343 5070
rect 25221 5067 25287 5070
rect 26233 4994 26299 4997
rect 20118 4992 26299 4994
rect 20118 4936 26238 4992
rect 26294 4936 26299 4992
rect 20118 4934 26299 4936
rect 12433 4931 12499 4934
rect 13997 4931 14063 4934
rect 15653 4931 15719 4934
rect 26233 4931 26299 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 2957 4858 3023 4861
rect 3550 4858 3556 4860
rect 2957 4856 3556 4858
rect 2957 4800 2962 4856
rect 3018 4800 3556 4856
rect 2957 4798 3556 4800
rect 2957 4795 3023 4798
rect 3550 4796 3556 4798
rect 3620 4858 3626 4860
rect 5073 4858 5139 4861
rect 3620 4856 5139 4858
rect 3620 4800 5078 4856
rect 5134 4800 5139 4856
rect 3620 4798 5139 4800
rect 3620 4796 3626 4798
rect 5073 4795 5139 4798
rect 5257 4858 5323 4861
rect 6494 4858 6500 4860
rect 5257 4856 6500 4858
rect 5257 4800 5262 4856
rect 5318 4800 6500 4856
rect 5257 4798 6500 4800
rect 5257 4795 5323 4798
rect 6494 4796 6500 4798
rect 6564 4858 6570 4860
rect 9857 4858 9923 4861
rect 6564 4856 9923 4858
rect 6564 4800 9862 4856
rect 9918 4800 9923 4856
rect 6564 4798 9923 4800
rect 6564 4796 6570 4798
rect 9857 4795 9923 4798
rect 10777 4858 10843 4861
rect 13077 4858 13143 4861
rect 10777 4856 13143 4858
rect 10777 4800 10782 4856
rect 10838 4800 13082 4856
rect 13138 4800 13143 4856
rect 10777 4798 13143 4800
rect 10777 4795 10843 4798
rect 13077 4795 13143 4798
rect 14590 4796 14596 4860
rect 14660 4858 14666 4860
rect 19425 4858 19491 4861
rect 14660 4856 19491 4858
rect 14660 4800 19430 4856
rect 19486 4800 19491 4856
rect 14660 4798 19491 4800
rect 14660 4796 14666 4798
rect 19425 4795 19491 4798
rect 25497 4858 25563 4861
rect 25497 4856 26802 4858
rect 25497 4800 25502 4856
rect 25558 4800 26802 4856
rect 25497 4798 26802 4800
rect 25497 4795 25563 4798
rect 2037 4722 2103 4725
rect 8753 4722 8819 4725
rect 10041 4722 10107 4725
rect 2037 4720 10107 4722
rect 2037 4664 2042 4720
rect 2098 4664 8758 4720
rect 8814 4664 10046 4720
rect 10102 4664 10107 4720
rect 2037 4662 10107 4664
rect 2037 4659 2103 4662
rect 8753 4659 8819 4662
rect 10041 4659 10107 4662
rect 12157 4722 12223 4725
rect 12433 4722 12499 4725
rect 12157 4720 12499 4722
rect 12157 4664 12162 4720
rect 12218 4664 12438 4720
rect 12494 4664 12499 4720
rect 12157 4662 12499 4664
rect 12157 4659 12223 4662
rect 12433 4659 12499 4662
rect 12617 4722 12683 4725
rect 23013 4722 23079 4725
rect 12617 4720 23079 4722
rect 12617 4664 12622 4720
rect 12678 4664 23018 4720
rect 23074 4664 23079 4720
rect 12617 4662 23079 4664
rect 26742 4722 26802 4798
rect 27520 4722 28000 4752
rect 26742 4662 28000 4722
rect 12617 4659 12683 4662
rect 23013 4659 23079 4662
rect 27520 4632 28000 4662
rect 6453 4586 6519 4589
rect 7741 4586 7807 4589
rect 20989 4586 21055 4589
rect 26325 4586 26391 4589
rect 6453 4584 21055 4586
rect 6453 4528 6458 4584
rect 6514 4528 7746 4584
rect 7802 4528 20994 4584
rect 21050 4528 21055 4584
rect 6453 4526 21055 4528
rect 6453 4523 6519 4526
rect 7741 4523 7807 4526
rect 20989 4523 21055 4526
rect 22832 4584 26391 4586
rect 22832 4528 26330 4584
rect 26386 4528 26391 4584
rect 22832 4526 26391 4528
rect 3877 4450 3943 4453
rect 9581 4450 9647 4453
rect 1902 4448 3943 4450
rect 1902 4392 3882 4448
rect 3938 4392 3943 4448
rect 1902 4390 3943 4392
rect 0 4314 480 4344
rect 1902 4314 1962 4390
rect 3877 4387 3943 4390
rect 6134 4448 9647 4450
rect 6134 4392 9586 4448
rect 9642 4392 9647 4448
rect 6134 4390 9647 4392
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 0 4254 1962 4314
rect 2129 4314 2195 4317
rect 4981 4314 5047 4317
rect 2129 4312 5047 4314
rect 2129 4256 2134 4312
rect 2190 4256 4986 4312
rect 5042 4256 5047 4312
rect 2129 4254 5047 4256
rect 0 4224 480 4254
rect 2129 4251 2195 4254
rect 4981 4251 5047 4254
rect 4337 4178 4403 4181
rect 6134 4178 6194 4390
rect 9581 4387 9647 4390
rect 17033 4450 17099 4453
rect 22832 4450 22892 4526
rect 26325 4523 26391 4526
rect 23473 4452 23539 4453
rect 17033 4448 22892 4450
rect 17033 4392 17038 4448
rect 17094 4392 22892 4448
rect 17033 4390 22892 4392
rect 17033 4387 17099 4390
rect 23422 4388 23428 4452
rect 23492 4450 23539 4452
rect 23492 4448 23584 4450
rect 23534 4392 23584 4448
rect 23492 4390 23584 4392
rect 23492 4388 23539 4390
rect 23473 4387 23539 4388
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 7005 4314 7071 4317
rect 7230 4314 7236 4316
rect 7005 4312 7236 4314
rect 7005 4256 7010 4312
rect 7066 4256 7236 4312
rect 7005 4254 7236 4256
rect 7005 4251 7071 4254
rect 7230 4252 7236 4254
rect 7300 4252 7306 4316
rect 9489 4314 9555 4317
rect 12525 4314 12591 4317
rect 9489 4312 12591 4314
rect 9489 4256 9494 4312
rect 9550 4256 12530 4312
rect 12586 4256 12591 4312
rect 9489 4254 12591 4256
rect 9489 4251 9555 4254
rect 12525 4251 12591 4254
rect 16389 4314 16455 4317
rect 17033 4314 17099 4317
rect 16389 4312 17099 4314
rect 16389 4256 16394 4312
rect 16450 4256 17038 4312
rect 17094 4256 17099 4312
rect 16389 4254 17099 4256
rect 16389 4251 16455 4254
rect 17033 4251 17099 4254
rect 21449 4314 21515 4317
rect 24117 4314 24183 4317
rect 21449 4312 24183 4314
rect 21449 4256 21454 4312
rect 21510 4256 24122 4312
rect 24178 4256 24183 4312
rect 21449 4254 24183 4256
rect 21449 4251 21515 4254
rect 24117 4251 24183 4254
rect 4337 4176 6194 4178
rect 4337 4120 4342 4176
rect 4398 4120 6194 4176
rect 4337 4118 6194 4120
rect 6361 4178 6427 4181
rect 17125 4178 17191 4181
rect 6361 4176 17191 4178
rect 6361 4120 6366 4176
rect 6422 4120 17130 4176
rect 17186 4120 17191 4176
rect 6361 4118 17191 4120
rect 4337 4115 4403 4118
rect 6361 4115 6427 4118
rect 17125 4115 17191 4118
rect 17309 4178 17375 4181
rect 21817 4178 21883 4181
rect 17309 4176 21883 4178
rect 17309 4120 17314 4176
rect 17370 4120 21822 4176
rect 21878 4120 21883 4176
rect 17309 4118 21883 4120
rect 17309 4115 17375 4118
rect 21817 4115 21883 4118
rect 22369 4178 22435 4181
rect 27520 4178 28000 4208
rect 22369 4176 28000 4178
rect 22369 4120 22374 4176
rect 22430 4120 28000 4176
rect 22369 4118 28000 4120
rect 22369 4115 22435 4118
rect 27520 4088 28000 4118
rect 1577 4042 1643 4045
rect 5993 4042 6059 4045
rect 1577 4040 6059 4042
rect 1577 3984 1582 4040
rect 1638 3984 5998 4040
rect 6054 3984 6059 4040
rect 1577 3982 6059 3984
rect 1577 3979 1643 3982
rect 5993 3979 6059 3982
rect 6310 3980 6316 4044
rect 6380 4042 6386 4044
rect 7005 4042 7071 4045
rect 6380 4040 7071 4042
rect 6380 3984 7010 4040
rect 7066 3984 7071 4040
rect 6380 3982 7071 3984
rect 6380 3980 6386 3982
rect 7005 3979 7071 3982
rect 8109 4042 8175 4045
rect 9029 4042 9095 4045
rect 8109 4040 9095 4042
rect 8109 3984 8114 4040
rect 8170 3984 9034 4040
rect 9090 3984 9095 4040
rect 8109 3982 9095 3984
rect 8109 3979 8175 3982
rect 9029 3979 9095 3982
rect 11094 3980 11100 4044
rect 11164 4042 11170 4044
rect 11789 4042 11855 4045
rect 11164 4040 11855 4042
rect 11164 3984 11794 4040
rect 11850 3984 11855 4040
rect 11164 3982 11855 3984
rect 11164 3980 11170 3982
rect 11789 3979 11855 3982
rect 12382 3980 12388 4044
rect 12452 4042 12458 4044
rect 20161 4042 20227 4045
rect 12452 4040 20227 4042
rect 12452 3984 20166 4040
rect 20222 3984 20227 4040
rect 12452 3982 20227 3984
rect 12452 3980 12458 3982
rect 20161 3979 20227 3982
rect 20529 4042 20595 4045
rect 22277 4042 22343 4045
rect 23749 4044 23815 4045
rect 23749 4042 23796 4044
rect 20529 4040 22343 4042
rect 20529 3984 20534 4040
rect 20590 3984 22282 4040
rect 22338 3984 22343 4040
rect 20529 3982 22343 3984
rect 23704 4040 23796 4042
rect 23704 3984 23754 4040
rect 23704 3982 23796 3984
rect 20529 3979 20595 3982
rect 22277 3979 22343 3982
rect 23749 3980 23796 3982
rect 23860 3980 23866 4044
rect 23933 4042 23999 4045
rect 24117 4042 24183 4045
rect 23933 4040 24183 4042
rect 23933 3984 23938 4040
rect 23994 3984 24122 4040
rect 24178 3984 24183 4040
rect 23933 3982 24183 3984
rect 23749 3979 23815 3980
rect 23933 3979 23999 3982
rect 24117 3979 24183 3982
rect 2865 3906 2931 3909
rect 5257 3906 5323 3909
rect 2865 3904 5323 3906
rect 2865 3848 2870 3904
rect 2926 3848 5262 3904
rect 5318 3848 5323 3904
rect 2865 3846 5323 3848
rect 2865 3843 2931 3846
rect 5257 3843 5323 3846
rect 6545 3906 6611 3909
rect 9990 3906 9996 3908
rect 6545 3904 9996 3906
rect 6545 3848 6550 3904
rect 6606 3848 9996 3904
rect 6545 3846 9996 3848
rect 6545 3843 6611 3846
rect 9990 3844 9996 3846
rect 10060 3844 10066 3908
rect 12893 3906 12959 3909
rect 15469 3906 15535 3909
rect 12893 3904 15535 3906
rect 12893 3848 12898 3904
rect 12954 3848 15474 3904
rect 15530 3848 15535 3904
rect 12893 3846 15535 3848
rect 12893 3843 12959 3846
rect 15469 3843 15535 3846
rect 16798 3844 16804 3908
rect 16868 3906 16874 3908
rect 17677 3906 17743 3909
rect 18229 3906 18295 3909
rect 16868 3904 18295 3906
rect 16868 3848 17682 3904
rect 17738 3848 18234 3904
rect 18290 3848 18295 3904
rect 16868 3846 18295 3848
rect 16868 3844 16874 3846
rect 17677 3843 17743 3846
rect 18229 3843 18295 3846
rect 20478 3844 20484 3908
rect 20548 3906 20554 3908
rect 20621 3906 20687 3909
rect 20897 3906 20963 3909
rect 20548 3904 20963 3906
rect 20548 3848 20626 3904
rect 20682 3848 20902 3904
rect 20958 3848 20963 3904
rect 20548 3846 20963 3848
rect 20548 3844 20554 3846
rect 20621 3843 20687 3846
rect 20897 3843 20963 3846
rect 22645 3906 22711 3909
rect 23933 3906 23999 3909
rect 22645 3904 23999 3906
rect 22645 3848 22650 3904
rect 22706 3848 23938 3904
rect 23994 3848 23999 3904
rect 22645 3846 23999 3848
rect 22645 3843 22711 3846
rect 23933 3843 23999 3846
rect 24577 3906 24643 3909
rect 26233 3906 26299 3909
rect 24577 3904 26299 3906
rect 24577 3848 24582 3904
rect 24638 3848 26238 3904
rect 26294 3848 26299 3904
rect 24577 3846 26299 3848
rect 24577 3843 24643 3846
rect 26233 3843 26299 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 3233 3770 3299 3773
rect 10041 3770 10107 3773
rect 13905 3770 13971 3773
rect 3233 3768 10107 3770
rect 3233 3712 3238 3768
rect 3294 3712 10046 3768
rect 10102 3712 10107 3768
rect 3233 3710 10107 3712
rect 3233 3707 3299 3710
rect 10041 3707 10107 3710
rect 11470 3768 13971 3770
rect 11470 3712 13910 3768
rect 13966 3712 13971 3768
rect 11470 3710 13971 3712
rect 0 3634 480 3664
rect 4429 3634 4495 3637
rect 0 3632 4495 3634
rect 0 3576 4434 3632
rect 4490 3576 4495 3632
rect 0 3574 4495 3576
rect 0 3544 480 3574
rect 4429 3571 4495 3574
rect 4889 3634 4955 3637
rect 6678 3634 6684 3636
rect 4889 3632 6684 3634
rect 4889 3576 4894 3632
rect 4950 3576 6684 3632
rect 4889 3574 6684 3576
rect 4889 3571 4955 3574
rect 6678 3572 6684 3574
rect 6748 3572 6754 3636
rect 7649 3634 7715 3637
rect 11470 3634 11530 3710
rect 13905 3707 13971 3710
rect 14181 3770 14247 3773
rect 15653 3770 15719 3773
rect 17125 3772 17191 3773
rect 17125 3770 17172 3772
rect 14181 3768 15719 3770
rect 14181 3712 14186 3768
rect 14242 3712 15658 3768
rect 15714 3712 15719 3768
rect 14181 3710 15719 3712
rect 17080 3768 17172 3770
rect 17236 3770 17242 3772
rect 19425 3770 19491 3773
rect 17236 3768 19491 3770
rect 17080 3712 17130 3768
rect 17236 3712 19430 3768
rect 19486 3712 19491 3768
rect 17080 3710 17172 3712
rect 14181 3707 14247 3710
rect 15653 3707 15719 3710
rect 17125 3708 17172 3710
rect 17236 3710 19491 3712
rect 17236 3708 17242 3710
rect 17125 3707 17191 3708
rect 19425 3707 19491 3710
rect 20805 3770 20871 3773
rect 21030 3770 21036 3772
rect 20805 3768 21036 3770
rect 20805 3712 20810 3768
rect 20866 3712 21036 3768
rect 20805 3710 21036 3712
rect 20805 3707 20871 3710
rect 21030 3708 21036 3710
rect 21100 3708 21106 3772
rect 21357 3770 21423 3773
rect 21357 3768 24962 3770
rect 21357 3712 21362 3768
rect 21418 3712 24962 3768
rect 21357 3710 24962 3712
rect 21357 3707 21423 3710
rect 7649 3632 11530 3634
rect 7649 3576 7654 3632
rect 7710 3576 11530 3632
rect 7649 3574 11530 3576
rect 11605 3634 11671 3637
rect 13813 3634 13879 3637
rect 11605 3632 13879 3634
rect 11605 3576 11610 3632
rect 11666 3576 13818 3632
rect 13874 3576 13879 3632
rect 11605 3574 13879 3576
rect 7649 3571 7715 3574
rect 11605 3571 11671 3574
rect 13813 3571 13879 3574
rect 14641 3634 14707 3637
rect 19333 3634 19399 3637
rect 14641 3632 19399 3634
rect 14641 3576 14646 3632
rect 14702 3576 19338 3632
rect 19394 3576 19399 3632
rect 14641 3574 19399 3576
rect 14641 3571 14707 3574
rect 19333 3571 19399 3574
rect 20161 3634 20227 3637
rect 22737 3634 22803 3637
rect 20161 3632 22803 3634
rect 20161 3576 20166 3632
rect 20222 3576 22742 3632
rect 22798 3576 22803 3632
rect 20161 3574 22803 3576
rect 20161 3571 20227 3574
rect 22737 3571 22803 3574
rect 24577 3634 24643 3637
rect 24710 3634 24716 3636
rect 24577 3632 24716 3634
rect 24577 3576 24582 3632
rect 24638 3576 24716 3632
rect 24577 3574 24716 3576
rect 24577 3571 24643 3574
rect 24710 3572 24716 3574
rect 24780 3572 24786 3636
rect 24902 3634 24962 3710
rect 27520 3634 28000 3664
rect 24902 3574 28000 3634
rect 27520 3544 28000 3574
rect 3417 3498 3483 3501
rect 9489 3498 9555 3501
rect 3417 3496 9555 3498
rect 3417 3440 3422 3496
rect 3478 3440 9494 3496
rect 9550 3440 9555 3496
rect 3417 3438 9555 3440
rect 3417 3435 3483 3438
rect 9489 3435 9555 3438
rect 9765 3498 9831 3501
rect 13629 3498 13695 3501
rect 13905 3500 13971 3501
rect 9765 3496 13695 3498
rect 9765 3440 9770 3496
rect 9826 3440 13634 3496
rect 13690 3440 13695 3496
rect 9765 3438 13695 3440
rect 9765 3435 9831 3438
rect 13629 3435 13695 3438
rect 13854 3436 13860 3500
rect 13924 3498 13971 3500
rect 14089 3498 14155 3501
rect 18137 3498 18203 3501
rect 13924 3496 14016 3498
rect 13966 3440 14016 3496
rect 13924 3438 14016 3440
rect 14089 3496 18203 3498
rect 14089 3440 14094 3496
rect 14150 3440 18142 3496
rect 18198 3440 18203 3496
rect 14089 3438 18203 3440
rect 13924 3436 13971 3438
rect 13905 3435 13971 3436
rect 14089 3435 14155 3438
rect 18137 3435 18203 3438
rect 18413 3498 18479 3501
rect 20253 3498 20319 3501
rect 18413 3496 20319 3498
rect 18413 3440 18418 3496
rect 18474 3440 20258 3496
rect 20314 3440 20319 3496
rect 18413 3438 20319 3440
rect 18413 3435 18479 3438
rect 20253 3435 20319 3438
rect 21173 3498 21239 3501
rect 25037 3498 25103 3501
rect 21173 3496 25103 3498
rect 21173 3440 21178 3496
rect 21234 3440 25042 3496
rect 25098 3440 25103 3496
rect 21173 3438 25103 3440
rect 21173 3435 21239 3438
rect 25037 3435 25103 3438
rect 7741 3362 7807 3365
rect 8017 3362 8083 3365
rect 10777 3362 10843 3365
rect 7741 3360 10843 3362
rect 7741 3304 7746 3360
rect 7802 3304 8022 3360
rect 8078 3304 10782 3360
rect 10838 3304 10843 3360
rect 7741 3302 10843 3304
rect 7741 3299 7807 3302
rect 8017 3299 8083 3302
rect 10777 3299 10843 3302
rect 16481 3362 16547 3365
rect 18597 3362 18663 3365
rect 16481 3360 18663 3362
rect 16481 3304 16486 3360
rect 16542 3304 18602 3360
rect 18658 3304 18663 3360
rect 16481 3302 18663 3304
rect 16481 3299 16547 3302
rect 18597 3299 18663 3302
rect 20345 3362 20411 3365
rect 22277 3362 22343 3365
rect 20345 3360 22343 3362
rect 20345 3304 20350 3360
rect 20406 3304 22282 3360
rect 22338 3304 22343 3360
rect 20345 3302 22343 3304
rect 20345 3299 20411 3302
rect 22277 3299 22343 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 16614 3164 16620 3228
rect 16684 3226 16690 3228
rect 16849 3226 16915 3229
rect 16684 3224 16915 3226
rect 16684 3168 16854 3224
rect 16910 3168 16915 3224
rect 16684 3166 16915 3168
rect 16684 3164 16690 3166
rect 16849 3163 16915 3166
rect 18689 3226 18755 3229
rect 22553 3226 22619 3229
rect 18689 3224 22619 3226
rect 18689 3168 18694 3224
rect 18750 3168 22558 3224
rect 22614 3168 22619 3224
rect 18689 3166 22619 3168
rect 18689 3163 18755 3166
rect 22553 3163 22619 3166
rect 24853 3226 24919 3229
rect 25262 3226 25268 3228
rect 24853 3224 25268 3226
rect 24853 3168 24858 3224
rect 24914 3168 25268 3224
rect 24853 3166 25268 3168
rect 24853 3163 24919 3166
rect 25262 3164 25268 3166
rect 25332 3226 25338 3228
rect 26325 3226 26391 3229
rect 25332 3224 26391 3226
rect 25332 3168 26330 3224
rect 26386 3168 26391 3224
rect 25332 3166 26391 3168
rect 25332 3164 25338 3166
rect 26325 3163 26391 3166
rect 5349 3090 5415 3093
rect 6913 3090 6979 3093
rect 12157 3090 12223 3093
rect 5349 3088 6979 3090
rect 5349 3032 5354 3088
rect 5410 3032 6918 3088
rect 6974 3032 6979 3088
rect 5349 3030 6979 3032
rect 5349 3027 5415 3030
rect 6913 3027 6979 3030
rect 9998 3088 12223 3090
rect 9998 3032 12162 3088
rect 12218 3032 12223 3088
rect 9998 3030 12223 3032
rect 0 2954 480 2984
rect 7649 2954 7715 2957
rect 0 2952 7715 2954
rect 0 2896 7654 2952
rect 7710 2896 7715 2952
rect 0 2894 7715 2896
rect 0 2864 480 2894
rect 7649 2891 7715 2894
rect 2497 2818 2563 2821
rect 9998 2818 10058 3030
rect 12157 3027 12223 3030
rect 20437 3090 20503 3093
rect 22829 3090 22895 3093
rect 20437 3088 22895 3090
rect 20437 3032 20442 3088
rect 20498 3032 22834 3088
rect 22890 3032 22895 3088
rect 20437 3030 22895 3032
rect 20437 3027 20503 3030
rect 22829 3027 22895 3030
rect 23381 3090 23447 3093
rect 25129 3090 25195 3093
rect 23381 3088 25195 3090
rect 23381 3032 23386 3088
rect 23442 3032 25134 3088
rect 25190 3032 25195 3088
rect 23381 3030 25195 3032
rect 23381 3027 23447 3030
rect 25129 3027 25195 3030
rect 26601 3090 26667 3093
rect 27520 3090 28000 3120
rect 26601 3088 28000 3090
rect 26601 3032 26606 3088
rect 26662 3032 28000 3088
rect 26601 3030 28000 3032
rect 26601 3027 26667 3030
rect 27520 3000 28000 3030
rect 10133 2954 10199 2957
rect 10726 2954 10732 2956
rect 10133 2952 10732 2954
rect 10133 2896 10138 2952
rect 10194 2896 10732 2952
rect 10133 2894 10732 2896
rect 10133 2891 10199 2894
rect 10726 2892 10732 2894
rect 10796 2892 10802 2956
rect 14549 2954 14615 2957
rect 22737 2954 22803 2957
rect 24117 2954 24183 2957
rect 25129 2954 25195 2957
rect 14549 2952 20178 2954
rect 14549 2896 14554 2952
rect 14610 2896 20178 2952
rect 14549 2894 20178 2896
rect 14549 2891 14615 2894
rect 2497 2816 10058 2818
rect 2497 2760 2502 2816
rect 2558 2760 10058 2816
rect 2497 2758 10058 2760
rect 10777 2818 10843 2821
rect 12382 2818 12388 2820
rect 10777 2816 12388 2818
rect 10777 2760 10782 2816
rect 10838 2760 12388 2816
rect 10777 2758 12388 2760
rect 2497 2755 2563 2758
rect 10777 2755 10843 2758
rect 12382 2756 12388 2758
rect 12452 2756 12458 2820
rect 12525 2818 12591 2821
rect 18689 2818 18755 2821
rect 12525 2816 18755 2818
rect 12525 2760 12530 2816
rect 12586 2760 18694 2816
rect 18750 2760 18755 2816
rect 12525 2758 18755 2760
rect 20118 2818 20178 2894
rect 22737 2952 25195 2954
rect 22737 2896 22742 2952
rect 22798 2896 24122 2952
rect 24178 2896 25134 2952
rect 25190 2896 25195 2952
rect 22737 2894 25195 2896
rect 22737 2891 22803 2894
rect 24117 2891 24183 2894
rect 25129 2891 25195 2894
rect 22461 2818 22527 2821
rect 20118 2816 22527 2818
rect 20118 2760 22466 2816
rect 22522 2760 22527 2816
rect 20118 2758 22527 2760
rect 12525 2755 12591 2758
rect 18689 2755 18755 2758
rect 22461 2755 22527 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 10685 2682 10751 2685
rect 16665 2682 16731 2685
rect 21725 2684 21791 2685
rect 21725 2682 21772 2684
rect 10685 2680 16731 2682
rect 10685 2624 10690 2680
rect 10746 2624 16670 2680
rect 16726 2624 16731 2680
rect 10685 2622 16731 2624
rect 21680 2680 21772 2682
rect 21680 2624 21730 2680
rect 21680 2622 21772 2624
rect 10685 2619 10751 2622
rect 16665 2619 16731 2622
rect 21725 2620 21772 2622
rect 21836 2620 21842 2684
rect 21725 2619 21791 2620
rect 3417 2546 3483 2549
rect 7373 2546 7439 2549
rect 3417 2544 7439 2546
rect 3417 2488 3422 2544
rect 3478 2488 7378 2544
rect 7434 2488 7439 2544
rect 3417 2486 7439 2488
rect 3417 2483 3483 2486
rect 7373 2483 7439 2486
rect 10317 2546 10383 2549
rect 12433 2546 12499 2549
rect 10317 2544 12499 2546
rect 10317 2488 10322 2544
rect 10378 2488 12438 2544
rect 12494 2488 12499 2544
rect 10317 2486 12499 2488
rect 10317 2483 10383 2486
rect 12433 2483 12499 2486
rect 16573 2546 16639 2549
rect 23657 2546 23723 2549
rect 16573 2544 23723 2546
rect 16573 2488 16578 2544
rect 16634 2488 23662 2544
rect 23718 2488 23723 2544
rect 16573 2486 23723 2488
rect 16573 2483 16639 2486
rect 23657 2483 23723 2486
rect 26509 2546 26575 2549
rect 27520 2546 28000 2576
rect 26509 2544 28000 2546
rect 26509 2488 26514 2544
rect 26570 2488 28000 2544
rect 26509 2486 28000 2488
rect 26509 2483 26575 2486
rect 27520 2456 28000 2486
rect 2957 2410 3023 2413
rect 3918 2410 3924 2412
rect 2957 2408 3924 2410
rect 2957 2352 2962 2408
rect 3018 2352 3924 2408
rect 2957 2350 3924 2352
rect 2957 2347 3023 2350
rect 3918 2348 3924 2350
rect 3988 2348 3994 2412
rect 5901 2410 5967 2413
rect 18873 2410 18939 2413
rect 21357 2410 21423 2413
rect 25405 2410 25471 2413
rect 5901 2408 17970 2410
rect 5901 2352 5906 2408
rect 5962 2352 17970 2408
rect 5901 2350 17970 2352
rect 5901 2347 5967 2350
rect 0 2274 480 2304
rect 3693 2274 3759 2277
rect 0 2272 3759 2274
rect 0 2216 3698 2272
rect 3754 2216 3759 2272
rect 0 2214 3759 2216
rect 0 2184 480 2214
rect 3693 2211 3759 2214
rect 7465 2274 7531 2277
rect 10501 2274 10567 2277
rect 7465 2272 10567 2274
rect 7465 2216 7470 2272
rect 7526 2216 10506 2272
rect 10562 2216 10567 2272
rect 7465 2214 10567 2216
rect 7465 2211 7531 2214
rect 10501 2211 10567 2214
rect 10685 2274 10751 2277
rect 13261 2274 13327 2277
rect 17910 2274 17970 2350
rect 18873 2408 25471 2410
rect 18873 2352 18878 2408
rect 18934 2352 21362 2408
rect 21418 2352 25410 2408
rect 25466 2352 25471 2408
rect 18873 2350 25471 2352
rect 18873 2347 18939 2350
rect 21357 2347 21423 2350
rect 25405 2347 25471 2350
rect 19149 2274 19215 2277
rect 10685 2272 13327 2274
rect 10685 2216 10690 2272
rect 10746 2216 13266 2272
rect 13322 2216 13327 2272
rect 10685 2214 13327 2216
rect 10685 2211 10751 2214
rect 13261 2211 13327 2214
rect 15334 2214 17786 2274
rect 17910 2272 19215 2274
rect 17910 2216 19154 2272
rect 19210 2216 19215 2272
rect 17910 2214 19215 2216
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 7557 2138 7623 2141
rect 14641 2138 14707 2141
rect 7557 2136 14707 2138
rect 7557 2080 7562 2136
rect 7618 2080 14646 2136
rect 14702 2080 14707 2136
rect 7557 2078 14707 2080
rect 7557 2075 7623 2078
rect 14641 2075 14707 2078
rect 3141 2002 3207 2005
rect 11145 2002 11211 2005
rect 3141 2000 11211 2002
rect 3141 1944 3146 2000
rect 3202 1944 11150 2000
rect 11206 1944 11211 2000
rect 3141 1942 11211 1944
rect 3141 1939 3207 1942
rect 11145 1939 11211 1942
rect 11329 2002 11395 2005
rect 15334 2002 15394 2214
rect 17401 2138 17467 2141
rect 11329 2000 15394 2002
rect 11329 1944 11334 2000
rect 11390 1944 15394 2000
rect 11329 1942 15394 1944
rect 15518 2136 17467 2138
rect 15518 2080 17406 2136
rect 17462 2080 17467 2136
rect 15518 2078 17467 2080
rect 17726 2138 17786 2214
rect 19149 2211 19215 2214
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 24117 2138 24183 2141
rect 17726 2136 24183 2138
rect 17726 2080 24122 2136
rect 24178 2080 24183 2136
rect 17726 2078 24183 2080
rect 11329 1939 11395 1942
rect 8937 1866 9003 1869
rect 15518 1866 15578 2078
rect 17401 2075 17467 2078
rect 24117 2075 24183 2078
rect 15745 2002 15811 2005
rect 25497 2002 25563 2005
rect 15745 2000 25563 2002
rect 15745 1944 15750 2000
rect 15806 1944 25502 2000
rect 25558 1944 25563 2000
rect 15745 1942 25563 1944
rect 15745 1939 15811 1942
rect 25497 1939 25563 1942
rect 25957 2002 26023 2005
rect 27520 2002 28000 2032
rect 25957 2000 28000 2002
rect 25957 1944 25962 2000
rect 26018 1944 28000 2000
rect 25957 1942 28000 1944
rect 25957 1939 26023 1942
rect 27520 1912 28000 1942
rect 8937 1864 15578 1866
rect 8937 1808 8942 1864
rect 8998 1808 15578 1864
rect 8937 1806 15578 1808
rect 15653 1866 15719 1869
rect 18413 1866 18479 1869
rect 15653 1864 18479 1866
rect 15653 1808 15658 1864
rect 15714 1808 18418 1864
rect 18474 1808 18479 1864
rect 15653 1806 18479 1808
rect 8937 1803 9003 1806
rect 15653 1803 15719 1806
rect 18413 1803 18479 1806
rect 18965 1866 19031 1869
rect 26417 1866 26483 1869
rect 18965 1864 26483 1866
rect 18965 1808 18970 1864
rect 19026 1808 26422 1864
rect 26478 1808 26483 1864
rect 18965 1806 26483 1808
rect 18965 1803 19031 1806
rect 26417 1803 26483 1806
rect 7925 1730 7991 1733
rect 14549 1730 14615 1733
rect 7925 1728 14615 1730
rect 7925 1672 7930 1728
rect 7986 1672 14554 1728
rect 14610 1672 14615 1728
rect 7925 1670 14615 1672
rect 7925 1667 7991 1670
rect 14549 1667 14615 1670
rect 14733 1730 14799 1733
rect 22369 1730 22435 1733
rect 14733 1728 22435 1730
rect 14733 1672 14738 1728
rect 14794 1672 22374 1728
rect 22430 1672 22435 1728
rect 14733 1670 22435 1672
rect 14733 1667 14799 1670
rect 22369 1667 22435 1670
rect 0 1594 480 1624
rect 2998 1594 3004 1596
rect 0 1534 3004 1594
rect 0 1504 480 1534
rect 2998 1532 3004 1534
rect 3068 1532 3074 1596
rect 3785 1594 3851 1597
rect 4429 1594 4495 1597
rect 13629 1594 13695 1597
rect 3785 1592 13695 1594
rect 3785 1536 3790 1592
rect 3846 1536 4434 1592
rect 4490 1536 13634 1592
rect 13690 1536 13695 1592
rect 3785 1534 13695 1536
rect 3785 1531 3851 1534
rect 4429 1531 4495 1534
rect 13629 1531 13695 1534
rect 14457 1594 14523 1597
rect 25589 1594 25655 1597
rect 14457 1592 25655 1594
rect 14457 1536 14462 1592
rect 14518 1536 25594 1592
rect 25650 1536 25655 1592
rect 14457 1534 25655 1536
rect 14457 1531 14523 1534
rect 25589 1531 25655 1534
rect 7782 1458 7788 1460
rect 1948 1398 7788 1458
rect 0 914 480 944
rect 1948 914 2008 1398
rect 7782 1396 7788 1398
rect 7852 1396 7858 1460
rect 12893 1458 12959 1461
rect 14917 1458 14983 1461
rect 12893 1456 14983 1458
rect 12893 1400 12898 1456
rect 12954 1400 14922 1456
rect 14978 1400 14983 1456
rect 12893 1398 14983 1400
rect 12893 1395 12959 1398
rect 14917 1395 14983 1398
rect 15101 1458 15167 1461
rect 19333 1458 19399 1461
rect 15101 1456 19399 1458
rect 15101 1400 15106 1456
rect 15162 1400 19338 1456
rect 19394 1400 19399 1456
rect 15101 1398 19399 1400
rect 15101 1395 15167 1398
rect 19333 1395 19399 1398
rect 20161 1458 20227 1461
rect 24945 1458 25011 1461
rect 20161 1456 25011 1458
rect 20161 1400 20166 1456
rect 20222 1400 24950 1456
rect 25006 1400 25011 1456
rect 20161 1398 25011 1400
rect 20161 1395 20227 1398
rect 24945 1395 25011 1398
rect 25681 1458 25747 1461
rect 27520 1458 28000 1488
rect 25681 1456 28000 1458
rect 25681 1400 25686 1456
rect 25742 1400 28000 1456
rect 25681 1398 28000 1400
rect 25681 1395 25747 1398
rect 27520 1368 28000 1398
rect 2129 1322 2195 1325
rect 17493 1322 17559 1325
rect 2129 1320 17559 1322
rect 2129 1264 2134 1320
rect 2190 1264 17498 1320
rect 17554 1264 17559 1320
rect 2129 1262 17559 1264
rect 2129 1259 2195 1262
rect 17493 1259 17559 1262
rect 17861 1322 17927 1325
rect 24669 1322 24735 1325
rect 17861 1320 24735 1322
rect 17861 1264 17866 1320
rect 17922 1264 24674 1320
rect 24730 1264 24735 1320
rect 17861 1262 24735 1264
rect 17861 1259 17927 1262
rect 24669 1259 24735 1262
rect 2814 1124 2820 1188
rect 2884 1186 2890 1188
rect 15285 1186 15351 1189
rect 2884 1184 15351 1186
rect 2884 1128 15290 1184
rect 15346 1128 15351 1184
rect 2884 1126 15351 1128
rect 2884 1124 2890 1126
rect 15285 1123 15351 1126
rect 22921 1186 22987 1189
rect 25313 1186 25379 1189
rect 22921 1184 25379 1186
rect 22921 1128 22926 1184
rect 22982 1128 25318 1184
rect 25374 1128 25379 1184
rect 22921 1126 25379 1128
rect 22921 1123 22987 1126
rect 25313 1123 25379 1126
rect 3693 1050 3759 1053
rect 20069 1050 20135 1053
rect 3693 1048 20135 1050
rect 3693 992 3698 1048
rect 3754 992 20074 1048
rect 20130 992 20135 1048
rect 3693 990 20135 992
rect 3693 987 3759 990
rect 20069 987 20135 990
rect 20478 988 20484 1052
rect 20548 1050 20554 1052
rect 23197 1050 23263 1053
rect 20548 1048 23263 1050
rect 20548 992 23202 1048
rect 23258 992 23263 1048
rect 20548 990 23263 992
rect 20548 988 20554 990
rect 23197 987 23263 990
rect 0 854 2008 914
rect 7373 914 7439 917
rect 20621 914 20687 917
rect 7373 912 20687 914
rect 7373 856 7378 912
rect 7434 856 20626 912
rect 20682 856 20687 912
rect 7373 854 20687 856
rect 0 824 480 854
rect 7373 851 7439 854
rect 20621 851 20687 854
rect 23289 914 23355 917
rect 27520 914 28000 944
rect 23289 912 28000 914
rect 23289 856 23294 912
rect 23350 856 28000 912
rect 23289 854 28000 856
rect 23289 851 23355 854
rect 27520 824 28000 854
rect 1393 778 1459 781
rect 23013 778 23079 781
rect 1393 776 23079 778
rect 1393 720 1398 776
rect 1454 720 23018 776
rect 23074 720 23079 776
rect 1393 718 23079 720
rect 1393 715 1459 718
rect 23013 715 23079 718
rect 7046 580 7052 644
rect 7116 642 7122 644
rect 27061 642 27127 645
rect 7116 640 27127 642
rect 7116 584 27066 640
rect 27122 584 27127 640
rect 7116 582 27127 584
rect 7116 580 7122 582
rect 27061 579 27127 582
rect 16389 506 16455 509
rect 22921 506 22987 509
rect 16389 504 22987 506
rect 16389 448 16394 504
rect 16450 448 22926 504
rect 22982 448 22987 504
rect 16389 446 22987 448
rect 16389 443 16455 446
rect 22921 443 22987 446
rect 0 370 480 400
rect 4429 370 4495 373
rect 0 368 4495 370
rect 0 312 4434 368
rect 4490 312 4495 368
rect 0 310 4495 312
rect 0 280 480 310
rect 4429 307 4495 310
rect 15561 370 15627 373
rect 26417 370 26483 373
rect 15561 368 26483 370
rect 15561 312 15566 368
rect 15622 312 26422 368
rect 26478 312 26483 368
rect 15561 310 26483 312
rect 15561 307 15627 310
rect 26417 307 26483 310
rect 26693 370 26759 373
rect 27520 370 28000 400
rect 26693 368 28000 370
rect 26693 312 26698 368
rect 26754 312 28000 368
rect 26693 310 28000 312
rect 26693 307 26759 310
rect 27520 280 28000 310
rect 13721 234 13787 237
rect 27337 234 27403 237
rect 13721 232 27403 234
rect 13721 176 13726 232
rect 13782 176 27342 232
rect 27398 176 27403 232
rect 13721 174 27403 176
rect 13721 171 13787 174
rect 27337 171 27403 174
rect 3969 98 4035 101
rect 20897 98 20963 101
rect 3969 96 20963 98
rect 3969 40 3974 96
rect 4030 40 20902 96
rect 20958 40 20963 96
rect 3969 38 20963 40
rect 3969 35 4035 38
rect 20897 35 20963 38
<< via3 >>
rect 3372 27644 3436 27708
rect 26372 26148 26436 26212
rect 20668 25876 20732 25940
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 5396 25468 5460 25532
rect 26924 25604 26988 25668
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 6316 25196 6380 25260
rect 21036 25196 21100 25260
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 3004 24848 3068 24852
rect 3004 24792 3054 24848
rect 3054 24792 3068 24848
rect 3004 24788 3068 24792
rect 3188 24788 3252 24852
rect 9812 24848 9876 24852
rect 9812 24792 9826 24848
rect 9826 24792 9876 24848
rect 9812 24788 9876 24792
rect 8708 24516 8772 24580
rect 20300 24516 20364 24580
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 9444 24244 9508 24308
rect 8156 23972 8220 24036
rect 22324 24108 22388 24172
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 20852 23896 20916 23900
rect 20852 23840 20866 23896
rect 20866 23840 20916 23896
rect 20852 23836 20916 23840
rect 21956 23836 22020 23900
rect 5028 23428 5092 23492
rect 9996 23428 10060 23492
rect 20484 23564 20548 23628
rect 16620 23428 16684 23492
rect 18644 23488 18708 23492
rect 18644 23432 18658 23488
rect 18658 23432 18708 23488
rect 18644 23428 18708 23432
rect 20116 23488 20180 23492
rect 20116 23432 20130 23488
rect 20130 23432 20180 23488
rect 20116 23428 20180 23432
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 6132 23292 6196 23356
rect 9076 23156 9140 23220
rect 23060 23428 23124 23492
rect 23796 23488 23860 23492
rect 23796 23432 23810 23488
rect 23810 23432 23860 23488
rect 23796 23428 23860 23432
rect 24716 23428 24780 23492
rect 21588 23292 21652 23356
rect 11652 23020 11716 23084
rect 23980 23020 24044 23084
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 9444 22748 9508 22812
rect 9582 22748 9646 22812
rect 8340 22612 8404 22676
rect 3924 22476 3988 22540
rect 6132 22340 6196 22404
rect 6500 22400 6564 22404
rect 6500 22344 6550 22400
rect 6550 22344 6564 22400
rect 6500 22340 6564 22344
rect 7972 22340 8036 22404
rect 8708 22400 8772 22404
rect 8708 22344 8722 22400
rect 8722 22344 8772 22400
rect 8708 22340 8772 22344
rect 4844 22204 4908 22268
rect 20668 22340 20732 22404
rect 21772 22340 21836 22404
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 8156 22068 8220 22132
rect 8708 22068 8772 22132
rect 20852 22128 20916 22132
rect 20852 22072 20866 22128
rect 20866 22072 20916 22128
rect 20852 22068 20916 22072
rect 22692 22068 22756 22132
rect 9996 21932 10060 21996
rect 18092 21932 18156 21996
rect 5396 21796 5460 21860
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 4476 21584 4540 21588
rect 8708 21660 8772 21724
rect 20668 21660 20732 21724
rect 21036 21660 21100 21724
rect 22876 21660 22940 21724
rect 25268 21660 25332 21724
rect 4476 21528 4526 21584
rect 4526 21528 4540 21584
rect 4476 21524 4540 21528
rect 21404 21524 21468 21588
rect 4660 21388 4724 21452
rect 6684 21252 6748 21316
rect 3924 21116 3988 21180
rect 7420 21116 7484 21180
rect 21036 21388 21100 21452
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 3740 20768 3804 20772
rect 3740 20712 3754 20768
rect 3754 20712 3804 20768
rect 3740 20708 3804 20712
rect 21404 20980 21468 21044
rect 15516 20708 15580 20772
rect 18092 20708 18156 20772
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 11652 20572 11716 20636
rect 8340 20436 8404 20500
rect 13308 20300 13372 20364
rect 20852 20360 20916 20364
rect 20852 20304 20902 20360
rect 20902 20304 20916 20360
rect 20852 20300 20916 20304
rect 8156 20164 8220 20228
rect 9628 20224 9692 20228
rect 9628 20168 9678 20224
rect 9678 20168 9692 20224
rect 9628 20164 9692 20168
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 2636 20028 2700 20092
rect 3188 20028 3252 20092
rect 9996 20088 10060 20092
rect 9996 20032 10010 20088
rect 10010 20032 10060 20088
rect 9996 20028 10060 20032
rect 10916 20028 10980 20092
rect 17172 20028 17236 20092
rect 21220 20164 21284 20228
rect 23428 20088 23492 20092
rect 23428 20032 23478 20088
rect 23478 20032 23492 20088
rect 23428 20028 23492 20032
rect 5396 19756 5460 19820
rect 9996 19756 10060 19820
rect 6316 19620 6380 19684
rect 12020 19620 12084 19684
rect 26004 19816 26068 19820
rect 26004 19760 26018 19816
rect 26018 19760 26068 19816
rect 26004 19756 26068 19760
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 11100 19484 11164 19548
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 22324 19484 22388 19548
rect 4292 19212 4356 19276
rect 7052 19272 7116 19276
rect 7052 19216 7066 19272
rect 7066 19216 7116 19272
rect 7052 19212 7116 19216
rect 23428 19212 23492 19276
rect 11836 19076 11900 19140
rect 12204 19076 12268 19140
rect 24900 19076 24964 19140
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5212 18940 5276 19004
rect 11652 18940 11716 19004
rect 20484 18940 20548 19004
rect 21220 18940 21284 19004
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 14596 18396 14660 18460
rect 3188 18184 3252 18188
rect 3188 18128 3238 18184
rect 3238 18128 3252 18184
rect 3188 18124 3252 18128
rect 3556 18124 3620 18188
rect 2268 18048 2332 18052
rect 2268 17992 2282 18048
rect 2282 17992 2332 18048
rect 2268 17988 2332 17992
rect 2820 18048 2884 18052
rect 2820 17992 2834 18048
rect 2834 17992 2884 18048
rect 2820 17988 2884 17992
rect 5028 17988 5092 18052
rect 9812 18124 9876 18188
rect 7052 17988 7116 18052
rect 16252 18048 16316 18052
rect 16252 17992 16266 18048
rect 16266 17992 16316 18048
rect 16252 17988 16316 17992
rect 21404 17988 21468 18052
rect 21772 17988 21836 18052
rect 22140 17988 22204 18052
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 2636 17912 2700 17916
rect 2636 17856 2650 17912
rect 2650 17856 2700 17912
rect 2636 17852 2700 17856
rect 6316 17852 6380 17916
rect 7788 17852 7852 17916
rect 8524 17852 8588 17916
rect 4844 17716 4908 17780
rect 20668 17852 20732 17916
rect 16620 17580 16684 17644
rect 14044 17444 14108 17508
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 10732 17308 10796 17372
rect 11468 17308 11532 17372
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 19012 17308 19076 17372
rect 10732 16900 10796 16964
rect 19380 17036 19444 17100
rect 20300 17036 20364 17100
rect 21772 17036 21836 17100
rect 23612 17096 23676 17100
rect 23612 17040 23626 17096
rect 23626 17040 23676 17096
rect 23612 17036 23676 17040
rect 24716 17036 24780 17100
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 1900 16628 1964 16692
rect 9812 16628 9876 16692
rect 11284 16628 11348 16692
rect 22324 16628 22388 16692
rect 4476 16492 4540 16556
rect 10732 16356 10796 16420
rect 10916 16356 10980 16420
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 8156 16220 8220 16284
rect 20668 16084 20732 16148
rect 10732 15812 10796 15876
rect 21404 15812 21468 15876
rect 21956 15812 22020 15876
rect 23980 15872 24044 15876
rect 23980 15816 24030 15872
rect 24030 15816 24044 15872
rect 23980 15812 24044 15816
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 4844 15676 4908 15740
rect 5396 15676 5460 15740
rect 9628 15736 9692 15740
rect 9628 15680 9642 15736
rect 9642 15680 9692 15736
rect 9628 15676 9692 15680
rect 22876 15540 22940 15604
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 20668 14996 20732 15060
rect 6316 14860 6380 14924
rect 6500 14860 6564 14924
rect 6868 14860 6932 14924
rect 4476 14724 4540 14788
rect 4292 14648 4356 14652
rect 4292 14592 4342 14648
rect 4342 14592 4356 14648
rect 4292 14588 4356 14592
rect 5212 14588 5276 14652
rect 22324 14860 22388 14924
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 8524 14512 8588 14516
rect 8524 14456 8574 14512
rect 8574 14456 8588 14512
rect 8524 14452 8588 14456
rect 16620 14452 16684 14516
rect 22140 14588 22204 14652
rect 23612 14588 23676 14652
rect 20300 14316 20364 14380
rect 22140 14180 22204 14244
rect 25084 14180 25148 14244
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 7052 13636 7116 13700
rect 16620 13908 16684 13972
rect 20300 13908 20364 13972
rect 20852 13908 20916 13972
rect 20116 13636 20180 13700
rect 20668 13636 20732 13700
rect 21036 13636 21100 13700
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 4844 13500 4908 13564
rect 5396 13500 5460 13564
rect 6316 13500 6380 13564
rect 19380 13500 19444 13564
rect 22508 13560 22572 13564
rect 22508 13504 22558 13560
rect 22558 13504 22572 13560
rect 22508 13500 22572 13504
rect 23428 13500 23492 13564
rect 24716 13500 24780 13564
rect 3924 13092 3988 13156
rect 5028 13092 5092 13156
rect 6684 13092 6748 13156
rect 7604 13092 7668 13156
rect 14044 13092 14108 13156
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 7052 12956 7116 13020
rect 7972 12956 8036 13020
rect 26004 13560 26068 13564
rect 26004 13504 26018 13560
rect 26018 13504 26068 13560
rect 26004 13500 26068 13504
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 19380 12880 19444 12884
rect 19380 12824 19394 12880
rect 19394 12824 19444 12880
rect 19380 12820 19444 12824
rect 3372 12608 3436 12612
rect 3372 12552 3386 12608
rect 3386 12552 3436 12608
rect 3372 12548 3436 12552
rect 11100 12548 11164 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 7972 12412 8036 12476
rect 8892 12412 8956 12476
rect 14596 12412 14660 12476
rect 23428 12548 23492 12612
rect 3556 12276 3620 12340
rect 8156 12276 8220 12340
rect 9444 12276 9508 12340
rect 12388 12276 12452 12340
rect 21036 12276 21100 12340
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 5028 11868 5092 11932
rect 6132 11868 6196 11932
rect 6500 11868 6564 11932
rect 4660 11732 4724 11796
rect 6132 11732 6196 11796
rect 21220 11928 21284 11932
rect 21220 11872 21270 11928
rect 21270 11872 21284 11928
rect 21220 11868 21284 11872
rect 24900 11928 24964 11932
rect 24900 11872 24914 11928
rect 24914 11872 24964 11928
rect 24900 11868 24964 11872
rect 21036 11732 21100 11796
rect 8892 11520 8956 11524
rect 8892 11464 8906 11520
rect 8906 11464 8956 11520
rect 8892 11460 8956 11464
rect 10732 11520 10796 11524
rect 10732 11464 10782 11520
rect 10782 11464 10796 11520
rect 10732 11460 10796 11464
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 12388 11324 12452 11388
rect 20300 11324 20364 11388
rect 24900 11324 24964 11388
rect 7052 10916 7116 10980
rect 15516 10976 15580 10980
rect 15516 10920 15530 10976
rect 15530 10920 15580 10976
rect 15516 10916 15580 10920
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 8524 10780 8588 10844
rect 14596 10840 14660 10844
rect 14596 10784 14646 10840
rect 14646 10784 14660 10840
rect 14596 10780 14660 10784
rect 22324 10780 22388 10844
rect 23980 10780 24044 10844
rect 2636 10644 2700 10708
rect 11284 10432 11348 10436
rect 20116 10644 20180 10708
rect 20484 10644 20548 10708
rect 11284 10376 11334 10432
rect 11334 10376 11348 10432
rect 11284 10372 11348 10376
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5396 10236 5460 10300
rect 9996 10236 10060 10300
rect 22140 10296 22204 10300
rect 22140 10240 22154 10296
rect 22154 10240 22204 10296
rect 22140 10236 22204 10240
rect 22324 10296 22388 10300
rect 22324 10240 22374 10296
rect 22374 10240 22388 10296
rect 22324 10236 22388 10240
rect 21404 9828 21468 9892
rect 22324 9828 22388 9892
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 23060 9828 23124 9892
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 9996 9284 10060 9348
rect 23980 9420 24044 9484
rect 24716 9420 24780 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 3004 9012 3068 9076
rect 4108 9012 4172 9076
rect 6684 9012 6748 9076
rect 5396 8876 5460 8940
rect 13860 8936 13924 8940
rect 13860 8880 13910 8936
rect 13910 8880 13924 8936
rect 13860 8876 13924 8880
rect 7052 8740 7116 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 25084 8604 25148 8668
rect 16804 8468 16868 8532
rect 3924 8196 3988 8260
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19012 8332 19076 8396
rect 11100 8234 11150 8260
rect 11150 8234 11164 8260
rect 11100 8196 11164 8234
rect 21220 8332 21284 8396
rect 22508 8332 22572 8396
rect 21588 8196 21652 8260
rect 23612 8196 23676 8260
rect 24716 8196 24780 8260
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 10732 7848 10796 7852
rect 10732 7792 10782 7848
rect 10782 7792 10796 7848
rect 10732 7788 10796 7792
rect 23980 7788 24044 7852
rect 14228 7652 14292 7716
rect 20484 7652 20548 7716
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 6132 7516 6196 7580
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 23428 7380 23492 7444
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 10732 6836 10796 6900
rect 20116 6972 20180 7036
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 8156 6700 8220 6764
rect 12204 6700 12268 6764
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 23980 6156 24044 6220
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5396 5748 5460 5812
rect 3188 5612 3252 5676
rect 10916 5612 10980 5676
rect 9444 5476 9508 5540
rect 9996 5476 10060 5540
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 13124 5340 13188 5404
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 24900 5340 24964 5404
rect 20852 5068 20916 5132
rect 21404 5068 21468 5132
rect 22140 5068 22204 5132
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 3556 4796 3620 4860
rect 6500 4796 6564 4860
rect 14596 4796 14660 4860
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 23428 4448 23492 4452
rect 23428 4392 23478 4448
rect 23478 4392 23492 4448
rect 23428 4388 23492 4392
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 7236 4252 7300 4316
rect 6316 3980 6380 4044
rect 11100 3980 11164 4044
rect 12388 3980 12452 4044
rect 23796 4040 23860 4044
rect 23796 3984 23810 4040
rect 23810 3984 23860 4040
rect 23796 3980 23860 3984
rect 9996 3844 10060 3908
rect 16804 3844 16868 3908
rect 20484 3844 20548 3908
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 6684 3572 6748 3636
rect 17172 3768 17236 3772
rect 17172 3712 17186 3768
rect 17186 3712 17236 3768
rect 17172 3708 17236 3712
rect 21036 3708 21100 3772
rect 24716 3572 24780 3636
rect 13860 3496 13924 3500
rect 13860 3440 13910 3496
rect 13910 3440 13924 3496
rect 13860 3436 13924 3440
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 16620 3164 16684 3228
rect 25268 3164 25332 3228
rect 10732 2892 10796 2956
rect 12388 2756 12452 2820
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 21772 2680 21836 2684
rect 21772 2624 21786 2680
rect 21786 2624 21836 2680
rect 21772 2620 21836 2624
rect 3924 2348 3988 2412
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 3004 1532 3068 1596
rect 7788 1396 7852 1460
rect 2820 1124 2884 1188
rect 20484 988 20548 1052
rect 7052 580 7116 644
<< metal4 >>
rect 3371 27708 3437 27709
rect 3371 27644 3372 27708
rect 3436 27644 3437 27708
rect 3371 27643 3437 27644
rect 3003 24852 3069 24853
rect 3003 24788 3004 24852
rect 3068 24788 3069 24852
rect 3003 24787 3069 24788
rect 3187 24852 3253 24853
rect 3187 24788 3188 24852
rect 3252 24788 3253 24852
rect 3187 24787 3253 24788
rect 2267 18052 2333 18053
rect 2267 17988 2268 18052
rect 2332 17988 2333 18052
rect 2267 17987 2333 17988
rect 2819 18052 2885 18053
rect 2819 17988 2820 18052
rect 2884 17988 2885 18052
rect 2819 17987 2885 17988
rect 2270 1818 2330 17987
rect 2635 17916 2701 17917
rect 2635 17852 2636 17916
rect 2700 17852 2701 17916
rect 2635 17851 2701 17852
rect 2638 10709 2698 17851
rect 2635 10708 2701 10709
rect 2635 10644 2636 10708
rect 2700 10644 2701 10708
rect 2635 10643 2701 10644
rect 2822 1189 2882 17987
rect 3006 9077 3066 24787
rect 3190 20093 3250 24787
rect 3187 20092 3253 20093
rect 3187 20028 3188 20092
rect 3252 20028 3253 20092
rect 3187 20027 3253 20028
rect 3187 18188 3253 18189
rect 3187 18124 3188 18188
rect 3252 18124 3253 18188
rect 3187 18123 3253 18124
rect 3003 9076 3069 9077
rect 3003 9012 3004 9076
rect 3068 9012 3069 9076
rect 3003 9011 3069 9012
rect 3190 5810 3250 18123
rect 3374 12613 3434 27643
rect 5395 25532 5461 25533
rect 5395 25468 5396 25532
rect 5460 25468 5461 25532
rect 5395 25467 5461 25468
rect 5027 23492 5093 23493
rect 5027 23428 5028 23492
rect 5092 23428 5093 23492
rect 5027 23427 5093 23428
rect 3923 22540 3989 22541
rect 3923 22476 3924 22540
rect 3988 22476 3989 22540
rect 3923 22475 3989 22476
rect 3926 21450 3986 22475
rect 4843 22268 4909 22269
rect 4843 22204 4844 22268
rect 4908 22204 4909 22268
rect 4843 22203 4909 22204
rect 4475 21588 4541 21589
rect 4475 21524 4476 21588
rect 4540 21524 4541 21588
rect 4475 21523 4541 21524
rect 3558 21390 3986 21450
rect 3558 18189 3618 21390
rect 3923 21180 3989 21181
rect 3923 21116 3924 21180
rect 3988 21116 3989 21180
rect 3923 21115 3989 21116
rect 3739 20772 3805 20773
rect 3739 20708 3740 20772
rect 3804 20708 3805 20772
rect 3739 20707 3805 20708
rect 3555 18188 3621 18189
rect 3555 18124 3556 18188
rect 3620 18124 3621 18188
rect 3555 18123 3621 18124
rect 3371 12612 3437 12613
rect 3371 12548 3372 12612
rect 3436 12548 3437 12612
rect 3371 12547 3437 12548
rect 3558 12341 3618 18123
rect 3555 12340 3621 12341
rect 3555 12276 3556 12340
rect 3620 12276 3621 12340
rect 3555 12275 3621 12276
rect 3742 8530 3802 20707
rect 3926 13157 3986 21115
rect 4291 19276 4357 19277
rect 4291 19212 4292 19276
rect 4356 19212 4357 19276
rect 4291 19211 4357 19212
rect 4294 14653 4354 19211
rect 4478 16557 4538 21523
rect 4659 21452 4725 21453
rect 4659 21388 4660 21452
rect 4724 21388 4725 21452
rect 4659 21387 4725 21388
rect 4475 16556 4541 16557
rect 4475 16492 4476 16556
rect 4540 16492 4541 16556
rect 4475 16491 4541 16492
rect 4478 14789 4538 16491
rect 4475 14788 4541 14789
rect 4475 14724 4476 14788
rect 4540 14724 4541 14788
rect 4475 14723 4541 14724
rect 4291 14652 4357 14653
rect 4291 14588 4292 14652
rect 4356 14588 4357 14652
rect 4291 14587 4357 14588
rect 3923 13156 3989 13157
rect 3923 13092 3924 13156
rect 3988 13092 3989 13156
rect 3923 13091 3989 13092
rect 4662 11797 4722 21387
rect 4846 17781 4906 22203
rect 5030 18053 5090 23427
rect 5398 21861 5458 25467
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 6134 23357 6194 26062
rect 20667 25940 20733 25941
rect 20667 25876 20668 25940
rect 20732 25876 20733 25940
rect 20667 25875 20733 25876
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 6315 25260 6381 25261
rect 6315 25196 6316 25260
rect 6380 25196 6381 25260
rect 6315 25195 6381 25196
rect 6131 23356 6197 23357
rect 6131 23292 6132 23356
rect 6196 23292 6197 23356
rect 6131 23291 6197 23292
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5395 21860 5461 21861
rect 5395 21796 5396 21860
rect 5460 21796 5461 21860
rect 5395 21795 5461 21796
rect 5610 21792 5931 22816
rect 6131 22404 6197 22405
rect 6131 22340 6132 22404
rect 6196 22340 6197 22404
rect 6131 22339 6197 22340
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5395 19820 5461 19821
rect 5395 19756 5396 19820
rect 5460 19756 5461 19820
rect 5395 19755 5461 19756
rect 5211 19004 5277 19005
rect 5211 18940 5212 19004
rect 5276 18940 5277 19004
rect 5211 18939 5277 18940
rect 5027 18052 5093 18053
rect 5027 17988 5028 18052
rect 5092 17988 5093 18052
rect 5027 17987 5093 17988
rect 4843 17780 4909 17781
rect 4843 17716 4844 17780
rect 4908 17716 4909 17780
rect 4843 17715 4909 17716
rect 4843 15740 4909 15741
rect 4843 15676 4844 15740
rect 4908 15676 4909 15740
rect 4843 15675 4909 15676
rect 4846 13565 4906 15675
rect 5214 14653 5274 18939
rect 5398 15741 5458 19755
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5395 15740 5461 15741
rect 5395 15676 5396 15740
rect 5460 15676 5461 15740
rect 5395 15675 5461 15676
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5211 14652 5277 14653
rect 5211 14588 5212 14652
rect 5276 14588 5277 14652
rect 5211 14587 5277 14588
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 4843 13564 4909 13565
rect 4843 13500 4844 13564
rect 4908 13500 4909 13564
rect 4843 13499 4909 13500
rect 5395 13564 5461 13565
rect 5395 13500 5396 13564
rect 5460 13500 5461 13564
rect 5395 13499 5461 13500
rect 5027 13156 5093 13157
rect 5027 13092 5028 13156
rect 5092 13092 5093 13156
rect 5027 13091 5093 13092
rect 5030 12698 5090 13091
rect 4659 11796 4725 11797
rect 4659 11732 4660 11796
rect 4724 11732 4725 11796
rect 4659 11731 4725 11732
rect 5398 10658 5458 13499
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 6134 11933 6194 22339
rect 6318 19685 6378 25195
rect 9811 24852 9877 24853
rect 9811 24788 9812 24852
rect 9876 24788 9877 24852
rect 9811 24787 9877 24788
rect 8707 24580 8773 24581
rect 8707 24516 8708 24580
rect 8772 24516 8773 24580
rect 8707 24515 8773 24516
rect 8155 24036 8221 24037
rect 8155 23972 8156 24036
rect 8220 23972 8221 24036
rect 8155 23971 8221 23972
rect 6499 22404 6565 22405
rect 6499 22340 6500 22404
rect 6564 22340 6565 22404
rect 6499 22339 6565 22340
rect 7971 22404 8037 22405
rect 7971 22340 7972 22404
rect 8036 22340 8037 22404
rect 7971 22339 8037 22340
rect 6315 19684 6381 19685
rect 6315 19620 6316 19684
rect 6380 19620 6381 19684
rect 6315 19619 6381 19620
rect 6318 17917 6378 19619
rect 6315 17916 6381 17917
rect 6315 17852 6316 17916
rect 6380 17852 6381 17916
rect 6315 17851 6381 17852
rect 6502 14925 6562 22339
rect 6683 21316 6749 21317
rect 6683 21252 6684 21316
rect 6748 21252 6749 21316
rect 6683 21251 6749 21252
rect 6315 14924 6381 14925
rect 6315 14860 6316 14924
rect 6380 14860 6381 14924
rect 6315 14859 6381 14860
rect 6499 14924 6565 14925
rect 6499 14860 6500 14924
rect 6564 14860 6565 14924
rect 6499 14859 6565 14860
rect 6318 13565 6378 14859
rect 6315 13564 6381 13565
rect 6315 13500 6316 13564
rect 6380 13500 6381 13564
rect 6315 13499 6381 13500
rect 6686 13290 6746 21251
rect 7238 20770 7298 21302
rect 7419 21180 7485 21181
rect 7419 21116 7420 21180
rect 7484 21116 7485 21180
rect 7419 21115 7485 21116
rect 7054 20710 7298 20770
rect 7054 19277 7114 20710
rect 7422 20634 7482 21115
rect 7238 20574 7482 20634
rect 7051 19276 7117 19277
rect 7051 19212 7052 19276
rect 7116 19212 7117 19276
rect 7051 19211 7117 19212
rect 7051 18052 7117 18053
rect 7051 17988 7052 18052
rect 7116 17988 7117 18052
rect 7051 17987 7117 17988
rect 6867 14924 6933 14925
rect 6867 14860 6868 14924
rect 6932 14860 6933 14924
rect 6867 14859 6933 14860
rect 6318 13230 6746 13290
rect 6131 11932 6197 11933
rect 6131 11868 6132 11932
rect 6196 11868 6197 11932
rect 6131 11867 6197 11868
rect 6131 11796 6197 11797
rect 6131 11732 6132 11796
rect 6196 11732 6197 11796
rect 6131 11731 6197 11732
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5398 10301 5458 10422
rect 5395 10300 5461 10301
rect 5395 10236 5396 10300
rect 5460 10236 5461 10300
rect 5395 10235 5461 10236
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 4107 9076 4173 9077
rect 4107 9012 4108 9076
rect 4172 9012 4173 9076
rect 4107 9011 4173 9012
rect 4110 8618 4170 9011
rect 5398 8941 5458 9062
rect 5395 8940 5461 8941
rect 5395 8876 5396 8940
rect 5460 8876 5461 8940
rect 5395 8875 5461 8876
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 3006 5750 3250 5810
rect 3558 8470 3802 8530
rect 3006 1597 3066 5750
rect 3187 5676 3253 5677
rect 3187 5612 3188 5676
rect 3252 5612 3253 5676
rect 3187 5611 3253 5612
rect 3003 1596 3069 1597
rect 3003 1532 3004 1596
rect 3068 1532 3069 1596
rect 3003 1531 3069 1532
rect 2819 1188 2885 1189
rect 2819 1124 2820 1188
rect 2884 1124 2885 1188
rect 3190 1138 3250 5611
rect 3558 4861 3618 8470
rect 3923 8260 3989 8261
rect 3923 8196 3924 8260
rect 3988 8196 3989 8260
rect 3923 8195 3989 8196
rect 3926 7938 3986 8195
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 6134 7581 6194 11731
rect 6131 7580 6197 7581
rect 6131 7516 6132 7580
rect 6196 7516 6197 7580
rect 6131 7515 6197 7516
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 3555 4860 3621 4861
rect 3555 4796 3556 4860
rect 3620 4796 3621 4860
rect 3555 4795 3621 4796
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 6318 4045 6378 13230
rect 6683 13156 6749 13157
rect 6683 13092 6684 13156
rect 6748 13092 6749 13156
rect 6683 13091 6749 13092
rect 6499 11932 6565 11933
rect 6499 11868 6500 11932
rect 6564 11868 6565 11932
rect 6499 11867 6565 11868
rect 6502 4861 6562 11867
rect 6686 9077 6746 13091
rect 6683 9076 6749 9077
rect 6683 9012 6684 9076
rect 6748 9012 6749 9076
rect 6683 9011 6749 9012
rect 6870 8938 6930 14859
rect 7054 13701 7114 17987
rect 7051 13700 7117 13701
rect 7051 13636 7052 13700
rect 7116 13636 7117 13700
rect 7051 13635 7117 13636
rect 7051 13020 7117 13021
rect 7051 12956 7052 13020
rect 7116 12956 7117 13020
rect 7051 12955 7117 12956
rect 7054 10981 7114 12955
rect 7051 10980 7117 10981
rect 7051 10916 7052 10980
rect 7116 10916 7117 10980
rect 7051 10915 7117 10916
rect 6686 8878 6930 8938
rect 6499 4860 6565 4861
rect 6499 4796 6500 4860
rect 6564 4796 6565 4860
rect 6499 4795 6565 4796
rect 6686 4538 6746 8878
rect 7051 8804 7117 8805
rect 7051 8740 7052 8804
rect 7116 8740 7117 8804
rect 7051 8739 7117 8740
rect 6315 4044 6381 4045
rect 6315 3980 6316 4044
rect 6380 3980 6381 4044
rect 6315 3979 6381 3980
rect 6686 3637 6746 4302
rect 6683 3636 6749 3637
rect 6683 3572 6684 3636
rect 6748 3572 6749 3636
rect 6683 3571 6749 3572
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 2819 1123 2885 1124
rect 7054 645 7114 8739
rect 7238 4317 7298 20574
rect 7606 13157 7666 19262
rect 7974 18730 8034 22339
rect 8158 22133 8218 23971
rect 8339 22676 8405 22677
rect 8339 22612 8340 22676
rect 8404 22612 8405 22676
rect 8339 22611 8405 22612
rect 8155 22132 8221 22133
rect 8155 22068 8156 22132
rect 8220 22068 8221 22132
rect 8155 22067 8221 22068
rect 8342 20501 8402 22611
rect 8710 22405 8770 24515
rect 9443 24308 9509 24309
rect 9443 24244 9444 24308
rect 9508 24244 9509 24308
rect 9443 24243 9509 24244
rect 9446 23354 9506 24243
rect 9446 23294 9644 23354
rect 9075 23220 9141 23221
rect 9075 23156 9076 23220
rect 9140 23156 9141 23220
rect 9075 23155 9141 23156
rect 8707 22404 8773 22405
rect 8707 22340 8708 22404
rect 8772 22340 8773 22404
rect 8707 22339 8773 22340
rect 9078 22218 9138 23155
rect 9584 22813 9644 23294
rect 9443 22812 9509 22813
rect 9443 22748 9444 22812
rect 9508 22748 9509 22812
rect 9443 22747 9509 22748
rect 9581 22812 9647 22813
rect 9581 22748 9582 22812
rect 9646 22748 9647 22812
rect 9581 22747 9647 22748
rect 8707 22132 8773 22133
rect 8707 22068 8708 22132
rect 8772 22068 8773 22132
rect 8707 22067 8773 22068
rect 8710 21725 8770 22067
rect 8707 21724 8773 21725
rect 8707 21660 8708 21724
rect 8772 21660 8773 21724
rect 8707 21659 8773 21660
rect 9446 21450 9506 22747
rect 9446 21390 9690 21450
rect 8339 20500 8405 20501
rect 8339 20436 8340 20500
rect 8404 20436 8405 20500
rect 8339 20435 8405 20436
rect 9630 20229 9690 21390
rect 8155 20228 8221 20229
rect 8155 20164 8156 20228
rect 8220 20164 8221 20228
rect 8155 20163 8221 20164
rect 9627 20228 9693 20229
rect 9627 20164 9628 20228
rect 9692 20164 9693 20228
rect 9627 20163 9693 20164
rect 7790 18670 8034 18730
rect 7790 17917 7850 18670
rect 7787 17916 7853 17917
rect 7787 17852 7788 17916
rect 7852 17852 7853 17916
rect 7787 17851 7853 17852
rect 7603 13156 7669 13157
rect 7603 13092 7604 13156
rect 7668 13092 7669 13156
rect 7603 13091 7669 13092
rect 7235 4316 7301 4317
rect 7235 4252 7236 4316
rect 7300 4252 7301 4316
rect 7235 4251 7301 4252
rect 7790 1461 7850 17851
rect 8158 16285 8218 20163
rect 9814 20090 9874 24787
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 9995 23492 10061 23493
rect 9995 23428 9996 23492
rect 10060 23428 10061 23492
rect 9995 23427 10061 23428
rect 9998 21997 10058 23427
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 11651 23084 11717 23085
rect 11651 23020 11652 23084
rect 11716 23020 11717 23084
rect 11651 23019 11717 23020
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 9995 21996 10061 21997
rect 9995 21932 9996 21996
rect 10060 21932 10061 21996
rect 9995 21931 10061 21932
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 11654 20637 11714 23019
rect 11651 20636 11717 20637
rect 11651 20572 11652 20636
rect 11716 20572 11717 20636
rect 11651 20571 11717 20572
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 9995 20092 10061 20093
rect 9995 20090 9996 20092
rect 9814 20030 9996 20090
rect 9995 20028 9996 20030
rect 10060 20028 10061 20092
rect 9995 20027 10061 20028
rect 9995 19820 10061 19821
rect 9995 19756 9996 19820
rect 10060 19756 10061 19820
rect 9995 19755 10061 19756
rect 9811 18188 9877 18189
rect 9811 18124 9812 18188
rect 9876 18124 9877 18188
rect 9811 18123 9877 18124
rect 8523 17852 8524 17902
rect 8588 17852 8589 17902
rect 8523 17851 8589 17852
rect 9814 16693 9874 18123
rect 9811 16692 9877 16693
rect 9811 16628 9812 16692
rect 9876 16628 9877 16692
rect 9811 16627 9877 16628
rect 8155 16284 8221 16285
rect 8155 16220 8156 16284
rect 8220 16220 8221 16284
rect 8155 16219 8221 16220
rect 9627 15740 9693 15741
rect 9627 15676 9628 15740
rect 9692 15676 9693 15740
rect 9627 15675 9693 15676
rect 9630 15418 9690 15675
rect 8523 14516 8589 14517
rect 8523 14452 8524 14516
rect 8588 14452 8589 14516
rect 8523 14451 8589 14452
rect 7971 13020 8037 13021
rect 7971 12956 7972 13020
rect 8036 12956 8037 13020
rect 7971 12955 8037 12956
rect 7974 12477 8034 12955
rect 7971 12476 8037 12477
rect 7971 12412 7972 12476
rect 8036 12412 8037 12476
rect 7971 12411 8037 12412
rect 8158 12341 8218 13142
rect 8155 12340 8221 12341
rect 8155 12276 8156 12340
rect 8220 12276 8221 12340
rect 8155 12275 8221 12276
rect 8526 10845 8586 14451
rect 8891 12476 8957 12477
rect 8891 12412 8892 12476
rect 8956 12412 8957 12476
rect 8891 12411 8957 12412
rect 8894 11525 8954 12411
rect 9443 12340 9509 12341
rect 9443 12276 9444 12340
rect 9508 12276 9509 12340
rect 9443 12275 9509 12276
rect 8891 11524 8957 11525
rect 8891 11460 8892 11524
rect 8956 11460 8957 11524
rect 8891 11459 8957 11460
rect 8523 10844 8589 10845
rect 8523 10780 8524 10844
rect 8588 10780 8589 10844
rect 8523 10779 8589 10780
rect 8158 6765 8218 7022
rect 8155 6764 8221 6765
rect 8155 6700 8156 6764
rect 8220 6700 8221 6764
rect 8155 6699 8221 6700
rect 9446 5541 9506 12275
rect 9998 10301 10058 19755
rect 10277 19072 10597 20096
rect 11099 19548 11165 19549
rect 11099 19484 11100 19548
rect 11164 19484 11165 19548
rect 11099 19483 11165 19484
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10731 17372 10797 17373
rect 10731 17308 10732 17372
rect 10796 17308 10797 17372
rect 10731 17307 10797 17308
rect 10734 16965 10794 17307
rect 10731 16964 10797 16965
rect 10731 16900 10732 16964
rect 10796 16900 10797 16964
rect 10731 16899 10797 16900
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10731 16420 10797 16421
rect 10731 16356 10732 16420
rect 10796 16356 10797 16420
rect 10731 16355 10797 16356
rect 10915 16420 10981 16421
rect 10915 16356 10916 16420
rect 10980 16356 10981 16420
rect 10915 16355 10981 16356
rect 10734 15877 10794 16355
rect 10731 15876 10797 15877
rect 10731 15812 10732 15876
rect 10796 15812 10797 15876
rect 10731 15811 10797 15812
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10734 11525 10794 15811
rect 10731 11524 10797 11525
rect 10731 11460 10732 11524
rect 10796 11460 10797 11524
rect 10731 11459 10797 11460
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9995 10300 10061 10301
rect 9995 10236 9996 10300
rect 10060 10236 10061 10300
rect 9995 10235 10061 10236
rect 9995 9348 10061 9349
rect 9995 9284 9996 9348
rect 10060 9284 10061 9348
rect 9995 9283 10061 9284
rect 9998 5541 10058 9283
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10731 7852 10797 7853
rect 10731 7788 10732 7852
rect 10796 7788 10797 7852
rect 10731 7787 10797 7788
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10734 6901 10794 7787
rect 10731 6900 10797 6901
rect 10731 6836 10732 6900
rect 10796 6836 10797 6900
rect 10731 6835 10797 6836
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 9443 5540 9509 5541
rect 9443 5476 9444 5540
rect 9508 5476 9509 5540
rect 9443 5475 9509 5476
rect 9995 5540 10061 5541
rect 9995 5476 9996 5540
rect 10060 5476 10061 5540
rect 9995 5475 10061 5476
rect 9998 3909 10058 5475
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 9995 3908 10061 3909
rect 9995 3844 9996 3908
rect 10060 3844 10061 3908
rect 9995 3843 10061 3844
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10734 2957 10794 6835
rect 10918 5677 10978 16355
rect 11102 12613 11162 19483
rect 11654 19005 11714 20571
rect 13307 20364 13373 20365
rect 13307 20300 13308 20364
rect 13372 20300 13373 20364
rect 13307 20299 13373 20300
rect 13310 20178 13370 20299
rect 12019 19684 12085 19685
rect 12019 19620 12020 19684
rect 12084 19620 12085 19684
rect 12019 19619 12085 19620
rect 11835 19140 11901 19141
rect 11835 19076 11836 19140
rect 11900 19076 11901 19140
rect 12022 19138 12082 19619
rect 12203 19140 12269 19141
rect 12203 19138 12204 19140
rect 12022 19078 12204 19138
rect 11835 19075 11901 19076
rect 12203 19076 12204 19078
rect 12268 19076 12269 19140
rect 12203 19075 12269 19076
rect 11651 19004 11717 19005
rect 11651 18940 11652 19004
rect 11716 18940 11717 19004
rect 11651 18939 11717 18940
rect 11283 16692 11349 16693
rect 11283 16628 11284 16692
rect 11348 16628 11349 16692
rect 11283 16627 11349 16628
rect 11099 12612 11165 12613
rect 11099 12548 11100 12612
rect 11164 12548 11165 12612
rect 11099 12547 11165 12548
rect 11286 10437 11346 16627
rect 11283 10436 11349 10437
rect 11283 10372 11284 10436
rect 11348 10372 11349 10436
rect 11283 10371 11349 10372
rect 11838 9298 11898 19075
rect 14046 17509 14106 25382
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 20299 24580 20365 24581
rect 20299 24516 20300 24580
rect 20364 24516 20365 24580
rect 20299 24515 20365 24516
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 16619 23492 16685 23493
rect 16619 23428 16620 23492
rect 16684 23428 16685 23492
rect 16619 23427 16685 23428
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 15515 20772 15581 20773
rect 15515 20708 15516 20772
rect 15580 20708 15581 20772
rect 15515 20707 15581 20708
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14595 18460 14661 18461
rect 14595 18396 14596 18460
rect 14660 18396 14661 18460
rect 14595 18395 14661 18396
rect 14043 17508 14109 17509
rect 14043 17444 14044 17508
rect 14108 17444 14109 17508
rect 14043 17443 14109 17444
rect 11099 8260 11165 8261
rect 11099 8196 11100 8260
rect 11164 8196 11165 8260
rect 11099 8195 11165 8196
rect 10915 5676 10981 5677
rect 10915 5612 10916 5676
rect 10980 5612 10981 5676
rect 10915 5611 10981 5612
rect 11102 4045 11162 8195
rect 11838 6578 11898 9062
rect 12206 6765 12266 16542
rect 14046 13157 14106 17443
rect 14043 13156 14109 13157
rect 14043 13092 14044 13156
rect 14108 13092 14109 13156
rect 14043 13091 14109 13092
rect 14598 12477 14658 18395
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14595 12476 14661 12477
rect 14595 12412 14596 12476
rect 14660 12412 14661 12476
rect 14595 12411 14661 12412
rect 12387 12340 12453 12341
rect 12387 12276 12388 12340
rect 12452 12276 12453 12340
rect 12387 12275 12453 12276
rect 12390 11389 12450 12275
rect 12387 11388 12453 11389
rect 12387 11324 12388 11388
rect 12452 11324 12453 11388
rect 12387 11323 12453 11324
rect 14598 10845 14658 12411
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 15518 10981 15578 20707
rect 16251 18052 16317 18053
rect 16251 17988 16252 18052
rect 16316 17988 16317 18052
rect 16251 17987 16317 17988
rect 15515 10980 15581 10981
rect 15515 10916 15516 10980
rect 15580 10916 15581 10980
rect 15515 10915 15581 10916
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14595 10844 14661 10845
rect 14595 10780 14596 10844
rect 14660 10780 14661 10844
rect 14595 10779 14661 10780
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 13859 8940 13925 8941
rect 13859 8876 13860 8940
rect 13924 8876 13925 8940
rect 13859 8875 13925 8876
rect 12203 6764 12269 6765
rect 12203 6700 12204 6764
rect 12268 6700 12269 6764
rect 12203 6699 12269 6700
rect 13123 5404 13189 5405
rect 13123 5340 13124 5404
rect 13188 5340 13189 5404
rect 13123 5339 13189 5340
rect 13126 5218 13186 5339
rect 11099 4044 11165 4045
rect 11099 3980 11100 4044
rect 11164 3980 11165 4044
rect 11099 3979 11165 3980
rect 12387 4044 12453 4045
rect 12387 3980 12388 4044
rect 12452 3980 12453 4044
rect 12387 3979 12453 3980
rect 10731 2956 10797 2957
rect 10731 2892 10732 2956
rect 10796 2892 10797 2956
rect 10731 2891 10797 2892
rect 12390 2821 12450 3979
rect 13862 3501 13922 8875
rect 14230 7717 14290 9742
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14227 7716 14293 7717
rect 14227 7652 14228 7716
rect 14292 7652 14293 7716
rect 14227 7651 14293 7652
rect 14598 4861 14658 7702
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 16254 5898 16314 17987
rect 16622 17645 16682 23427
rect 19610 23424 19930 24448
rect 20115 23492 20181 23493
rect 20115 23428 20116 23492
rect 20180 23428 20181 23492
rect 20115 23427 20181 23428
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 18091 21996 18157 21997
rect 18091 21932 18092 21996
rect 18156 21932 18157 21996
rect 18091 21931 18157 21932
rect 18094 20773 18154 21931
rect 18091 20772 18157 20773
rect 18091 20708 18092 20772
rect 18156 20708 18157 20772
rect 18091 20707 18157 20708
rect 17171 20092 17237 20093
rect 17171 20028 17172 20092
rect 17236 20028 17237 20092
rect 17171 20027 17237 20028
rect 16619 17644 16685 17645
rect 16619 17580 16620 17644
rect 16684 17580 16685 17644
rect 16619 17579 16685 17580
rect 16619 14516 16685 14517
rect 16619 14452 16620 14516
rect 16684 14452 16685 14516
rect 16619 14451 16685 14452
rect 16622 13973 16682 14451
rect 16619 13972 16685 13973
rect 16619 13908 16620 13972
rect 16684 13908 16685 13972
rect 16619 13907 16685 13908
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14595 4860 14661 4861
rect 14595 4796 14596 4860
rect 14660 4796 14661 4860
rect 14595 4795 14661 4796
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 13859 3500 13925 3501
rect 13859 3436 13860 3500
rect 13924 3436 13925 3500
rect 13859 3435 13925 3436
rect 14944 3296 15264 4320
rect 16806 3909 16866 6342
rect 16803 3908 16869 3909
rect 16803 3844 16804 3908
rect 16868 3844 16869 3908
rect 16803 3843 16869 3844
rect 17174 3773 17234 20027
rect 19011 17372 19077 17373
rect 19011 17308 19012 17372
rect 19076 17308 19077 17372
rect 19011 17307 19077 17308
rect 19014 8397 19074 17307
rect 19382 17101 19442 21982
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19379 17100 19445 17101
rect 19379 17036 19380 17100
rect 19444 17036 19445 17100
rect 19379 17035 19445 17036
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 20118 13701 20178 23427
rect 20302 17370 20362 24515
rect 20483 23628 20549 23629
rect 20483 23564 20484 23628
rect 20548 23564 20549 23628
rect 20483 23563 20549 23564
rect 20486 19005 20546 23563
rect 20670 22405 20730 25875
rect 26923 25668 26989 25669
rect 26923 25618 26924 25668
rect 26988 25618 26989 25668
rect 21035 25260 21101 25261
rect 21035 25196 21036 25260
rect 21100 25196 21101 25260
rect 21035 25195 21101 25196
rect 20851 23900 20917 23901
rect 20851 23836 20852 23900
rect 20916 23836 20917 23900
rect 20851 23835 20917 23836
rect 20667 22404 20733 22405
rect 20667 22340 20668 22404
rect 20732 22340 20733 22404
rect 20667 22339 20733 22340
rect 20854 22133 20914 23835
rect 20851 22132 20917 22133
rect 20851 22068 20852 22132
rect 20916 22068 20917 22132
rect 20851 22067 20917 22068
rect 21038 21725 21098 25195
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 22323 24172 22389 24173
rect 22323 24108 22324 24172
rect 22388 24108 22389 24172
rect 22323 24107 22389 24108
rect 21955 23900 22021 23901
rect 21955 23836 21956 23900
rect 22020 23836 22021 23900
rect 21955 23835 22021 23836
rect 21958 23578 22018 23835
rect 21587 23356 21653 23357
rect 21587 23292 21588 23356
rect 21652 23292 21653 23356
rect 21587 23291 21653 23292
rect 20667 21724 20733 21725
rect 20667 21660 20668 21724
rect 20732 21660 20733 21724
rect 20667 21659 20733 21660
rect 21035 21724 21101 21725
rect 21035 21660 21036 21724
rect 21100 21660 21101 21724
rect 21035 21659 21101 21660
rect 20483 19004 20549 19005
rect 20483 18940 20484 19004
rect 20548 18940 20549 19004
rect 20483 18939 20549 18940
rect 20670 17917 20730 21659
rect 21403 21588 21469 21589
rect 21403 21524 21404 21588
rect 21468 21524 21469 21588
rect 21403 21523 21469 21524
rect 21406 21045 21466 21523
rect 21403 21044 21469 21045
rect 21403 20980 21404 21044
rect 21468 20980 21469 21044
rect 21403 20979 21469 20980
rect 20851 20364 20917 20365
rect 20851 20300 20852 20364
rect 20916 20300 20917 20364
rect 20851 20299 20917 20300
rect 20854 18730 20914 20299
rect 21219 20228 21285 20229
rect 21219 20164 21220 20228
rect 21284 20164 21285 20228
rect 21219 20163 21285 20164
rect 21222 19498 21282 20163
rect 21219 19004 21285 19005
rect 21219 18940 21220 19004
rect 21284 18940 21285 19004
rect 21219 18939 21285 18940
rect 20854 18670 21098 18730
rect 20667 17916 20733 17917
rect 20667 17852 20668 17916
rect 20732 17852 20733 17916
rect 20667 17851 20733 17852
rect 20302 17310 20546 17370
rect 20299 17100 20365 17101
rect 20299 17036 20300 17100
rect 20364 17036 20365 17100
rect 20299 17035 20365 17036
rect 20302 14381 20362 17035
rect 20299 14380 20365 14381
rect 20299 14316 20300 14380
rect 20364 14316 20365 14380
rect 20299 14315 20365 14316
rect 20299 13972 20365 13973
rect 20299 13908 20300 13972
rect 20364 13908 20365 13972
rect 20299 13907 20365 13908
rect 20115 13700 20181 13701
rect 20115 13636 20116 13700
rect 20180 13636 20181 13700
rect 20115 13635 20181 13636
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19379 13564 19445 13565
rect 19379 13500 19380 13564
rect 19444 13500 19445 13564
rect 19379 13499 19445 13500
rect 19382 13378 19442 13499
rect 19379 12884 19445 12885
rect 19379 12820 19380 12884
rect 19444 12820 19445 12884
rect 19379 12819 19445 12820
rect 19382 12018 19442 12819
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 20302 11389 20362 13907
rect 20299 11388 20365 11389
rect 20299 11324 20300 11388
rect 20364 11324 20365 11388
rect 20299 11323 20365 11324
rect 20486 10709 20546 17310
rect 20667 16148 20733 16149
rect 20667 16084 20668 16148
rect 20732 16084 20733 16148
rect 20667 16083 20733 16084
rect 20670 15061 20730 16083
rect 20667 15060 20733 15061
rect 20667 14996 20668 15060
rect 20732 14996 20733 15060
rect 20667 14995 20733 14996
rect 20851 13972 20917 13973
rect 20851 13908 20852 13972
rect 20916 13908 20917 13972
rect 20851 13907 20917 13908
rect 20667 13700 20733 13701
rect 20667 13636 20668 13700
rect 20732 13636 20733 13700
rect 20667 13635 20733 13636
rect 20115 10708 20181 10709
rect 20115 10644 20116 10708
rect 20180 10644 20181 10708
rect 20115 10643 20181 10644
rect 20483 10708 20549 10709
rect 20483 10644 20484 10708
rect 20548 10644 20549 10708
rect 20483 10643 20549 10644
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19011 8396 19077 8397
rect 19011 8332 19012 8396
rect 19076 8332 19077 8396
rect 19011 8331 19077 8332
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 20118 7037 20178 10643
rect 20670 10570 20730 13635
rect 20486 10510 20730 10570
rect 20486 7717 20546 10510
rect 20483 7716 20549 7717
rect 20483 7652 20484 7716
rect 20548 7652 20549 7716
rect 20483 7651 20549 7652
rect 20115 7036 20181 7037
rect 20115 6972 20116 7036
rect 20180 6972 20181 7036
rect 20115 6971 20181 6972
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 20854 5133 20914 13907
rect 21038 13701 21098 18670
rect 21035 13700 21101 13701
rect 21035 13636 21036 13700
rect 21100 13636 21101 13700
rect 21035 13635 21101 13636
rect 21035 12340 21101 12341
rect 21035 12276 21036 12340
rect 21100 12276 21101 12340
rect 21222 12338 21282 18939
rect 21403 18052 21469 18053
rect 21403 17988 21404 18052
rect 21468 17988 21469 18052
rect 21403 17987 21469 17988
rect 21406 15877 21466 17987
rect 21403 15876 21469 15877
rect 21403 15812 21404 15876
rect 21468 15812 21469 15876
rect 21403 15811 21469 15812
rect 21222 12278 21466 12338
rect 21035 12275 21101 12276
rect 21038 11797 21098 12275
rect 21219 11932 21285 11933
rect 21219 11868 21220 11932
rect 21284 11868 21285 11932
rect 21219 11867 21285 11868
rect 21035 11796 21101 11797
rect 21035 11732 21036 11796
rect 21100 11732 21101 11796
rect 21035 11731 21101 11732
rect 20851 5132 20917 5133
rect 20851 5068 20852 5132
rect 20916 5068 20917 5132
rect 20851 5067 20917 5068
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 20483 3908 20549 3909
rect 20483 3844 20484 3908
rect 20548 3844 20549 3908
rect 20483 3843 20549 3844
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 17171 3772 17237 3773
rect 17171 3708 17172 3772
rect 17236 3708 17237 3772
rect 17171 3707 17237 3708
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 12387 2820 12453 2821
rect 12387 2756 12388 2820
rect 12452 2756 12453 2820
rect 12387 2755 12453 2756
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 2208 15264 3232
rect 16619 3228 16685 3229
rect 16619 3164 16620 3228
rect 16684 3164 16685 3228
rect 16619 3163 16685 3164
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 16622 1818 16682 3163
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 20486 2498 20546 3843
rect 21038 3773 21098 11731
rect 21222 8397 21282 11867
rect 21406 9893 21466 12278
rect 21403 9892 21469 9893
rect 21403 9828 21404 9892
rect 21468 9828 21469 9892
rect 21403 9827 21469 9828
rect 21219 8396 21285 8397
rect 21219 8332 21220 8396
rect 21284 8332 21285 8396
rect 21219 8331 21285 8332
rect 21590 8261 21650 23291
rect 21771 22404 21837 22405
rect 21771 22340 21772 22404
rect 21836 22340 21837 22404
rect 21771 22339 21837 22340
rect 21774 18053 21834 22339
rect 22326 19549 22386 24107
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 23059 23492 23125 23493
rect 23059 23428 23060 23492
rect 23124 23428 23125 23492
rect 23059 23427 23125 23428
rect 23795 23492 23861 23493
rect 23795 23428 23796 23492
rect 23860 23428 23861 23492
rect 23795 23427 23861 23428
rect 22691 22132 22757 22133
rect 22691 22068 22692 22132
rect 22756 22068 22757 22132
rect 22691 22067 22757 22068
rect 22323 19548 22389 19549
rect 22323 19484 22324 19548
rect 22388 19484 22389 19548
rect 22323 19483 22389 19484
rect 21771 18052 21837 18053
rect 21771 17988 21772 18052
rect 21836 17988 21837 18052
rect 22139 18052 22205 18053
rect 22139 18050 22140 18052
rect 21771 17987 21837 17988
rect 21958 17990 22140 18050
rect 21958 17458 22018 17990
rect 22139 17988 22140 17990
rect 22204 17988 22205 18052
rect 22139 17987 22205 17988
rect 21771 17100 21837 17101
rect 21771 17036 21772 17100
rect 21836 17036 21837 17100
rect 21771 17035 21837 17036
rect 21587 8260 21653 8261
rect 21587 8196 21588 8260
rect 21652 8196 21653 8260
rect 21587 8195 21653 8196
rect 21035 3772 21101 3773
rect 21035 3708 21036 3772
rect 21100 3708 21101 3772
rect 21035 3707 21101 3708
rect 21774 2685 21834 17035
rect 22323 16692 22389 16693
rect 22323 16690 22324 16692
rect 22142 16630 22324 16690
rect 21955 15876 22021 15877
rect 21955 15812 21956 15876
rect 22020 15812 22021 15876
rect 21955 15811 22021 15812
rect 21958 5130 22018 15811
rect 22142 14653 22202 16630
rect 22323 16628 22324 16630
rect 22388 16628 22389 16692
rect 22323 16627 22389 16628
rect 22694 15418 22754 22067
rect 22875 21724 22941 21725
rect 22875 21660 22876 21724
rect 22940 21660 22941 21724
rect 22875 21659 22941 21660
rect 22878 15605 22938 21659
rect 23062 17370 23122 23427
rect 23427 19276 23493 19277
rect 23427 19212 23428 19276
rect 23492 19212 23493 19276
rect 23427 19211 23493 19212
rect 23430 18138 23490 19211
rect 23062 17310 23490 17370
rect 22875 15604 22941 15605
rect 22875 15540 22876 15604
rect 22940 15540 22941 15604
rect 22875 15539 22941 15540
rect 22323 14924 22389 14925
rect 22323 14860 22324 14924
rect 22388 14860 22389 14924
rect 22323 14859 22389 14860
rect 22139 14652 22205 14653
rect 22139 14588 22140 14652
rect 22204 14588 22205 14652
rect 22139 14587 22205 14588
rect 22139 14244 22205 14245
rect 22139 14180 22140 14244
rect 22204 14180 22205 14244
rect 22139 14179 22205 14180
rect 22142 10301 22202 14179
rect 22326 10845 22386 14859
rect 22507 13564 22573 13565
rect 22507 13500 22508 13564
rect 22572 13500 22573 13564
rect 22507 13499 22573 13500
rect 22323 10844 22389 10845
rect 22323 10780 22324 10844
rect 22388 10780 22389 10844
rect 22323 10779 22389 10780
rect 22139 10300 22205 10301
rect 22139 10236 22140 10300
rect 22204 10236 22205 10300
rect 22139 10235 22205 10236
rect 22323 10300 22389 10301
rect 22323 10236 22324 10300
rect 22388 10236 22389 10300
rect 22323 10235 22389 10236
rect 22326 9893 22386 10235
rect 22323 9892 22389 9893
rect 22323 9828 22324 9892
rect 22388 9828 22389 9892
rect 22323 9827 22389 9828
rect 22510 8397 22570 13499
rect 22694 11930 22754 15182
rect 23430 13565 23490 17310
rect 23611 17100 23677 17101
rect 23611 17036 23612 17100
rect 23676 17036 23677 17100
rect 23611 17035 23677 17036
rect 23614 14653 23674 17035
rect 23611 14652 23677 14653
rect 23611 14588 23612 14652
rect 23676 14588 23677 14652
rect 23611 14587 23677 14588
rect 23427 13564 23493 13565
rect 23427 13500 23428 13564
rect 23492 13500 23493 13564
rect 23427 13499 23493 13500
rect 22694 11870 23490 11930
rect 22507 8396 22573 8397
rect 22507 8332 22508 8396
rect 22572 8332 22573 8396
rect 22507 8331 22573 8332
rect 23430 7445 23490 11870
rect 23798 11250 23858 23427
rect 23979 23084 24045 23085
rect 23979 23020 23980 23084
rect 24044 23020 24045 23084
rect 23979 23019 24045 23020
rect 23982 15877 24042 23019
rect 24277 22880 24597 23904
rect 24715 23492 24781 23493
rect 24715 23428 24716 23492
rect 24780 23428 24781 23492
rect 24715 23427 24781 23428
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24718 17101 24778 23427
rect 25267 21724 25333 21725
rect 25267 21660 25268 21724
rect 25332 21660 25333 21724
rect 25267 21659 25333 21660
rect 24899 19140 24965 19141
rect 24899 19076 24900 19140
rect 24964 19076 24965 19140
rect 24899 19075 24965 19076
rect 24715 17100 24781 17101
rect 24715 17036 24716 17100
rect 24780 17036 24781 17100
rect 24715 17035 24781 17036
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 23979 15876 24045 15877
rect 23979 15812 23980 15876
rect 24044 15812 24045 15876
rect 23979 15811 24045 15812
rect 23614 11190 23858 11250
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24715 13564 24781 13565
rect 24715 13500 24716 13564
rect 24780 13500 24781 13564
rect 24715 13499 24781 13500
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 23614 8261 23674 11190
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 23979 10844 24045 10845
rect 23979 10780 23980 10844
rect 24044 10780 24045 10844
rect 23979 10779 24045 10780
rect 23982 10658 24042 10779
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 23979 9484 24045 9485
rect 23979 9420 23980 9484
rect 24044 9420 24045 9484
rect 23979 9419 24045 9420
rect 23982 8530 24042 9419
rect 23798 8470 24042 8530
rect 24277 8736 24597 9760
rect 24718 9485 24778 13499
rect 24902 11933 24962 19075
rect 25083 14244 25149 14245
rect 25083 14180 25084 14244
rect 25148 14180 25149 14244
rect 25083 14179 25149 14180
rect 24899 11932 24965 11933
rect 24899 11868 24900 11932
rect 24964 11868 24965 11932
rect 24899 11867 24965 11868
rect 24899 11388 24965 11389
rect 24899 11324 24900 11388
rect 24964 11324 24965 11388
rect 24899 11323 24965 11324
rect 24715 9484 24781 9485
rect 24715 9420 24716 9484
rect 24780 9420 24781 9484
rect 24715 9419 24781 9420
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 23611 8260 23677 8261
rect 23611 8196 23612 8260
rect 23676 8196 23677 8260
rect 23611 8195 23677 8196
rect 23798 7850 23858 8470
rect 23614 7790 23858 7850
rect 23979 7852 24045 7853
rect 23427 7444 23493 7445
rect 23427 7380 23428 7444
rect 23492 7380 23493 7444
rect 23427 7379 23493 7380
rect 22139 5132 22205 5133
rect 22139 5130 22140 5132
rect 21958 5070 22140 5130
rect 22139 5068 22140 5070
rect 22204 5068 22205 5132
rect 23614 5130 23674 7790
rect 23979 7788 23980 7852
rect 24044 7788 24045 7852
rect 23979 7787 24045 7788
rect 23982 7258 24042 7787
rect 24277 7648 24597 8672
rect 24715 8260 24781 8261
rect 24715 8196 24716 8260
rect 24780 8196 24781 8260
rect 24715 8195 24781 8196
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 23979 6220 24045 6221
rect 23979 6156 23980 6220
rect 24044 6156 24045 6220
rect 23979 6155 24045 6156
rect 23982 5898 24042 6155
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 23614 5070 23858 5130
rect 22139 5067 22205 5068
rect 23798 4045 23858 5070
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 23795 4044 23861 4045
rect 23795 3980 23796 4044
rect 23860 3980 23861 4044
rect 23795 3979 23861 3980
rect 24277 3296 24597 4320
rect 24718 3637 24778 8195
rect 24902 5405 24962 11323
rect 25086 8669 25146 14179
rect 25083 8668 25149 8669
rect 25083 8604 25084 8668
rect 25148 8604 25149 8668
rect 25083 8603 25149 8604
rect 24899 5404 24965 5405
rect 24899 5340 24900 5404
rect 24964 5340 24965 5404
rect 24899 5339 24965 5340
rect 24715 3636 24781 3637
rect 24715 3572 24716 3636
rect 24780 3572 24781 3636
rect 24715 3571 24781 3572
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 21771 2684 21837 2685
rect 21771 2620 21772 2684
rect 21836 2620 21837 2684
rect 21771 2619 21837 2620
rect 24277 2208 24597 3232
rect 25270 3229 25330 21659
rect 26003 19820 26069 19821
rect 26003 19756 26004 19820
rect 26068 19756 26069 19820
rect 26003 19755 26069 19756
rect 26006 13565 26066 19755
rect 26003 13564 26069 13565
rect 26003 13500 26004 13564
rect 26068 13500 26069 13564
rect 26003 13499 26069 13500
rect 25267 3228 25333 3229
rect 25267 3164 25268 3228
rect 25332 3164 25333 3228
rect 25267 3163 25333 3164
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 7787 1460 7853 1461
rect 7787 1396 7788 1460
rect 7852 1396 7853 1460
rect 7787 1395 7853 1396
rect 7051 644 7117 645
rect 7051 580 7052 644
rect 7116 580 7117 644
rect 7051 579 7117 580
<< via4 >>
rect 2550 20092 2786 20178
rect 2550 20028 2636 20092
rect 2636 20028 2700 20092
rect 2700 20028 2786 20092
rect 2550 19942 2786 20028
rect 1814 16692 2050 16778
rect 1814 16628 1900 16692
rect 1900 16628 1964 16692
rect 1964 16628 2050 16692
rect 1814 16542 2050 16628
rect 2182 1582 2418 1818
rect 6046 26062 6282 26298
rect 26286 26212 26522 26298
rect 26286 26148 26372 26212
rect 26372 26148 26436 26212
rect 26436 26148 26522 26212
rect 26286 26062 26522 26148
rect 4942 12462 5178 12698
rect 4942 11932 5178 12018
rect 4942 11868 5028 11932
rect 5028 11868 5092 11932
rect 5092 11868 5178 11932
rect 4942 11782 5178 11868
rect 7150 21302 7386 21538
rect 5310 10422 5546 10658
rect 5310 9062 5546 9298
rect 4022 8382 4258 8618
rect 3838 7702 4074 7938
rect 5310 5812 5546 5898
rect 5310 5748 5396 5812
rect 5396 5748 5460 5812
rect 5460 5748 5546 5812
rect 5310 5662 5546 5748
rect 6598 4302 6834 4538
rect 3838 2412 4074 2498
rect 3838 2348 3924 2412
rect 3924 2348 3988 2412
rect 3988 2348 4074 2412
rect 3838 2262 4074 2348
rect 3102 902 3338 1138
rect 7518 19262 7754 19498
rect 8990 21982 9226 22218
rect 13958 25382 14194 25618
rect 8438 17916 8674 18138
rect 8438 17902 8524 17916
rect 8524 17902 8588 17916
rect 8588 17902 8674 17916
rect 9542 15182 9778 15418
rect 8070 13142 8306 13378
rect 8070 7022 8306 7258
rect 10830 20092 11066 20178
rect 10830 20028 10916 20092
rect 10916 20028 10980 20092
rect 10980 20028 11066 20092
rect 10830 19942 11066 20028
rect 13222 19942 13458 20178
rect 11382 17372 11618 17458
rect 11382 17308 11468 17372
rect 11468 17308 11532 17372
rect 11532 17308 11618 17372
rect 11382 17222 11618 17308
rect 18558 23492 18794 23578
rect 18558 23428 18644 23492
rect 18644 23428 18708 23492
rect 18708 23428 18794 23492
rect 12118 16542 12354 16778
rect 11750 9062 11986 9298
rect 14142 9742 14378 9978
rect 11750 6342 11986 6578
rect 13038 4982 13274 5218
rect 14510 7702 14746 7938
rect 18558 23342 18794 23428
rect 19294 21982 19530 22218
rect 16718 8532 16954 8618
rect 16718 8468 16804 8532
rect 16804 8468 16868 8532
rect 16868 8468 16954 8532
rect 16718 8382 16954 8468
rect 16718 6342 16954 6578
rect 16166 5662 16402 5898
rect 26838 25604 26924 25618
rect 26924 25604 26988 25618
rect 26988 25604 27074 25618
rect 26838 25382 27074 25604
rect 21870 23342 22106 23578
rect 20950 21452 21186 21538
rect 20950 21388 21036 21452
rect 21036 21388 21100 21452
rect 21100 21388 21186 21452
rect 20950 21302 21186 21388
rect 21134 19262 21370 19498
rect 19294 13142 19530 13378
rect 19294 11782 19530 12018
rect 21870 17222 22106 17458
rect 21318 5132 21554 5218
rect 21318 5068 21404 5132
rect 21404 5068 21468 5132
rect 21468 5068 21554 5132
rect 21318 4982 21554 5068
rect 23342 20092 23578 20178
rect 23342 20028 23428 20092
rect 23428 20028 23492 20092
rect 23492 20028 23578 20092
rect 23342 19942 23578 20028
rect 23342 17902 23578 18138
rect 22606 15182 22842 15418
rect 23342 12612 23578 12698
rect 23342 12548 23428 12612
rect 23428 12548 23492 12612
rect 23492 12548 23578 12612
rect 23342 12462 23578 12548
rect 22974 9892 23210 9978
rect 22974 9828 23060 9892
rect 23060 9828 23124 9892
rect 23124 9828 23210 9892
rect 22974 9742 23210 9828
rect 23894 10422 24130 10658
rect 23894 7022 24130 7258
rect 23894 5662 24130 5898
rect 23342 4452 23578 4538
rect 23342 4388 23428 4452
rect 23428 4388 23492 4452
rect 23492 4388 23578 4452
rect 23342 4302 23578 4388
rect 20398 2262 20634 2498
rect 16534 1582 16770 1818
rect 20398 1052 20634 1138
rect 20398 988 20484 1052
rect 20484 988 20548 1052
rect 20548 988 20634 1052
rect 20398 902 20634 988
<< metal5 >>
rect 6004 26298 26564 26340
rect 6004 26062 6046 26298
rect 6282 26062 26286 26298
rect 26522 26062 26564 26298
rect 6004 26020 26564 26062
rect 13916 25618 27116 25660
rect 13916 25382 13958 25618
rect 14194 25382 26838 25618
rect 27074 25382 27116 25618
rect 13916 25340 27116 25382
rect 18516 23578 22148 23620
rect 18516 23342 18558 23578
rect 18794 23342 21870 23578
rect 22106 23342 22148 23578
rect 18516 23300 22148 23342
rect 8948 22218 19572 22260
rect 8948 21982 8990 22218
rect 9226 21982 19294 22218
rect 19530 21982 19572 22218
rect 8948 21940 19572 21982
rect 7108 21538 21228 21580
rect 7108 21302 7150 21538
rect 7386 21302 20950 21538
rect 21186 21302 21228 21538
rect 7108 21260 21228 21302
rect 2508 20178 11108 20220
rect 2508 19942 2550 20178
rect 2786 19942 10830 20178
rect 11066 19942 11108 20178
rect 2508 19900 11108 19942
rect 13180 20178 23620 20220
rect 13180 19942 13222 20178
rect 13458 19942 23342 20178
rect 23578 19942 23620 20178
rect 13180 19900 23620 19942
rect 7476 19498 21412 19540
rect 7476 19262 7518 19498
rect 7754 19262 21134 19498
rect 21370 19262 21412 19498
rect 7476 19220 21412 19262
rect 8396 18138 23620 18180
rect 8396 17902 8438 18138
rect 8674 17902 23342 18138
rect 23578 17902 23620 18138
rect 8396 17860 23620 17902
rect 11340 17458 22148 17500
rect 11340 17222 11382 17458
rect 11618 17222 21870 17458
rect 22106 17222 22148 17458
rect 11340 17180 22148 17222
rect 1772 16778 12396 16820
rect 1772 16542 1814 16778
rect 2050 16542 12118 16778
rect 12354 16542 12396 16778
rect 1772 16500 12396 16542
rect 9500 15418 22884 15460
rect 9500 15182 9542 15418
rect 9778 15182 22606 15418
rect 22842 15182 22884 15418
rect 9500 15140 22884 15182
rect 8028 13378 19572 13420
rect 8028 13142 8070 13378
rect 8306 13142 19294 13378
rect 19530 13142 19572 13378
rect 8028 13100 19572 13142
rect 4900 12698 23620 12740
rect 4900 12462 4942 12698
rect 5178 12462 23342 12698
rect 23578 12462 23620 12698
rect 4900 12420 23620 12462
rect 4900 12018 19572 12060
rect 4900 11782 4942 12018
rect 5178 11782 19294 12018
rect 19530 11782 19572 12018
rect 4900 11740 19572 11782
rect 5268 10658 24172 10700
rect 5268 10422 5310 10658
rect 5546 10422 23894 10658
rect 24130 10422 24172 10658
rect 5268 10380 24172 10422
rect 14100 9978 23252 10020
rect 14100 9742 14142 9978
rect 14378 9742 22974 9978
rect 23210 9742 23252 9978
rect 14100 9700 23252 9742
rect 5268 9298 12028 9340
rect 5268 9062 5310 9298
rect 5546 9062 11750 9298
rect 11986 9062 12028 9298
rect 5268 9020 12028 9062
rect 3980 8618 16996 8660
rect 3980 8382 4022 8618
rect 4258 8382 16718 8618
rect 16954 8382 16996 8618
rect 3980 8340 16996 8382
rect 3796 7938 14788 7980
rect 3796 7702 3838 7938
rect 4074 7702 14510 7938
rect 14746 7702 14788 7938
rect 3796 7660 14788 7702
rect 8028 7258 24172 7300
rect 8028 7022 8070 7258
rect 8306 7022 23894 7258
rect 24130 7022 24172 7258
rect 8028 6980 24172 7022
rect 11708 6578 16996 6620
rect 11708 6342 11750 6578
rect 11986 6342 16718 6578
rect 16954 6342 16996 6578
rect 11708 6300 16996 6342
rect 5268 5898 24172 5940
rect 5268 5662 5310 5898
rect 5546 5662 16166 5898
rect 16402 5662 23894 5898
rect 24130 5662 24172 5898
rect 5268 5620 24172 5662
rect 12996 5218 21596 5260
rect 12996 4982 13038 5218
rect 13274 4982 21318 5218
rect 21554 4982 21596 5218
rect 12996 4940 21596 4982
rect 6556 4538 23620 4580
rect 6556 4302 6598 4538
rect 6834 4302 23342 4538
rect 23578 4302 23620 4538
rect 6556 4260 23620 4302
rect 3796 2498 20676 2540
rect 3796 2262 3838 2498
rect 4074 2262 20398 2498
rect 20634 2262 20676 2498
rect 3796 2220 20676 2262
rect 2140 1818 16812 1860
rect 2140 1582 2182 1818
rect 2418 1582 16534 1818
rect 16770 1582 16812 1818
rect 2140 1540 16812 1582
rect 3060 1138 20676 1180
rect 3060 902 3102 1138
rect 3338 902 20398 1138
rect 20634 902 20676 1138
rect 3060 860 20676 902
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_3_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_16 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_12
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_16
timestamp 1586364061
transform 1 0 2576 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_12
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A0
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_3.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 590 592
use scs8hd_conb_1  _046_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_3_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_49 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_45
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _107_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 10028 0 -1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_111 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_115
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 12696 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_130
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_4_
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_146
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_169
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_173
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_201
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_4_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_227
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_231
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_234
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_234
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_238
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_242
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_243
timestamp 1586364061
transform 1 0 23460 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__S
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__S
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l5_in_0_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_268
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A1
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_272
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A0
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_5_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__S
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_11
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_53
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_57
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_61
timestamp 1586364061
transform 1 0 6716 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9752 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_87
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_100
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_176
timestamp 1586364061
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_189
timestamp 1586364061
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_193
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l3_in_3_
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__S
timestamp 1586364061
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_241
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_247
timestamp 1586364061
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_262
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_266
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A1
timestamp 1586364061
transform 1 0 25760 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A0
timestamp 1586364061
transform 1 0 26128 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l4_in_1_
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A1
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A0
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_24
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_28
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12052 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_111
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_169
timestamp 1586364061
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_203
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_207
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_224
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_234
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l3_in_2_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_242
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_266
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_270
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l3_in_2_
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__S
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_4_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__S
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_21
timestamp 1586364061
transform 1 0 3036 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_2_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_69
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_112
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_116
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_3_
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_4_169
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_3_
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_2_
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23736 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_241
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_245
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_248
timestamp 1586364061
transform 1 0 23920 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_258
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_262
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_266
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_163
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_200
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 130 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21896 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 26312 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_268
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_272
timestamp 1586364061
transform 1 0 26128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_12
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__S
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l5_in_0_
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_44
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_48
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_54
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_55
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_82
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_90
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_102
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_2_
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 866 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_119
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_126
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_conb_1  _031_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_130
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_157
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 15364 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_161
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_159
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_4_
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_176
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_197
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_193
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19504 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21068 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_214
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_238
timestamp 1586364061
transform 1 0 23000 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_238
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_242
timestamp 1586364061
transform 1 0 23368 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23552 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23736 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_255
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 25116 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_267
timestamp 1586364061
transform 1 0 25668 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_272
timestamp 1586364061
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_268
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_271
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25852 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_276
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 26312 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A0
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__S
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_48
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_52
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_116
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_120
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_3_
timestamp 1586364061
transform 1 0 15364 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_147
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_168
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_191
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_195
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_241
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_245
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_258
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_262
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25392 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_266
timestamp 1586364061
transform 1 0 25576 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25760 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_270
timestamp 1586364061
transform 1 0 25944 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A1
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 1786 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_9
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_32
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_49
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_85
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_106
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _033_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_126
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_192
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 26128 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_270
timestamp 1586364061
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 314 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_7_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__S
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__S
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_6_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_114
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_171
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_179
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_191
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_195
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_207
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_222
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_245
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_249
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_262
timestamp 1586364061
transform 1 0 25208 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25392 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_266
timestamp 1586364061
transform 1 0 25576 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A0
timestamp 1586364061
transform 1 0 25760 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l3_in_3_
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_9
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_22
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_43
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_79
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_82
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_146
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_150
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_167
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_188
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_254
timestamp 1586364061
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 26128 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_266
timestamp 1586364061
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_270
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_274
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A0
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A1
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A1
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_76
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A1
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_33.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_114
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_184
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_32.mux_l1_in_3_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_257
timestamp 1586364061
transform 1 0 24748 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 25116 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_265
timestamp 1586364061
transform 1 0 25484 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_269
timestamp 1586364061
transform 1 0 25852 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__S
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A1
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_6_
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_48
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A0
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_2_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_75
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_85
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A0
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_3_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_32.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_115
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_111
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_133
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_3_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_146
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_150
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15364 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_164
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_185
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 18492 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18768 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_211
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_13_228
timestamp 1586364061
transform 1 0 22080 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_234
timestamp 1586364061
transform 1 0 22632 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_238
timestamp 1586364061
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23368 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_261
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_269
timestamp 1586364061
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_265
timestamp 1586364061
transform 1 0 25484 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_268
timestamp 1586364061
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_272
timestamp 1586364061
transform 1 0 26128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 26312 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_43
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A0
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_4_
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_162
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18492 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_198
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_215
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 590 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_268
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_272
timestamp 1586364061
transform 1 0 26128 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__S
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_51
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_116
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_158
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16192 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_162
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_183
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_209
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_228
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_241
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_262
timestamp 1586364061
transform 1 0 25208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_258
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__S
timestamp 1586364061
transform 1 0 25024 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_266
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25392 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_270
timestamp 1586364061
transform 1 0 25944 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25760 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use scs8hd_mux2_2  mux_left_track_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__S
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_9
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_13
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_30
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_88
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_116
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 406 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_3_
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_200
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_213
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_230
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A1
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_264
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_268
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_272
timestamp 1586364061
transform 1 0 26128 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l3_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l3_in_3_
timestamp 1586364061
transform 1 0 4232 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_43
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_conb_1  _029_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_96
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_100
timestamp 1586364061
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_148
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15824 0 -1 12512
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_179
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_183
timestamp 1586364061
transform 1 0 17940 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_187
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_203
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A1
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 20976 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21528 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_4.mux_l4_in_1_
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_250
timestamp 1586364061
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A0
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_267 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 866 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l4_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A1
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_38
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_4  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_42
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_4_
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 866 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_78
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_2_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8648 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_95
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_91
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_103
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_101
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_4_
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_149
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_153
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_157
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_24.mux_l4_in_0_
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_164
timestamp 1586364061
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l3_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16928 0 -1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_195
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_191
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A1
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_207
timestamp 1586364061
transform 1 0 20148 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_201
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19964 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 866 592
use scs8hd_conb_1  _032_
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_218
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_228
timestamp 1586364061
transform 1 0 22080 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_231
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 22632 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_253
timestamp 1586364061
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_257
timestamp 1586364061
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_265
timestamp 1586364061
transform 1 0 25484 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_266
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_274
timestamp 1586364061
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_270
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 26128 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 1786 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_29
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_56
timestamp 1586364061
transform 1 0 6256 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_17.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 1786 592
use scs8hd_conb_1  _030_
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_100
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_104
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_149
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_2_
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_209
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_213
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_226
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_3_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_266
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_270 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25944 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 1472 0 -1 14688
box -38 -48 1786 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_53
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_57
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_69
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__S
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_114
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_173
timestamp 1586364061
transform 1 0 17020 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17756 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_197
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_201
timestamp 1586364061
transform 1 0 19596 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 22632 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_228
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_232
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_236
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_22_240
timestamp 1586364061
transform 1 0 23184 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_260
timestamp 1586364061
transform 1 0 25024 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_264
timestamp 1586364061
transform 1 0 25392 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_272
timestamp 1586364061
transform 1 0 26128 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_5.mux_l5_in_0_
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A0
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_18
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A1
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__S
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_22
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_49
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_70
timestamp 1586364061
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A0
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_4_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A1
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_137
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_2_
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_157
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_3_
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_214
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_218
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_235
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_268
timestamp 1586364061
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_272
timestamp 1586364061
transform 1 0 26128 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_7_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__S
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_11
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_51
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_85
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_101
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_127
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_172
timestamp 1586364061
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_185
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21620 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_219
timestamp 1586364061
transform 1 0 21252 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24104 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23552 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 23920 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_242
timestamp 1586364061
transform 1 0 23368 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_246
timestamp 1586364061
transform 1 0 23736 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25116 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_263 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _063_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 1786 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_12
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_67
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_91
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_108
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_137
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_141
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_176
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_180
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_211
timestamp 1586364061
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_234
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_254
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 406 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_261
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_266
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_270
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_9
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_13
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_26
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_43
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_55
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_75
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_102
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_101
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_148
timestamp 1586364061
transform 1 0 14720 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_165
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_161
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_171
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _127_
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18952 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 18768 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_197
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_190
timestamp 1586364061
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_207
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_203
timestamp 1586364061
transform 1 0 19780 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_201
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20148 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_209
timestamp 1586364061
transform 1 0 20332 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_16.mux_l4_in_0_
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_27_224
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21528 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_238
timestamp 1586364061
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_234
timestamp 1586364061
transform 1 0 22632 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23368 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_254
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_255
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24748 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 24380 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_266
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 24932 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_270
timestamp 1586364061
transform 1 0 25944 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_conb_1  _028_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_10
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l4_in_0_
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A0
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_65
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9752 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_3_
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_103
timestamp 1586364061
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_120
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_137
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_2  _129_
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_161
timestamp 1586364061
transform 1 0 15916 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_165
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_2_
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_196
timestamp 1586364061
transform 1 0 19136 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 22264 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_228
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 24012 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_241
timestamp 1586364061
transform 1 0 23276 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_247
timestamp 1586364061
transform 1 0 23828 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_262
timestamp 1586364061
transform 1 0 25208 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_258
timestamp 1586364061
transform 1 0 24840 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 25024 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_266
timestamp 1586364061
transform 1 0 25576 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 25392 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_270
timestamp 1586364061
transform 1 0 25944 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25760 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_274
timestamp 1586364061
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 866 592
use scs8hd_buf_4  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 590 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_9
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_13
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_26
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_30
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A1
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _066_
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 130 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_162
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_166
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_201
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 22264 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 21896 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_224
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_228
timestamp 1586364061
transform 1 0 22080 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_254
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _083_
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 26128 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_270
timestamp 1586364061
transform 1 0 25944 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_274
timestamp 1586364061
transform 1 0 26312 0 1 17952
box -38 -48 314 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_10
timestamp 1586364061
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_29
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_5_
timestamp 1586364061
transform 1 0 6440 0 -1 19040
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__S
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_40
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_50
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_54
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_67
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_71
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_97
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_33.mux_l1_in_3_
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_120
timestamp 1586364061
transform 1 0 12144 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_124
timestamp 1586364061
transform 1 0 12512 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_137
timestamp 1586364061
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_2_
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_4_
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_180
timestamp 1586364061
transform 1 0 17664 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_197
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19412 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20148 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_201
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_205
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_209
timestamp 1586364061
transform 1 0 20332 0 -1 19040
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_2_
timestamp 1586364061
transform 1 0 22448 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 22264 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_228
timestamp 1586364061
transform 1 0 22080 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24012 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_241
timestamp 1586364061
transform 1 0 23276 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_247
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25024 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25392 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_258
timestamp 1586364061
transform 1 0 24840 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_262
timestamp 1586364061
transform 1 0 25208 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_266
timestamp 1586364061
transform 1 0 25576 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _064_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_70
timestamp 1586364061
transform 1 0 7544 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_111
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_115
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_119
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use scs8hd_buf_2  _131_
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_128
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_155
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_3_
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_172
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_176
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 20700 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 20148 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_205
timestamp 1586364061
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_236
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_254
timestamp 1586364061
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 25208 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 26128 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_258
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_266
timestamp 1586364061
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_270
timestamp 1586364061
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_274
timestamp 1586364061
transform 1 0 26312 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_8
timestamp 1586364061
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_12
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4324 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_29
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5888 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_48
timestamp 1586364061
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_71
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_75
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_79
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_25.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_106
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_110
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_122
timestamp 1586364061
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14536 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_148
timestamp 1586364061
transform 1 0 14720 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_157
timestamp 1586364061
transform 1 0 15548 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15732 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_161
timestamp 1586364061
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_184
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_188
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 21068 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_203
timestamp 1586364061
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_207
timestamp 1586364061
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_211
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21344 0 -1 20128
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_32_219
timestamp 1586364061
transform 1 0 21252 0 -1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_2_
timestamp 1586364061
transform 1 0 23828 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23644 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 23276 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_243
timestamp 1586364061
transform 1 0 23460 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_256
timestamp 1586364061
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_260
timestamp 1586364061
transform 1 0 25024 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25208 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_267
timestamp 1586364061
transform 1 0 25668 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 25392 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 25852 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_8
timestamp 1586364061
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_12
timestamp 1586364061
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_19
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_29
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_39
timestamp 1586364061
transform 1 0 4692 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_35
timestamp 1586364061
transform 1 0 4324 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A0
timestamp 1586364061
transform 1 0 4508 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_40
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_52
timestamp 1586364061
transform 1 0 5888 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 6624 0 -1 21216
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_67
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_79
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_87
timestamp 1586364061
transform 1 0 9108 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_83
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_84
timestamp 1586364061
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_80
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A0
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_97
timestamp 1586364061
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__S
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_33_101
timestamp 1586364061
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_116
timestamp 1586364061
transform 1 0 11776 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_112
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 11960 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 11592 0 -1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12512 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12328 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_120
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_133
timestamp 1586364061
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_137
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_146
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_buf_2  _123_
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14904 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_168
timestamp 1586364061
transform 1 0 16560 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_167
timestamp 1586364061
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_163
timestamp 1586364061
transform 1 0 16100 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16836 0 -1 21216
box -38 -48 866 592
use scs8hd_buf_2  _120_
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_186
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_180
timestamp 1586364061
transform 1 0 17664 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18400 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_197
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_190
timestamp 1586364061
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_207
timestamp 1586364061
transform 1 0 20148 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_201
timestamp 1586364061
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_205
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_201
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19412 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20148 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_211
timestamp 1586364061
transform 1 0 20516 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_218
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20332 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_228
timestamp 1586364061
transform 1 0 22080 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_224
timestamp 1586364061
transform 1 0 21712 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_222
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21896 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_3_
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_33_235
timestamp 1586364061
transform 1 0 22724 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 22264 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l4_in_0_
timestamp 1586364061
transform 1 0 22448 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_247
timestamp 1586364061
transform 1 0 23828 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_241
timestamp 1586364061
transform 1 0 23276 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23644 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_254
timestamp 1586364061
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24012 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_262
timestamp 1586364061
transform 1 0 25208 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_258
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_258
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25392 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_270
timestamp 1586364061
transform 1 0 25944 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_266
timestamp 1586364061
transform 1 0 25576 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_268
timestamp 1586364061
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25760 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_276
timestamp 1586364061
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_272
timestamp 1586364061
transform 1 0 26128 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 26128 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 26312 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_13
timestamp 1586364061
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_17
timestamp 1586364061
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3404 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_21
timestamp 1586364061
transform 1 0 3036 0 1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_35_36
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_40
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_43
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 1786 592
use scs8hd_buf_4  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_60
timestamp 1586364061
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_69
timestamp 1586364061
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_73
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A1
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_96
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A0
timestamp 1586364061
transform 1 0 10488 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_100
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_104
timestamp 1586364061
transform 1 0 10672 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_buf_2  _121_
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15088 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14720 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_142
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_146
timestamp 1586364061
transform 1 0 14536 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_150
timestamp 1586364061
transform 1 0 14904 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_158
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l3_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18768 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18584 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_188
timestamp 1586364061
transform 1 0 18400 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_217
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21252 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_228
timestamp 1586364061
transform 1 0 22080 0 1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_35_234
timestamp 1586364061
transform 1 0 22632 0 1 21216
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_240
timestamp 1586364061
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_254
timestamp 1586364061
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 25944 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 26312 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_258
timestamp 1586364061
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_268
timestamp 1586364061
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_272
timestamp 1586364061
transform 1 0 26128 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_276
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use scs8hd_buf_2  _060_
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 406 592
use scs8hd_buf_2  _065_
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 1932 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2300 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_7
timestamp 1586364061
transform 1 0 1748 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_11
timestamp 1586364061
transform 1 0 2116 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_19
timestamp 1586364061
transform 1 0 2852 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A1
timestamp 1586364061
transform 1 0 3036 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_29
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_6_
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 4876 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__S
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_40
timestamp 1586364061
transform 1 0 4784 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_50
timestamp 1586364061
transform 1 0 5704 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_54
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__S
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_67
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_73
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_7_
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 11592 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 11132 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_107
timestamp 1586364061
transform 1 0 10948 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_111
timestamp 1586364061
transform 1 0 11316 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_123
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_127
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_140
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_144
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16008 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_160
timestamp 1586364061
transform 1 0 15824 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_164
timestamp 1586364061
transform 1 0 16192 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19044 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 18492 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 18860 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_187
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_191
timestamp 1586364061
transform 1 0 18676 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_204
timestamp 1586364061
transform 1 0 19872 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_208
timestamp 1586364061
transform 1 0 20240 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_213
timestamp 1586364061
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 22448 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 21896 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22264 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_224
timestamp 1586364061
transform 1 0 21712 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_228
timestamp 1586364061
transform 1 0 22080 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 24012 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_241
timestamp 1586364061
transform 1 0 23276 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_247
timestamp 1586364061
transform 1 0 23828 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_262
timestamp 1586364061
transform 1 0 25208 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_258
timestamp 1586364061
transform 1 0 24840 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_266
timestamp 1586364061
transform 1 0 25576 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 25392 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_270
timestamp 1586364061
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25760 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_buf_2  _059_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_buf_2  _061_
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _067_
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 3036 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_23
timestamp 1586364061
transform 1 0 3220 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_36
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_3_
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_40
timestamp 1586364061
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l3_in_3_
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 7360 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_60
timestamp 1586364061
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_66
timestamp 1586364061
transform 1 0 7176 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_70
timestamp 1586364061
transform 1 0 7544 0 1 22304
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l3_in_2_
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__S
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__S
timestamp 1586364061
transform 1 0 8648 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_84
timestamp 1586364061
transform 1 0 8832 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_97
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_101
timestamp 1586364061
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13340 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 12604 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_127
timestamp 1586364061
transform 1 0 12788 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_152
timestamp 1586364061
transform 1 0 15088 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l4_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20516 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 20332 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19964 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_203
timestamp 1586364061
transform 1 0 19780 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_207
timestamp 1586364061
transform 1 0 20148 0 1 22304
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22080 0 1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 21528 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 21896 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_224
timestamp 1586364061
transform 1 0 21712 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_234
timestamp 1586364061
transform 1 0 22632 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_254
timestamp 1586364061
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 590 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25944 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_268
timestamp 1586364061
transform 1 0 25760 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_272
timestamp 1586364061
transform 1 0 26128 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_276
timestamp 1586364061
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use scs8hd_buf_2  _058_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_buf_2  _062_
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A1
timestamp 1586364061
transform 1 0 1932 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A0
timestamp 1586364061
transform 1 0 2300 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_11
timestamp 1586364061
transform 1 0 2116 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A0
timestamp 1586364061
transform 1 0 3036 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_38
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_2  _116_
timestamp 1586364061
transform 1 0 5336 0 -1 23392
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_4_
timestamp 1586364061
transform 1 0 6440 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4784 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5888 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_42
timestamp 1586364061
transform 1 0 4968 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_50
timestamp 1586364061
transform 1 0 5704 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_54
timestamp 1586364061
transform 1 0 6072 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l4_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__S
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_67
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_71
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_88
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11592 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11960 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_112
timestamp 1586364061
transform 1 0 11408 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_116
timestamp 1586364061
transform 1 0 11776 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_120
timestamp 1586364061
transform 1 0 12144 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_130
timestamp 1586364061
transform 1 0 13064 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_134
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_138
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use scs8hd_buf_4  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13892 0 -1 23392
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_149
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_2_
timestamp 1586364061
transform 1 0 16836 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 16652 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_167
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_3_
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_180
timestamp 1586364061
transform 1 0 17664 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_186
timestamp 1586364061
transform 1 0 18216 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_197
timestamp 1586364061
transform 1 0 19228 0 -1 23392
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__S
timestamp 1586364061
transform 1 0 20056 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20516 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_201
timestamp 1586364061
transform 1 0 19596 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_204
timestamp 1586364061
transform 1 0 19872 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_208
timestamp 1586364061
transform 1 0 20240 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 22724 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22448 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_224
timestamp 1586364061
transform 1 0 21712 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_228
timestamp 1586364061
transform 1 0 22080 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_234
timestamp 1586364061
transform 1 0 22632 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 24288 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23920 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_244
timestamp 1586364061
transform 1 0 23552 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_250
timestamp 1586364061
transform 1 0 24104 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25668 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_261
timestamp 1586364061
transform 1 0 25116 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_265
timestamp 1586364061
transform 1 0 25484 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_269
timestamp 1586364061
transform 1 0 25852 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_buf_2  _057_
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _056_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_decap_6  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_24
timestamp 1586364061
transform 1 0 3312 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_21
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_28
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_32
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3864 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_38
timestamp 1586364061
transform 1 0 4600 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_36
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_42
timestamp 1586364061
transform 1 0 4968 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4784 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5060 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_46
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_45
timestamp 1586364061
transform 1 0 5244 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5612 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _132_
timestamp 1586364061
transform 1 0 5612 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _135_
timestamp 1586364061
transform 1 0 5796 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_59
timestamp 1586364061
transform 1 0 6532 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_55
timestamp 1586364061
transform 1 0 6164 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 6348 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_67
timestamp 1586364061
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A1
timestamp 1586364061
transform 1 0 6716 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__S
timestamp 1586364061
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_5_
timestamp 1586364061
transform 1 0 7452 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _130_
timestamp 1586364061
transform 1 0 6900 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_71
timestamp 1586364061
transform 1 0 7636 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_78
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 7820 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_4_
timestamp 1586364061
transform 1 0 8004 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_88
timestamp 1586364061
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_97
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10580 0 -1 24480
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_109
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_113
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_127
timestamp 1586364061
transform 1 0 12788 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_122
timestamp 1586364061
transform 1 0 12328 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13156 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_148
timestamp 1586364061
transform 1 0 14720 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_144
timestamp 1586364061
transform 1 0 14352 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14536 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14168 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_152
timestamp 1586364061
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14904 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 15456 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_40_162
timestamp 1586364061
transform 1 0 16008 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_161
timestamp 1586364061
transform 1 0 15916 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16192 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_177
timestamp 1586364061
transform 1 0 17388 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_173
timestamp 1586364061
transform 1 0 17020 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17204 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17572 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 17756 0 -1 24480
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_3_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_198
timestamp 1586364061
transform 1 0 19320 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_194
timestamp 1586364061
transform 1 0 18952 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_198
timestamp 1586364061
transform 1 0 19320 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19136 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 18768 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A0
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_206
timestamp 1586364061
transform 1 0 20056 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_5_
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_210
timestamp 1586364061
transform 1 0 20424 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_215
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_211
timestamp 1586364061
transform 1 0 20516 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21068 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_228
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21252 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21252 0 1 23392
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21436 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_234
timestamp 1586364061
transform 1 0 22632 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_230
timestamp 1586364061
transform 1 0 22264 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_237
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_233
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22448 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 22816 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__S
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_238
timestamp 1586364061
transform 1 0 23000 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_241
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_6_
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_252
timestamp 1586364061
transform 1 0 24288 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_248
timestamp 1586364061
transform 1 0 23920 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 24472 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 24104 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23920 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 24656 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_261
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 25484 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_272
timestamp 1586364061
transform 1 0 26128 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_39_273
timestamp 1586364061
transform 1 0 26220 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 26036 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_260
timestamp 1586364061
transform 1 0 25024 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_42
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_46
timestamp 1586364061
transform 1 0 5336 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5520 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_54
timestamp 1586364061
transform 1 0 6072 0 1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_41_50
timestamp 1586364061
transform 1 0 5704 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A0
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _134_
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_66
timestamp 1586364061
transform 1 0 7176 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_70
timestamp 1586364061
transform 1 0 7544 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l5_in_0_
timestamp 1586364061
transform 1 0 9476 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__S
timestamp 1586364061
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_83
timestamp 1586364061
transform 1 0 8740 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_87
timestamp 1586364061
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _124_
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10948 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_100
timestamp 1586364061
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_104
timestamp 1586364061
transform 1 0 10672 0 1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_41_109
timestamp 1586364061
transform 1 0 11132 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 14720 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_146
timestamp 1586364061
transform 1 0 14536 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_150
timestamp 1586364061
transform 1 0 14904 0 1 24480
box -38 -48 314 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 16928 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16744 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_164
timestamp 1586364061
transform 1 0 16192 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_168
timestamp 1586364061
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _117_
timestamp 1586364061
transform 1 0 18860 0 1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 18400 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_179
timestamp 1586364061
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_41_190
timestamp 1586364061
transform 1 0 18584 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_197
timestamp 1586364061
transform 1 0 19228 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19964 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 19412 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 19780 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A1
timestamp 1586364061
transform 1 0 21068 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_201
timestamp 1586364061
transform 1 0 19596 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_214
timestamp 1586364061
transform 1 0 20792 0 1 24480
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_4_
timestamp 1586364061
transform 1 0 21620 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 21436 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A0
timestamp 1586364061
transform 1 0 22632 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__S
timestamp 1586364061
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_219
timestamp 1586364061
transform 1 0 21252 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_236
timestamp 1586364061
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_7_
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1586364061
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 24656 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_240
timestamp 1586364061
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_254
timestamp 1586364061
transform 1 0 24472 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 25208 0 1 24480
box -38 -48 406 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 25760 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_258
timestamp 1586364061
transform 1 0 24840 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_266
timestamp 1586364061
transform 1 0 25576 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_270
timestamp 1586364061
transform 1 0 25944 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_276
timestamp 1586364061
transform 1 0 26496 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _133_
timestamp 1586364061
transform 1 0 7452 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A0
timestamp 1586364061
transform 1 0 8372 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A1
timestamp 1586364061
transform 1 0 7268 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_73
timestamp 1586364061
transform 1 0 7820 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_77
timestamp 1586364061
transform 1 0 8188 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _125_
timestamp 1586364061
transform 1 0 9844 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _128_
timestamp 1586364061
transform 1 0 8556 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A1
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A1
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_85
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_89
timestamp 1586364061
transform 1 0 9292 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_99
timestamp 1586364061
transform 1 0 10212 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10948 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A0
timestamp 1586364061
transform 1 0 10396 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_103
timestamp 1586364061
transform 1 0 10580 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_116
timestamp 1586364061
transform 1 0 11776 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 13616 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_120
timestamp 1586364061
transform 1 0 12144 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_134
timestamp 1586364061
transform 1 0 13432 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_138
timestamp 1586364061
transform 1 0 13800 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _122_
timestamp 1586364061
transform 1 0 14260 0 -1 25568
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13984 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_142
timestamp 1586364061
transform 1 0 14168 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_147
timestamp 1586364061
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_151
timestamp 1586364061
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _119_
timestamp 1586364061
transform 1 0 17112 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_8  FILLER_42_165
timestamp 1586364061
transform 1 0 16284 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_173
timestamp 1586364061
transform 1 0 17020 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_178
timestamp 1586364061
transform 1 0 17480 0 -1 25568
box -38 -48 314 592
use scs8hd_buf_2  _118_
timestamp 1586364061
transform 1 0 18400 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_183
timestamp 1586364061
transform 1 0 17940 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_192
timestamp 1586364061
transform 1 0 18768 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _126_
timestamp 1586364061
transform 1 0 19504 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20056 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20424 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_204
timestamp 1586364061
transform 1 0 19872 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_208
timestamp 1586364061
transform 1 0 20240 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_212
timestamp 1586364061
transform 1 0 20608 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_216
timestamp 1586364061
transform 1 0 20976 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 21712 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 22816 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__S
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 21344 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_222
timestamp 1586364061
transform 1 0 21528 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_228
timestamp 1586364061
transform 1 0 22080 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_232
timestamp 1586364061
transform 1 0 22448 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A0
timestamp 1586364061
transform 1 0 23644 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_240
timestamp 1586364061
transform 1 0 23184 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_244
timestamp 1586364061
transform 1 0 23552 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_247
timestamp 1586364061
transform 1 0 23828 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_259
timestamp 1586364061
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_271
timestamp 1586364061
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1214 0 1270 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 1766 0 1822 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2226 0 2282 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 2778 0 2834 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 3882 0 3938 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 25502 0 25558 480 6 ccff_head
port 8 nsew default input
rlabel metal2 s 26054 0 26110 480 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 280 480 400 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 10208 480 10328 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 1504 480 1624 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 2184 480 2304 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 2864 480 2984 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 3544 480 3664 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 22856 480 22976 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 24896 480 25016 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 25576 480 25696 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 26256 480 26376 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 27520 4632 28000 4752 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 27520 10344 28000 10464 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 27520 10888 28000 11008 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 27520 11432 28000 11552 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 27520 11976 28000 12096 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 27520 5856 28000 5976 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 27520 6400 28000 6520 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 27520 7488 28000 7608 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 27520 8032 28000 8152 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 27520 8576 28000 8696 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 27520 9120 28000 9240 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 27520 21496 28000 21616 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 27520 22040 28000 22160 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 27520 22584 28000 22704 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 27520 23808 28000 23928 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 27520 24352 28000 24472 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 27520 24896 28000 25016 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 27520 25440 28000 25560 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 27520 25984 28000 26104 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 27520 16464 28000 16584 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 27520 17008 28000 17128 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 27520 17552 28000 17672 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 27520 18096 28000 18216 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 27520 18640 28000 18760 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 27520 19320 28000 19440 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 27520 19864 28000 19984 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 27520 20408 28000 20528 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 27520 20952 28000 21072 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 10690 0 10746 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 11242 0 11298 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 4894 0 4950 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 5446 0 5502 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 6458 0 6514 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 7010 0 7066 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 20166 0 20222 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 21270 0 21326 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 21822 0 21878 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 22282 0 22338 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 22834 0 22890 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 23386 0 23442 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 23938 0 23994 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 24398 0 24454 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 24950 0 25006 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal2 s 294 27520 350 28000 6 chany_top_in[0]
port 130 nsew default input
rlabel metal2 s 5814 27520 5870 28000 6 chany_top_in[10]
port 131 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[11]
port 132 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 chany_top_in[12]
port 133 nsew default input
rlabel metal2 s 7562 27520 7618 28000 6 chany_top_in[13]
port 134 nsew default input
rlabel metal2 s 8114 27520 8170 28000 6 chany_top_in[14]
port 135 nsew default input
rlabel metal2 s 8666 27520 8722 28000 6 chany_top_in[15]
port 136 nsew default input
rlabel metal2 s 9218 27520 9274 28000 6 chany_top_in[16]
port 137 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[17]
port 138 nsew default input
rlabel metal2 s 10322 27520 10378 28000 6 chany_top_in[18]
port 139 nsew default input
rlabel metal2 s 10874 27520 10930 28000 6 chany_top_in[19]
port 140 nsew default input
rlabel metal2 s 846 27520 902 28000 6 chany_top_in[1]
port 141 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 chany_top_in[2]
port 142 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 chany_top_in[3]
port 143 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 chany_top_in[4]
port 144 nsew default input
rlabel metal2 s 3054 27520 3110 28000 6 chany_top_in[5]
port 145 nsew default input
rlabel metal2 s 3606 27520 3662 28000 6 chany_top_in[6]
port 146 nsew default input
rlabel metal2 s 4158 27520 4214 28000 6 chany_top_in[7]
port 147 nsew default input
rlabel metal2 s 4710 27520 4766 28000 6 chany_top_in[8]
port 148 nsew default input
rlabel metal2 s 5262 27520 5318 28000 6 chany_top_in[9]
port 149 nsew default input
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[0]
port 150 nsew default tristate
rlabel metal2 s 21546 27520 21602 28000 6 chany_top_out[10]
port 151 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[11]
port 152 nsew default tristate
rlabel metal2 s 22650 27520 22706 28000 6 chany_top_out[12]
port 153 nsew default tristate
rlabel metal2 s 23202 27520 23258 28000 6 chany_top_out[13]
port 154 nsew default tristate
rlabel metal2 s 23754 27520 23810 28000 6 chany_top_out[14]
port 155 nsew default tristate
rlabel metal2 s 24306 27520 24362 28000 6 chany_top_out[15]
port 156 nsew default tristate
rlabel metal2 s 24858 27520 24914 28000 6 chany_top_out[16]
port 157 nsew default tristate
rlabel metal2 s 25410 27520 25466 28000 6 chany_top_out[17]
port 158 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[18]
port 159 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[19]
port 160 nsew default tristate
rlabel metal2 s 16486 27520 16542 28000 6 chany_top_out[1]
port 161 nsew default tristate
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_out[2]
port 162 nsew default tristate
rlabel metal2 s 17590 27520 17646 28000 6 chany_top_out[3]
port 163 nsew default tristate
rlabel metal2 s 18142 27520 18198 28000 6 chany_top_out[4]
port 164 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[5]
port 165 nsew default tristate
rlabel metal2 s 19246 27520 19302 28000 6 chany_top_out[6]
port 166 nsew default tristate
rlabel metal2 s 19798 27520 19854 28000 6 chany_top_out[7]
port 167 nsew default tristate
rlabel metal2 s 20350 27520 20406 28000 6 chany_top_out[8]
port 168 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[9]
port 169 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 left_top_grid_pin_42_
port 170 nsew default input
rlabel metal2 s 26514 0 26570 480 6 left_top_grid_pin_43_
port 171 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 left_top_grid_pin_44_
port 172 nsew default input
rlabel metal3 s 0 26936 480 27056 6 left_top_grid_pin_45_
port 173 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 left_top_grid_pin_46_
port 174 nsew default input
rlabel metal2 s 27066 0 27122 480 6 left_top_grid_pin_47_
port 175 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_48_
port 176 nsew default input
rlabel metal2 s 27618 0 27674 480 6 left_top_grid_pin_49_
port 177 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 prog_clk
port 178 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_top_grid_pin_42_
port 179 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_top_grid_pin_43_
port 180 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_top_grid_pin_44_
port 181 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_top_grid_pin_45_
port 182 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 right_top_grid_pin_46_
port 183 nsew default input
rlabel metal3 s 27520 3000 28000 3120 6 right_top_grid_pin_47_
port 184 nsew default input
rlabel metal3 s 27520 3544 28000 3664 6 right_top_grid_pin_48_
port 185 nsew default input
rlabel metal3 s 27520 4088 28000 4208 6 right_top_grid_pin_49_
port 186 nsew default input
rlabel metal2 s 11426 27520 11482 28000 6 top_left_grid_pin_34_
port 187 nsew default input
rlabel metal2 s 11978 27520 12034 28000 6 top_left_grid_pin_35_
port 188 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 top_left_grid_pin_36_
port 189 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 top_left_grid_pin_37_
port 190 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 top_left_grid_pin_38_
port 191 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 top_left_grid_pin_39_
port 192 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 top_left_grid_pin_40_
port 193 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 top_left_grid_pin_41_
port 194 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 195 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 196 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
