VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1178.580 BY 1266.000 ;
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 220.280 51.880 220.880 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1127.080 1026.760 1129.480 1027.360 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 102.640 51.880 103.240 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 338.600 51.880 339.200 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.270 1221.720 139.550 1224.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 604.330 44.120 604.610 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 634.230 44.120 634.510 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 664.130 44.120 664.410 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 694.030 44.120 694.310 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 723.930 44.120 724.210 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 754.290 44.120 754.570 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 456.240 51.880 456.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 810.520 51.880 811.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 319.130 1221.720 319.410 1224.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1127.080 240.000 1129.480 240.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1127.080 633.720 1129.480 634.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.290 44.120 64.570 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.190 44.120 94.470 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.090 44.120 124.370 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 153.990 44.120 154.270 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.890 44.120 184.170 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 214.250 44.120 214.530 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 498.990 1221.720 499.270 1224.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 784.190 44.120 784.470 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 814.090 44.120 814.370 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 843.990 44.120 844.270 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.350 44.120 874.630 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 904.250 44.120 904.530 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 934.150 44.120 934.430 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 574.560 51.880 575.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 928.160 51.880 928.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.310 1221.720 679.590 1224.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1127.080 371.240 1129.480 371.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1127.080 764.280 1129.480 764.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.150 44.120 244.430 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.050 44.120 274.330 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 303.950 44.120 304.230 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.310 44.120 334.590 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.210 44.120 364.490 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 394.110 44.120 394.390 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 859.170 1221.720 859.450 1224.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 964.050 44.120 964.330 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 993.950 44.120 994.230 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.310 44.120 1024.590 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1054.210 44.120 1054.490 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1084.110 44.120 1084.390 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1114.010 44.120 1114.290 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 692.200 51.880 692.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1046.480 51.880 1047.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1039.030 1221.720 1039.310 1224.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1127.080 502.480 1129.480 503.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1127.080 895.520 1129.480 896.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 424.010 44.120 424.290 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 453.910 44.120 454.190 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.270 44.120 484.550 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 514.170 44.120 514.450 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 544.070 44.120 544.350 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.970 44.120 574.250 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1127.080 109.440 1129.480 110.040 ;
    END
  END prog_clk
  PIN sc_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1164.120 51.880 1164.720 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1127.080 1158.000 1129.480 1158.600 ;
    END
  END sc_tail
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 1153.580 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 1178.580 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 105.000 89.765 1073.800 1185.075 ;
      LAYER met1 ;
        RECT 63.810 60.480 1114.310 1221.500 ;
      LAYER met2 ;
        RECT 63.830 1221.440 138.990 1221.720 ;
        RECT 139.830 1221.440 318.850 1221.720 ;
        RECT 319.690 1221.440 498.710 1221.720 ;
        RECT 499.550 1221.440 679.030 1221.720 ;
        RECT 679.870 1221.440 858.890 1221.720 ;
        RECT 859.730 1221.440 1038.750 1221.720 ;
        RECT 1039.590 1221.440 1114.280 1221.720 ;
        RECT 63.830 46.800 1114.280 1221.440 ;
        RECT 63.830 46.520 64.010 46.800 ;
        RECT 64.850 46.520 93.910 46.800 ;
        RECT 94.750 46.520 123.810 46.800 ;
        RECT 124.650 46.520 153.710 46.800 ;
        RECT 154.550 46.520 183.610 46.800 ;
        RECT 184.450 46.520 213.970 46.800 ;
        RECT 214.810 46.520 243.870 46.800 ;
        RECT 244.710 46.520 273.770 46.800 ;
        RECT 274.610 46.520 303.670 46.800 ;
        RECT 304.510 46.520 334.030 46.800 ;
        RECT 334.870 46.520 363.930 46.800 ;
        RECT 364.770 46.520 393.830 46.800 ;
        RECT 394.670 46.520 423.730 46.800 ;
        RECT 424.570 46.520 453.630 46.800 ;
        RECT 454.470 46.520 483.990 46.800 ;
        RECT 484.830 46.520 513.890 46.800 ;
        RECT 514.730 46.520 543.790 46.800 ;
        RECT 544.630 46.520 573.690 46.800 ;
        RECT 574.530 46.520 604.050 46.800 ;
        RECT 604.890 46.520 633.950 46.800 ;
        RECT 634.790 46.520 663.850 46.800 ;
        RECT 664.690 46.520 693.750 46.800 ;
        RECT 694.590 46.520 723.650 46.800 ;
        RECT 724.490 46.520 754.010 46.800 ;
        RECT 754.850 46.520 783.910 46.800 ;
        RECT 784.750 46.520 813.810 46.800 ;
        RECT 814.650 46.520 843.710 46.800 ;
        RECT 844.550 46.520 874.070 46.800 ;
        RECT 874.910 46.520 903.970 46.800 ;
        RECT 904.810 46.520 933.870 46.800 ;
        RECT 934.710 46.520 963.770 46.800 ;
        RECT 964.610 46.520 993.670 46.800 ;
        RECT 994.510 46.520 1024.030 46.800 ;
        RECT 1024.870 46.520 1053.930 46.800 ;
        RECT 1054.770 46.520 1083.830 46.800 ;
        RECT 1084.670 46.520 1113.730 46.800 ;
      LAYER met3 ;
        RECT 51.880 1165.120 1127.080 1182.945 ;
        RECT 52.280 1163.720 1127.080 1165.120 ;
        RECT 51.880 1159.000 1127.080 1163.720 ;
        RECT 51.880 1157.600 1126.680 1159.000 ;
        RECT 51.880 1047.480 1127.080 1157.600 ;
        RECT 52.280 1046.080 1127.080 1047.480 ;
        RECT 51.880 1027.760 1127.080 1046.080 ;
        RECT 51.880 1026.360 1126.680 1027.760 ;
        RECT 51.880 929.160 1127.080 1026.360 ;
        RECT 52.280 927.760 1127.080 929.160 ;
        RECT 51.880 896.520 1127.080 927.760 ;
        RECT 51.880 895.120 1126.680 896.520 ;
        RECT 51.880 811.520 1127.080 895.120 ;
        RECT 52.280 810.120 1127.080 811.520 ;
        RECT 51.880 765.280 1127.080 810.120 ;
        RECT 51.880 763.880 1126.680 765.280 ;
        RECT 51.880 693.200 1127.080 763.880 ;
        RECT 52.280 691.800 1127.080 693.200 ;
        RECT 51.880 634.720 1127.080 691.800 ;
        RECT 51.880 633.320 1126.680 634.720 ;
        RECT 51.880 575.560 1127.080 633.320 ;
        RECT 52.280 574.160 1127.080 575.560 ;
        RECT 51.880 503.480 1127.080 574.160 ;
        RECT 51.880 502.080 1126.680 503.480 ;
        RECT 51.880 457.240 1127.080 502.080 ;
        RECT 52.280 455.840 1127.080 457.240 ;
        RECT 51.880 372.240 1127.080 455.840 ;
        RECT 51.880 370.840 1126.680 372.240 ;
        RECT 51.880 339.600 1127.080 370.840 ;
        RECT 52.280 338.200 1127.080 339.600 ;
        RECT 51.880 241.000 1127.080 338.200 ;
        RECT 51.880 239.600 1126.680 241.000 ;
        RECT 51.880 221.280 1127.080 239.600 ;
        RECT 52.280 219.880 1127.080 221.280 ;
        RECT 51.880 110.440 1127.080 219.880 ;
        RECT 51.880 109.040 1126.680 110.440 ;
        RECT 51.880 103.640 1127.080 109.040 ;
        RECT 52.280 102.240 1127.080 103.640 ;
        RECT 51.880 85.095 1127.080 102.240 ;
      LAYER met4 ;
        RECT 0.000 0.000 1178.580 1266.000 ;
      LAYER met5 ;
        RECT 0.000 79.200 1178.580 1266.000 ;
  END
END fpga_core
END LIBRARY

