magic
tech EFS8A
magscale 1 2
timestamp 1602269361
<< locali >>
rect 16163 23137 16290 23171
rect 1443 22049 1478 22083
rect 6687 21029 6732 21063
rect 18279 20961 18314 20995
rect 12259 20009 12265 20043
rect 12259 19941 12293 20009
rect 22879 19873 22914 19907
rect 12759 19193 12804 19227
rect 8159 18785 8194 18819
rect 8401 18207 8435 18377
rect 14105 18275 14139 18377
rect 8435 18173 8562 18207
rect 8401 18124 8435 18173
rect 6463 17833 6469 17867
rect 6463 17765 6497 17833
rect 23949 17697 24110 17731
rect 23949 17527 23983 17697
rect 11299 17153 11437 17187
rect 22971 16609 23006 16643
rect 23983 16609 24018 16643
rect 3151 15895 3185 15963
rect 3151 15861 3157 15895
rect 17693 14943 17727 15113
rect 10051 14569 10057 14603
rect 13639 14569 13645 14603
rect 10051 14501 10085 14569
rect 13639 14501 13673 14569
rect 4077 14263 4111 14433
rect 12541 13855 12575 14025
rect 12541 13821 12655 13855
rect 20815 13719 20849 13787
rect 20815 13685 20821 13719
rect 18515 13481 18521 13515
rect 18515 13413 18549 13481
rect 12817 13175 12851 13413
rect 17083 13345 17118 13379
rect 14013 13175 14047 13345
rect 13823 12393 13829 12427
rect 25099 12393 25145 12427
rect 13823 12325 13857 12393
rect 22971 12257 23006 12291
rect 23983 12257 24018 12291
rect 8125 11543 8159 11849
rect 8619 11169 8654 11203
rect 11287 11169 11322 11203
rect 7481 9911 7515 10081
rect 15663 9129 15669 9163
rect 15663 9061 15697 9129
rect 24627 8993 24662 9027
rect 16991 8381 17026 8415
rect 4623 8279 4657 8347
rect 9631 8313 9676 8347
rect 15571 8279 15605 8347
rect 17325 8279 17359 8381
rect 18889 8279 18923 8517
rect 4623 8245 4629 8279
rect 15571 8245 15577 8279
rect 4623 8041 4629 8075
rect 11155 8041 11161 8075
rect 4623 7973 4657 8041
rect 11155 7973 11189 8041
rect 2455 7905 2582 7939
rect 2881 6817 3042 6851
rect 2881 6647 2915 6817
<< viali >>
rect 13553 24361 13587 24395
rect 5432 24225 5466 24259
rect 13369 24225 13403 24259
rect 5503 24021 5537 24055
rect 5825 23817 5859 23851
rect 13369 23817 13403 23851
rect 13645 23817 13679 23851
rect 18245 23817 18279 23851
rect 21465 23817 21499 23851
rect 5400 23613 5434 23647
rect 6193 23613 6227 23647
rect 13461 23613 13495 23647
rect 18061 23613 18095 23647
rect 18613 23613 18647 23647
rect 21281 23613 21315 23647
rect 21833 23613 21867 23647
rect 5503 23477 5537 23511
rect 14105 23477 14139 23511
rect 6837 23273 6871 23307
rect 13967 23273 14001 23307
rect 16359 23273 16393 23307
rect 13896 23137 13930 23171
rect 16129 23137 16163 23171
rect 24660 23137 24694 23171
rect 13645 22933 13679 22967
rect 24731 22933 24765 22967
rect 1869 22729 1903 22763
rect 14565 22729 14599 22763
rect 20131 22729 20165 22763
rect 25513 22729 25547 22763
rect 6653 22661 6687 22695
rect 25145 22661 25179 22695
rect 6929 22593 6963 22627
rect 1460 22525 1494 22559
rect 8744 22525 8778 22559
rect 13553 22525 13587 22559
rect 14013 22525 14047 22559
rect 20060 22525 20094 22559
rect 24660 22525 24694 22559
rect 1547 22457 1581 22491
rect 7021 22457 7055 22491
rect 7573 22457 7607 22491
rect 14289 22457 14323 22491
rect 8815 22389 8849 22423
rect 9229 22389 9263 22423
rect 13369 22389 13403 22423
rect 16221 22389 16255 22423
rect 20453 22389 20487 22423
rect 24731 22389 24765 22423
rect 8953 22185 8987 22219
rect 21465 22185 21499 22219
rect 6469 22117 6503 22151
rect 7021 22117 7055 22151
rect 8033 22117 8067 22151
rect 12449 22117 12483 22151
rect 13001 22117 13035 22151
rect 16865 22117 16899 22151
rect 1409 22049 1443 22083
rect 9756 22049 9790 22083
rect 18312 22049 18346 22083
rect 21992 22049 22026 22083
rect 23556 22049 23590 22083
rect 24660 22049 24694 22083
rect 6377 21981 6411 22015
rect 7941 21981 7975 22015
rect 8585 21981 8619 22015
rect 12909 21981 12943 22015
rect 13553 21981 13587 22015
rect 15577 21981 15611 22015
rect 16773 21981 16807 22015
rect 17049 21981 17083 22015
rect 20913 21981 20947 22015
rect 23627 21913 23661 21947
rect 1547 21845 1581 21879
rect 9827 21845 9861 21879
rect 14473 21845 14507 21879
rect 18383 21845 18417 21879
rect 22063 21845 22097 21879
rect 24731 21845 24765 21879
rect 1593 21641 1627 21675
rect 5549 21641 5583 21675
rect 8309 21641 8343 21675
rect 10241 21641 10275 21675
rect 15945 21641 15979 21675
rect 22385 21641 22419 21675
rect 23949 21641 23983 21675
rect 24685 21641 24719 21675
rect 8033 21573 8067 21607
rect 9781 21573 9815 21607
rect 8585 21505 8619 21539
rect 12541 21505 12575 21539
rect 12909 21505 12943 21539
rect 16497 21505 16531 21539
rect 16773 21505 16807 21539
rect 19165 21505 19199 21539
rect 21465 21505 21499 21539
rect 21741 21505 21775 21539
rect 10057 21437 10091 21471
rect 10609 21437 10643 21471
rect 14381 21437 14415 21471
rect 14473 21437 14507 21471
rect 14933 21437 14967 21471
rect 17877 21437 17911 21471
rect 18061 21437 18095 21471
rect 18521 21437 18555 21471
rect 19660 21437 19694 21471
rect 20085 21437 20119 21471
rect 6561 21369 6595 21403
rect 7021 21369 7055 21403
rect 7113 21369 7147 21403
rect 7665 21369 7699 21403
rect 8677 21369 8711 21403
rect 9229 21369 9263 21403
rect 12633 21369 12667 21403
rect 15209 21369 15243 21403
rect 16589 21369 16623 21403
rect 18797 21369 18831 21403
rect 21557 21369 21591 21403
rect 5917 21301 5951 21335
rect 6285 21301 6319 21335
rect 12265 21301 12299 21335
rect 13461 21301 13495 21335
rect 16221 21301 16255 21335
rect 17417 21301 17451 21335
rect 19763 21301 19797 21335
rect 21281 21301 21315 21335
rect 8723 21097 8757 21131
rect 15439 21097 15473 21131
rect 16497 21097 16531 21131
rect 19073 21097 19107 21131
rect 22201 21097 22235 21131
rect 6653 21029 6687 21063
rect 11989 21029 12023 21063
rect 12173 21029 12207 21063
rect 12265 21029 12299 21063
rect 13093 21029 13127 21063
rect 13829 21029 13863 21063
rect 16773 21029 16807 21063
rect 19441 21029 19475 21063
rect 21189 21029 21223 21063
rect 21281 21029 21315 21063
rect 22845 21029 22879 21063
rect 5400 20961 5434 20995
rect 5503 20961 5537 20995
rect 8620 20961 8654 20995
rect 10701 20961 10735 20995
rect 11069 20961 11103 20995
rect 15336 20961 15370 20995
rect 18245 20961 18279 20995
rect 24660 20961 24694 20995
rect 6377 20893 6411 20927
rect 11253 20893 11287 20927
rect 12817 20893 12851 20927
rect 13737 20893 13771 20927
rect 16681 20893 16715 20927
rect 17325 20893 17359 20927
rect 19349 20893 19383 20927
rect 21465 20893 21499 20927
rect 22753 20893 22787 20927
rect 23029 20893 23063 20927
rect 14289 20825 14323 20859
rect 18383 20825 18417 20859
rect 19901 20825 19935 20859
rect 5273 20757 5307 20791
rect 6193 20757 6227 20791
rect 7297 20757 7331 20791
rect 7941 20757 7975 20791
rect 15761 20757 15795 20791
rect 18061 20757 18095 20791
rect 18705 20757 18739 20791
rect 24731 20757 24765 20791
rect 1593 20553 1627 20587
rect 8401 20553 8435 20587
rect 13369 20553 13403 20587
rect 13645 20553 13679 20587
rect 14013 20553 14047 20587
rect 15025 20553 15059 20587
rect 17095 20553 17129 20587
rect 21465 20553 21499 20587
rect 23397 20553 23431 20587
rect 25145 20553 25179 20587
rect 25513 20553 25547 20587
rect 7757 20485 7791 20519
rect 16129 20485 16163 20519
rect 23029 20485 23063 20519
rect 4169 20417 4203 20451
rect 5917 20417 5951 20451
rect 8953 20417 8987 20451
rect 15209 20417 15243 20451
rect 16681 20417 16715 20451
rect 18705 20417 18739 20451
rect 20545 20417 20579 20451
rect 20821 20417 20855 20451
rect 22109 20417 22143 20451
rect 22385 20417 22419 20451
rect 1409 20349 1443 20383
rect 5089 20349 5123 20383
rect 5181 20349 5215 20383
rect 5641 20349 5675 20383
rect 6837 20349 6871 20383
rect 8033 20349 8067 20383
rect 9873 20349 9907 20383
rect 10241 20349 10275 20383
rect 11069 20349 11103 20383
rect 11253 20349 11287 20383
rect 11805 20349 11839 20383
rect 12449 20349 12483 20383
rect 14248 20349 14282 20383
rect 14657 20349 14691 20383
rect 17024 20349 17058 20383
rect 17417 20349 17451 20383
rect 19625 20349 19659 20383
rect 24660 20349 24694 20383
rect 6653 20281 6687 20315
rect 7199 20281 7233 20315
rect 8677 20281 8711 20315
rect 8769 20281 8803 20315
rect 11529 20281 11563 20315
rect 12811 20281 12845 20315
rect 14335 20281 14369 20315
rect 15571 20281 15605 20315
rect 19026 20281 19060 20315
rect 20361 20281 20395 20315
rect 20637 20281 20671 20315
rect 21925 20281 21959 20315
rect 22201 20281 22235 20315
rect 2053 20213 2087 20247
rect 6285 20213 6319 20247
rect 10609 20213 10643 20247
rect 12265 20213 12299 20247
rect 18245 20213 18279 20247
rect 19993 20213 20027 20247
rect 24731 20213 24765 20247
rect 1593 20009 1627 20043
rect 7665 20009 7699 20043
rect 8585 20009 8619 20043
rect 8953 20009 8987 20043
rect 12265 20009 12299 20043
rect 12817 20009 12851 20043
rect 13553 20009 13587 20043
rect 15117 20009 15151 20043
rect 16865 20009 16899 20043
rect 19533 20009 19567 20043
rect 19901 20009 19935 20043
rect 20545 20009 20579 20043
rect 23995 20009 24029 20043
rect 6187 19941 6221 19975
rect 7481 19941 7515 19975
rect 13829 19941 13863 19975
rect 14381 19941 14415 19975
rect 15622 19941 15656 19975
rect 16589 19941 16623 19975
rect 17233 19941 17267 19975
rect 18934 19941 18968 19975
rect 21189 19941 21223 19975
rect 21465 19941 21499 19975
rect 1409 19873 1443 19907
rect 4880 19873 4914 19907
rect 7113 19873 7147 19907
rect 7849 19873 7883 19907
rect 8033 19873 8067 19907
rect 10333 19873 10367 19907
rect 10885 19873 10919 19907
rect 22017 19873 22051 19907
rect 22845 19873 22879 19907
rect 23924 19873 23958 19907
rect 5825 19805 5859 19839
rect 11069 19805 11103 19839
rect 11897 19805 11931 19839
rect 13737 19805 13771 19839
rect 15301 19805 15335 19839
rect 17141 19805 17175 19839
rect 17601 19805 17635 19839
rect 18613 19805 18647 19839
rect 21373 19805 21407 19839
rect 5273 19737 5307 19771
rect 6745 19737 6779 19771
rect 11437 19737 11471 19771
rect 3617 19669 3651 19703
rect 4951 19669 4985 19703
rect 5641 19669 5675 19703
rect 13093 19669 13127 19703
rect 16221 19669 16255 19703
rect 22983 19669 23017 19703
rect 2651 19465 2685 19499
rect 4905 19465 4939 19499
rect 10333 19465 10367 19499
rect 15301 19465 15335 19499
rect 15669 19465 15703 19499
rect 17049 19465 17083 19499
rect 17877 19465 17911 19499
rect 20637 19465 20671 19499
rect 22109 19465 22143 19499
rect 9965 19397 9999 19431
rect 5917 19329 5951 19363
rect 6561 19329 6595 19363
rect 7389 19329 7423 19363
rect 7849 19329 7883 19363
rect 9229 19329 9263 19363
rect 11529 19329 11563 19363
rect 13645 19329 13679 19363
rect 14565 19329 14599 19363
rect 15945 19329 15979 19363
rect 18613 19329 18647 19363
rect 20269 19329 20303 19363
rect 21189 19329 21223 19363
rect 1409 19261 1443 19295
rect 2580 19261 2614 19295
rect 2973 19261 3007 19295
rect 3617 19261 3651 19295
rect 3709 19261 3743 19295
rect 3893 19261 3927 19295
rect 5181 19261 5215 19295
rect 5641 19261 5675 19295
rect 7113 19261 7147 19295
rect 10793 19261 10827 19295
rect 11345 19261 11379 19295
rect 12449 19261 12483 19295
rect 13369 19261 13403 19295
rect 14013 19261 14047 19295
rect 18889 19261 18923 19295
rect 4353 19193 4387 19227
rect 7481 19193 7515 19227
rect 8953 19193 8987 19227
rect 9045 19193 9079 19227
rect 12725 19193 12759 19227
rect 14289 19193 14323 19227
rect 14381 19193 14415 19227
rect 16037 19193 16071 19227
rect 16589 19193 16623 19227
rect 19210 19193 19244 19227
rect 21281 19193 21315 19227
rect 21833 19193 21867 19227
rect 1593 19125 1627 19159
rect 1961 19125 1995 19159
rect 3433 19125 3467 19159
rect 6285 19125 6319 19159
rect 8309 19125 8343 19159
rect 8769 19125 8803 19159
rect 11897 19125 11931 19159
rect 12173 19125 12207 19159
rect 17509 19125 17543 19159
rect 18245 19125 18279 19159
rect 19809 19125 19843 19159
rect 21005 19125 21039 19159
rect 22845 19125 22879 19159
rect 23949 19125 23983 19159
rect 1685 18921 1719 18955
rect 7573 18921 7607 18955
rect 8953 18921 8987 18955
rect 11897 18921 11931 18955
rect 13001 18921 13035 18955
rect 13645 18921 13679 18955
rect 14013 18921 14047 18955
rect 18889 18921 18923 18955
rect 6698 18853 6732 18887
rect 11253 18853 11287 18887
rect 12443 18853 12477 18887
rect 14657 18853 14691 18887
rect 15945 18853 15979 18887
rect 16497 18853 16531 18887
rect 18429 18853 18463 18887
rect 19441 18853 19475 18887
rect 19993 18853 20027 18887
rect 21557 18853 21591 18887
rect 23121 18853 23155 18887
rect 2973 18785 3007 18819
rect 4905 18785 4939 18819
rect 5273 18785 5307 18819
rect 7297 18785 7331 18819
rect 8125 18785 8159 18819
rect 10793 18785 10827 18819
rect 11069 18785 11103 18819
rect 14264 18785 14298 18819
rect 17693 18785 17727 18819
rect 18153 18785 18187 18819
rect 5549 18717 5583 18751
rect 6193 18717 6227 18751
rect 6377 18717 6411 18751
rect 10425 18717 10459 18751
rect 12081 18717 12115 18751
rect 15853 18717 15887 18751
rect 19349 18717 19383 18751
rect 21465 18717 21499 18751
rect 23029 18717 23063 18751
rect 23305 18717 23339 18751
rect 14335 18649 14369 18683
rect 15025 18649 15059 18683
rect 22017 18649 22051 18683
rect 2697 18581 2731 18615
rect 3709 18581 3743 18615
rect 8263 18581 8297 18615
rect 15577 18581 15611 18615
rect 21189 18581 21223 18615
rect 8401 18377 8435 18411
rect 8631 18377 8665 18411
rect 11483 18377 11517 18411
rect 14105 18377 14139 18411
rect 14289 18377 14323 18411
rect 15945 18377 15979 18411
rect 16313 18377 16347 18411
rect 18199 18377 18233 18411
rect 19073 18377 19107 18411
rect 21925 18377 21959 18411
rect 23029 18377 23063 18411
rect 4077 18309 4111 18343
rect 3433 18241 3467 18275
rect 5273 18241 5307 18275
rect 5917 18241 5951 18275
rect 7021 18241 7055 18275
rect 11161 18309 11195 18343
rect 20545 18309 20579 18343
rect 9781 18241 9815 18275
rect 13829 18241 13863 18275
rect 14105 18241 14139 18275
rect 8401 18173 8435 18207
rect 8953 18173 8987 18207
rect 10425 18173 10459 18207
rect 11412 18173 11446 18207
rect 12449 18173 12483 18207
rect 13001 18173 13035 18207
rect 16681 18173 16715 18207
rect 16865 18173 16899 18207
rect 18128 18173 18162 18207
rect 19257 18173 19291 18207
rect 21005 18173 21039 18207
rect 23397 18173 23431 18207
rect 23673 18173 23707 18207
rect 24133 18173 24167 18207
rect 3157 18105 3191 18139
rect 3249 18105 3283 18139
rect 4537 18105 4571 18139
rect 5365 18105 5399 18139
rect 7113 18105 7147 18139
rect 7665 18105 7699 18139
rect 9597 18105 9631 18139
rect 9873 18105 9907 18139
rect 10793 18105 10827 18139
rect 14933 18105 14967 18139
rect 15025 18105 15059 18139
rect 15577 18105 15611 18139
rect 17693 18105 17727 18139
rect 19578 18105 19612 18139
rect 20821 18105 20855 18139
rect 21326 18105 21360 18139
rect 2053 18037 2087 18071
rect 2605 18037 2639 18071
rect 2973 18037 3007 18071
rect 4905 18037 4939 18071
rect 6469 18037 6503 18071
rect 8125 18037 8159 18071
rect 12173 18037 12207 18071
rect 12541 18037 12575 18071
rect 13461 18037 13495 18071
rect 14657 18037 14691 18071
rect 16497 18037 16531 18071
rect 18613 18037 18647 18071
rect 20177 18037 20211 18071
rect 22201 18037 22235 18071
rect 22661 18037 22695 18071
rect 23765 18037 23799 18071
rect 1547 17833 1581 17867
rect 5273 17833 5307 17867
rect 6469 17833 6503 17867
rect 7021 17833 7055 17867
rect 7297 17833 7331 17867
rect 7757 17833 7791 17867
rect 9965 17833 9999 17867
rect 11437 17833 11471 17867
rect 13001 17833 13035 17867
rect 14381 17833 14415 17867
rect 14933 17833 14967 17867
rect 16405 17833 16439 17867
rect 18981 17833 19015 17867
rect 20729 17833 20763 17867
rect 22569 17833 22603 17867
rect 25191 17833 25225 17867
rect 2513 17765 2547 17799
rect 2605 17765 2639 17799
rect 3157 17765 3191 17799
rect 4261 17765 4295 17799
rect 8033 17765 8067 17799
rect 8585 17765 8619 17799
rect 10241 17765 10275 17799
rect 11805 17765 11839 17799
rect 12725 17765 12759 17799
rect 13823 17765 13857 17799
rect 15485 17765 15519 17799
rect 18245 17765 18279 17799
rect 21097 17765 21131 17799
rect 1476 17697 1510 17731
rect 13461 17697 13495 17731
rect 17509 17697 17543 17731
rect 17969 17697 18003 17731
rect 18521 17697 18555 17731
rect 19073 17697 19107 17731
rect 19533 17697 19567 17731
rect 22477 17697 22511 17731
rect 22937 17697 22971 17731
rect 23673 17697 23707 17731
rect 25120 17697 25154 17731
rect 1961 17629 1995 17663
rect 4169 17629 4203 17663
rect 4445 17629 4479 17663
rect 6101 17629 6135 17663
rect 7941 17629 7975 17663
rect 10149 17629 10183 17663
rect 11713 17629 11747 17663
rect 11989 17629 12023 17663
rect 15393 17629 15427 17663
rect 15669 17629 15703 17663
rect 19625 17629 19659 17663
rect 21005 17629 21039 17663
rect 10701 17561 10735 17595
rect 20177 17561 20211 17595
rect 21557 17561 21591 17595
rect 24179 17629 24213 17663
rect 3433 17493 3467 17527
rect 5549 17493 5583 17527
rect 6009 17493 6043 17527
rect 16773 17493 16807 17527
rect 21925 17493 21959 17527
rect 23949 17493 23983 17527
rect 2421 17289 2455 17323
rect 3801 17289 3835 17323
rect 4077 17289 4111 17323
rect 7757 17289 7791 17323
rect 8033 17289 8067 17323
rect 11069 17289 11103 17323
rect 15485 17289 15519 17323
rect 15761 17289 15795 17323
rect 17509 17289 17543 17323
rect 17785 17289 17819 17323
rect 19073 17289 19107 17323
rect 22845 17289 22879 17323
rect 24041 17289 24075 17323
rect 25513 17289 25547 17323
rect 1547 17221 1581 17255
rect 10333 17221 10367 17255
rect 11989 17221 12023 17255
rect 14105 17221 14139 17255
rect 14473 17221 14507 17255
rect 20545 17221 20579 17255
rect 4537 17153 4571 17187
rect 11437 17153 11471 17187
rect 12817 17153 12851 17187
rect 14565 17153 14599 17187
rect 16405 17153 16439 17187
rect 19625 17153 19659 17187
rect 21741 17153 21775 17187
rect 1444 17085 1478 17119
rect 1869 17085 1903 17119
rect 2881 17085 2915 17119
rect 5089 17085 5123 17119
rect 5457 17085 5491 17119
rect 5733 17085 5767 17119
rect 5917 17085 5951 17119
rect 6837 17085 6871 17119
rect 9413 17085 9447 17119
rect 10609 17085 10643 17119
rect 11228 17085 11262 17119
rect 11621 17085 11655 17119
rect 18061 17085 18095 17119
rect 18521 17085 18555 17119
rect 22477 17085 22511 17119
rect 24660 17085 24694 17119
rect 3202 17017 3236 17051
rect 7158 17017 7192 17051
rect 9229 17017 9263 17051
rect 9775 17017 9809 17051
rect 12725 17017 12759 17051
rect 13179 17017 13213 17051
rect 14886 17017 14920 17051
rect 16474 17017 16508 17051
rect 17049 17017 17083 17051
rect 18797 17017 18831 17051
rect 19946 17017 19980 17051
rect 21005 17017 21039 17051
rect 21465 17017 21499 17051
rect 21557 17017 21591 17051
rect 2789 16949 2823 16983
rect 6193 16949 6227 16983
rect 6561 16949 6595 16983
rect 8401 16949 8435 16983
rect 13737 16949 13771 16983
rect 16221 16949 16255 16983
rect 19441 16949 19475 16983
rect 24731 16949 24765 16983
rect 25145 16949 25179 16983
rect 2237 16745 2271 16779
rect 5917 16745 5951 16779
rect 6837 16745 6871 16779
rect 10609 16745 10643 16779
rect 14657 16745 14691 16779
rect 18061 16745 18095 16779
rect 19073 16745 19107 16779
rect 20269 16745 20303 16779
rect 20729 16745 20763 16779
rect 24087 16745 24121 16779
rect 2605 16677 2639 16711
rect 3157 16677 3191 16711
rect 4077 16677 4111 16711
rect 8769 16677 8803 16711
rect 9413 16677 9447 16711
rect 10051 16677 10085 16711
rect 13553 16677 13587 16711
rect 13829 16677 13863 16711
rect 14381 16677 14415 16711
rect 15663 16677 15697 16711
rect 17233 16677 17267 16711
rect 19441 16677 19475 16711
rect 19993 16677 20027 16711
rect 21097 16677 21131 16711
rect 21557 16677 21591 16711
rect 1476 16609 1510 16643
rect 4169 16609 4203 16643
rect 5641 16609 5675 16643
rect 6101 16609 6135 16643
rect 8309 16609 8343 16643
rect 8493 16609 8527 16643
rect 12081 16609 12115 16643
rect 12357 16609 12391 16643
rect 22937 16609 22971 16643
rect 23949 16609 23983 16643
rect 2513 16541 2547 16575
rect 9045 16541 9079 16575
rect 9689 16541 9723 16575
rect 12817 16541 12851 16575
rect 13737 16541 13771 16575
rect 15301 16541 15335 16575
rect 17141 16541 17175 16575
rect 19349 16541 19383 16575
rect 21465 16541 21499 16575
rect 1547 16473 1581 16507
rect 12173 16473 12207 16507
rect 15117 16473 15151 16507
rect 17693 16473 17727 16507
rect 22017 16473 22051 16507
rect 1961 16405 1995 16439
rect 3433 16405 3467 16439
rect 5181 16405 5215 16439
rect 11345 16405 11379 16439
rect 11621 16405 11655 16439
rect 16221 16405 16255 16439
rect 16497 16405 16531 16439
rect 18429 16405 18463 16439
rect 23075 16405 23109 16439
rect 1685 16201 1719 16235
rect 1915 16201 1949 16235
rect 3709 16201 3743 16235
rect 4077 16201 4111 16235
rect 4721 16201 4755 16235
rect 6193 16201 6227 16235
rect 8769 16201 8803 16235
rect 12173 16201 12207 16235
rect 15439 16201 15473 16235
rect 20177 16201 20211 16235
rect 21649 16201 21683 16235
rect 22385 16201 22419 16235
rect 23029 16201 23063 16235
rect 23949 16201 23983 16235
rect 7573 16133 7607 16167
rect 15117 16133 15151 16167
rect 16129 16133 16163 16167
rect 18889 16133 18923 16167
rect 5917 16065 5951 16099
rect 8401 16065 8435 16099
rect 9965 16065 9999 16099
rect 11529 16065 11563 16099
rect 13645 16065 13679 16099
rect 14565 16065 14599 16099
rect 17049 16065 17083 16099
rect 17785 16065 17819 16099
rect 18521 16065 18555 16099
rect 20729 16065 20763 16099
rect 1812 15997 1846 16031
rect 2237 15997 2271 16031
rect 2789 15997 2823 16031
rect 7849 15997 7883 16031
rect 8125 15997 8159 16031
rect 10609 15997 10643 16031
rect 11069 15997 11103 16031
rect 11253 15997 11287 16031
rect 14289 15997 14323 16031
rect 15368 15997 15402 16031
rect 15853 15997 15887 16031
rect 18981 15997 19015 16031
rect 19901 15997 19935 16031
rect 5273 15929 5307 15963
rect 5365 15929 5399 15963
rect 9321 15929 9355 15963
rect 9413 15929 9447 15963
rect 13737 15929 13771 15963
rect 16405 15929 16439 15963
rect 16497 15929 16531 15963
rect 19302 15929 19336 15963
rect 20545 15929 20579 15963
rect 21050 15929 21084 15963
rect 22477 15929 22511 15963
rect 2697 15861 2731 15895
rect 3157 15861 3191 15895
rect 4997 15861 5031 15895
rect 7205 15861 7239 15895
rect 9137 15861 9171 15895
rect 10241 15861 10275 15895
rect 12449 15861 12483 15895
rect 12909 15861 12943 15895
rect 13461 15861 13495 15895
rect 17325 15861 17359 15895
rect 22017 15861 22051 15895
rect 1961 15657 1995 15691
rect 6009 15657 6043 15691
rect 9505 15657 9539 15691
rect 10885 15657 10919 15691
rect 13277 15657 13311 15691
rect 13829 15657 13863 15691
rect 14289 15657 14323 15691
rect 19901 15657 19935 15691
rect 24777 15657 24811 15691
rect 3157 15589 3191 15623
rect 7665 15589 7699 15623
rect 9781 15589 9815 15623
rect 9873 15589 9907 15623
rect 11437 15589 11471 15623
rect 11989 15589 12023 15623
rect 15761 15589 15795 15623
rect 21189 15589 21223 15623
rect 21281 15589 21315 15623
rect 2421 15521 2455 15555
rect 2697 15521 2731 15555
rect 5457 15521 5491 15555
rect 6469 15521 6503 15555
rect 6745 15521 6779 15555
rect 8033 15521 8067 15555
rect 8493 15521 8527 15555
rect 12725 15521 12759 15555
rect 12817 15521 12851 15555
rect 13093 15521 13127 15555
rect 17785 15521 17819 15555
rect 18245 15521 18279 15555
rect 19349 15521 19383 15555
rect 22661 15521 22695 15555
rect 22937 15521 22971 15555
rect 24593 15521 24627 15555
rect 2329 15453 2363 15487
rect 4905 15453 4939 15487
rect 7205 15453 7239 15487
rect 8769 15453 8803 15487
rect 10057 15453 10091 15487
rect 11345 15453 11379 15487
rect 15669 15453 15703 15487
rect 18521 15453 18555 15487
rect 21557 15453 21591 15487
rect 23121 15453 23155 15487
rect 2513 15385 2547 15419
rect 6285 15385 6319 15419
rect 6561 15385 6595 15419
rect 12909 15385 12943 15419
rect 16221 15385 16255 15419
rect 22753 15385 22787 15419
rect 3433 15317 3467 15351
rect 9045 15317 9079 15351
rect 12265 15317 12299 15351
rect 16681 15317 16715 15351
rect 18981 15317 19015 15351
rect 20453 15317 20487 15351
rect 22201 15317 22235 15351
rect 1777 15113 1811 15147
rect 9597 15113 9631 15147
rect 11345 15113 11379 15147
rect 14197 15113 14231 15147
rect 16313 15113 16347 15147
rect 17693 15113 17727 15147
rect 17785 15113 17819 15147
rect 21373 15113 21407 15147
rect 21741 15113 21775 15147
rect 11069 15045 11103 15079
rect 11713 15045 11747 15079
rect 15577 15045 15611 15079
rect 2145 14977 2179 15011
rect 2513 14977 2547 15011
rect 8401 14977 8435 15011
rect 17141 14977 17175 15011
rect 22569 15045 22603 15079
rect 20453 14977 20487 15011
rect 22017 14977 22051 15011
rect 23811 14977 23845 15011
rect 2881 14909 2915 14943
rect 3341 14909 3375 14943
rect 3617 14909 3651 14943
rect 3985 14909 4019 14943
rect 4997 14909 5031 14943
rect 5641 14909 5675 14943
rect 6101 14909 6135 14943
rect 6469 14909 6503 14943
rect 6929 14909 6963 14943
rect 10149 14909 10183 14943
rect 12265 14909 12299 14943
rect 13277 14909 13311 14943
rect 13553 14909 13587 14943
rect 13829 14909 13863 14943
rect 14657 14909 14691 14943
rect 16497 14909 16531 14943
rect 16865 14909 16899 14943
rect 17693 14909 17727 14943
rect 18061 14909 18095 14943
rect 18521 14909 18555 14943
rect 19073 14909 19107 14943
rect 23724 14909 23758 14943
rect 24593 14909 24627 14943
rect 5089 14841 5123 14875
rect 6837 14841 6871 14875
rect 8309 14841 8343 14875
rect 8763 14841 8797 14875
rect 10057 14841 10091 14875
rect 10511 14841 10545 14875
rect 14473 14841 14507 14875
rect 14978 14841 15012 14875
rect 18797 14841 18831 14875
rect 20545 14841 20579 14875
rect 21097 14841 21131 14875
rect 22109 14841 22143 14875
rect 2697 14773 2731 14807
rect 4629 14773 4663 14807
rect 7849 14773 7883 14807
rect 9321 14773 9355 14807
rect 12909 14773 12943 14807
rect 15853 14773 15887 14807
rect 17509 14773 17543 14807
rect 20269 14773 20303 14807
rect 22937 14773 22971 14807
rect 23305 14773 23339 14807
rect 24225 14773 24259 14807
rect 2329 14569 2363 14603
rect 5181 14569 5215 14603
rect 7067 14569 7101 14603
rect 9413 14569 9447 14603
rect 10057 14569 10091 14603
rect 10609 14569 10643 14603
rect 12909 14569 12943 14603
rect 13645 14569 13679 14603
rect 14657 14569 14691 14603
rect 15117 14569 15151 14603
rect 18797 14569 18831 14603
rect 19901 14569 19935 14603
rect 20453 14569 20487 14603
rect 21925 14569 21959 14603
rect 1961 14501 1995 14535
rect 10885 14501 10919 14535
rect 11621 14501 11655 14535
rect 15761 14501 15795 14535
rect 19302 14501 19336 14535
rect 21097 14501 21131 14535
rect 22661 14501 22695 14535
rect 2421 14433 2455 14467
rect 2697 14433 2731 14467
rect 3801 14433 3835 14467
rect 4077 14433 4111 14467
rect 5365 14433 5399 14467
rect 5641 14433 5675 14467
rect 6996 14433 7030 14467
rect 8033 14433 8067 14467
rect 8493 14433 8527 14467
rect 11253 14433 11287 14467
rect 17417 14433 17451 14467
rect 17877 14433 17911 14467
rect 18429 14433 18463 14467
rect 18981 14433 19015 14467
rect 1409 14365 1443 14399
rect 3157 14365 3191 14399
rect 2513 14297 2547 14331
rect 3525 14297 3559 14331
rect 6101 14365 6135 14399
rect 8769 14365 8803 14399
rect 9689 14365 9723 14399
rect 11529 14365 11563 14399
rect 11989 14365 12023 14399
rect 12541 14365 12575 14399
rect 13277 14365 13311 14399
rect 15669 14365 15703 14399
rect 16313 14365 16347 14399
rect 18153 14365 18187 14399
rect 21005 14365 21039 14399
rect 21281 14365 21315 14399
rect 22569 14365 22603 14399
rect 22845 14365 22879 14399
rect 5457 14297 5491 14331
rect 6469 14297 6503 14331
rect 4077 14229 4111 14263
rect 4261 14229 4295 14263
rect 4905 14229 4939 14263
rect 7389 14229 7423 14263
rect 9045 14229 9079 14263
rect 14197 14229 14231 14263
rect 16589 14229 16623 14263
rect 8033 14025 8067 14059
rect 9597 14025 9631 14059
rect 11437 14025 11471 14059
rect 12265 14025 12299 14059
rect 12541 14025 12575 14059
rect 13737 14025 13771 14059
rect 14473 14025 14507 14059
rect 15945 14025 15979 14059
rect 17417 14025 17451 14059
rect 17785 14025 17819 14059
rect 19625 14025 19659 14059
rect 21649 14025 21683 14059
rect 22753 14025 22787 14059
rect 23029 14025 23063 14059
rect 2145 13957 2179 13991
rect 5273 13957 5307 13991
rect 5641 13889 5675 13923
rect 7113 13889 7147 13923
rect 7757 13889 7791 13923
rect 8677 13889 8711 13923
rect 10333 13889 10367 13923
rect 10517 13889 10551 13923
rect 11161 13889 11195 13923
rect 14013 13957 14047 13991
rect 15669 13957 15703 13991
rect 19901 13957 19935 13991
rect 20269 13957 20303 13991
rect 13369 13889 13403 13923
rect 15301 13889 15335 13923
rect 16497 13889 16531 13923
rect 18705 13889 18739 13923
rect 20453 13889 20487 13923
rect 1409 13821 1443 13855
rect 3157 13821 3191 13855
rect 3617 13821 3651 13855
rect 3709 13821 3743 13855
rect 4261 13821 4295 13855
rect 5181 13821 5215 13855
rect 5457 13821 5491 13855
rect 7021 13821 7055 13855
rect 7297 13821 7331 13855
rect 12725 13821 12759 13855
rect 12909 13821 12943 13855
rect 22268 13821 22302 13855
rect 23724 13821 23758 13855
rect 24133 13821 24167 13855
rect 2421 13753 2455 13787
rect 4629 13753 4663 13787
rect 8585 13753 8619 13787
rect 9039 13753 9073 13787
rect 10609 13753 10643 13787
rect 14657 13753 14691 13787
rect 14749 13753 14783 13787
rect 16221 13753 16255 13787
rect 16313 13753 16347 13787
rect 19026 13753 19060 13787
rect 23811 13753 23845 13787
rect 1593 13685 1627 13719
rect 2973 13685 3007 13719
rect 4997 13685 5031 13719
rect 6193 13685 6227 13719
rect 6653 13685 6687 13719
rect 9965 13685 9999 13719
rect 11897 13685 11931 13719
rect 18521 13685 18555 13719
rect 20821 13685 20855 13719
rect 21373 13685 21407 13719
rect 22109 13685 22143 13719
rect 22339 13685 22373 13719
rect 1685 13481 1719 13515
rect 9505 13481 9539 13515
rect 13185 13481 13219 13515
rect 15117 13481 15151 13515
rect 16497 13481 16531 13515
rect 18521 13481 18555 13515
rect 19349 13481 19383 13515
rect 20177 13481 20211 13515
rect 20453 13481 20487 13515
rect 24179 13481 24213 13515
rect 2599 13413 2633 13447
rect 4261 13413 4295 13447
rect 10701 13413 10735 13447
rect 11713 13413 11747 13447
rect 12817 13413 12851 13447
rect 15669 13413 15703 13447
rect 19809 13413 19843 13447
rect 21097 13413 21131 13447
rect 22661 13413 22695 13447
rect 3157 13345 3191 13379
rect 5641 13345 5675 13379
rect 5733 13345 5767 13379
rect 5917 13345 5951 13379
rect 7849 13345 7883 13379
rect 8309 13345 8343 13379
rect 8861 13345 8895 13379
rect 10149 13345 10183 13379
rect 2237 13277 2271 13311
rect 4169 13277 4203 13311
rect 4445 13277 4479 13311
rect 6377 13277 6411 13311
rect 8401 13277 8435 13311
rect 11621 13277 11655 13311
rect 11897 13277 11931 13311
rect 7021 13209 7055 13243
rect 13277 13345 13311 13379
rect 13645 13345 13679 13379
rect 14013 13345 14047 13379
rect 17049 13345 17083 13379
rect 24108 13345 24142 13379
rect 15577 13277 15611 13311
rect 15853 13277 15887 13311
rect 18153 13277 18187 13311
rect 21005 13277 21039 13311
rect 22569 13277 22603 13311
rect 22845 13277 22879 13311
rect 14657 13209 14691 13243
rect 17187 13209 17221 13243
rect 21557 13209 21591 13243
rect 2145 13141 2179 13175
rect 3433 13141 3467 13175
rect 3893 13141 3927 13175
rect 5181 13141 5215 13175
rect 6745 13141 6779 13175
rect 7389 13141 7423 13175
rect 10977 13141 11011 13175
rect 11345 13141 11379 13175
rect 12633 13141 12667 13175
rect 12817 13141 12851 13175
rect 13001 13141 13035 13175
rect 14013 13141 14047 13175
rect 14197 13141 14231 13175
rect 19073 13141 19107 13175
rect 3157 12937 3191 12971
rect 5457 12937 5491 12971
rect 7849 12937 7883 12971
rect 11805 12937 11839 12971
rect 14381 12937 14415 12971
rect 16635 12937 16669 12971
rect 20729 12937 20763 12971
rect 21097 12937 21131 12971
rect 22569 12937 22603 12971
rect 24133 12937 24167 12971
rect 24777 12937 24811 12971
rect 2789 12869 2823 12903
rect 8309 12869 8343 12903
rect 16037 12869 16071 12903
rect 18429 12869 18463 12903
rect 1777 12801 1811 12835
rect 2421 12801 2455 12835
rect 5779 12801 5813 12835
rect 6929 12801 6963 12835
rect 7205 12801 7239 12835
rect 9045 12801 9079 12835
rect 11529 12801 11563 12835
rect 15301 12801 15335 12835
rect 19441 12801 19475 12835
rect 20085 12801 20119 12835
rect 3249 12733 3283 12767
rect 3709 12733 3743 12767
rect 4261 12733 4295 12767
rect 4445 12733 4479 12767
rect 5181 12733 5215 12767
rect 5692 12733 5726 12767
rect 8401 12733 8435 12767
rect 8861 12733 8895 12767
rect 12541 12733 12575 12767
rect 13185 12733 13219 12767
rect 13369 12733 13403 12767
rect 13737 12733 13771 12767
rect 16405 12733 16439 12767
rect 16532 12733 16566 12767
rect 18245 12733 18279 12767
rect 24593 12733 24627 12767
rect 25145 12733 25179 12767
rect 1869 12665 1903 12699
rect 6469 12665 6503 12699
rect 7021 12665 7055 12699
rect 10885 12665 10919 12699
rect 10977 12665 11011 12699
rect 14013 12665 14047 12699
rect 15025 12665 15059 12699
rect 15117 12665 15151 12699
rect 19533 12665 19567 12699
rect 21281 12665 21315 12699
rect 21373 12665 21407 12699
rect 21925 12665 21959 12699
rect 3525 12597 3559 12631
rect 6101 12597 6135 12631
rect 10057 12597 10091 12631
rect 10701 12597 10735 12631
rect 12173 12597 12207 12631
rect 14749 12597 14783 12631
rect 17049 12597 17083 12631
rect 17877 12597 17911 12631
rect 18797 12597 18831 12631
rect 19257 12597 19291 12631
rect 22845 12597 22879 12631
rect 3341 12393 3375 12427
rect 3709 12393 3743 12427
rect 4997 12393 5031 12427
rect 6929 12393 6963 12427
rect 8125 12393 8159 12427
rect 8493 12393 8527 12427
rect 8723 12393 8757 12427
rect 11161 12393 11195 12427
rect 12909 12393 12943 12427
rect 13829 12393 13863 12427
rect 15025 12393 15059 12427
rect 16681 12393 16715 12427
rect 18797 12393 18831 12427
rect 21833 12393 21867 12427
rect 22063 12393 22097 12427
rect 25145 12393 25179 12427
rect 6469 12325 6503 12359
rect 7205 12325 7239 12359
rect 10603 12325 10637 12359
rect 12173 12325 12207 12359
rect 15485 12325 15519 12359
rect 17325 12325 17359 12359
rect 18337 12325 18371 12359
rect 24087 12325 24121 12359
rect 1777 12257 1811 12291
rect 2053 12257 2087 12291
rect 2697 12257 2731 12291
rect 4721 12257 4755 12291
rect 5181 12257 5215 12291
rect 5549 12257 5583 12291
rect 5917 12257 5951 12291
rect 8620 12257 8654 12291
rect 12265 12257 12299 12291
rect 14381 12257 14415 12291
rect 18981 12257 19015 12291
rect 19257 12257 19291 12291
rect 21992 12257 22026 12291
rect 22937 12257 22971 12291
rect 23949 12257 23983 12291
rect 25028 12257 25062 12291
rect 4537 12189 4571 12223
rect 7113 12189 7147 12223
rect 10241 12189 10275 12223
rect 13461 12189 13495 12223
rect 15393 12189 15427 12223
rect 15669 12189 15703 12223
rect 17233 12189 17267 12223
rect 17877 12189 17911 12223
rect 20913 12189 20947 12223
rect 7665 12121 7699 12155
rect 11529 12121 11563 12155
rect 12449 12121 12483 12155
rect 21465 12121 21499 12155
rect 23075 12121 23109 12155
rect 9965 12053 9999 12087
rect 13369 12053 13403 12087
rect 16405 12053 16439 12087
rect 19809 12053 19843 12087
rect 2145 11849 2179 11883
rect 4077 11849 4111 11883
rect 6193 11849 6227 11883
rect 8125 11849 8159 11883
rect 8953 11849 8987 11883
rect 12725 11849 12759 11883
rect 15025 11849 15059 11883
rect 15669 11849 15703 11883
rect 19073 11849 19107 11883
rect 19441 11849 19475 11883
rect 23949 11849 23983 11883
rect 3801 11781 3835 11815
rect 1869 11713 1903 11747
rect 2421 11713 2455 11747
rect 4997 11713 5031 11747
rect 6653 11713 6687 11747
rect 6837 11713 6871 11747
rect 2329 11645 2363 11679
rect 2605 11645 2639 11679
rect 3893 11645 3927 11679
rect 5917 11645 5951 11679
rect 7021 11645 7055 11679
rect 7941 11645 7975 11679
rect 3065 11577 3099 11611
rect 5359 11577 5393 11611
rect 12173 11781 12207 11815
rect 14657 11781 14691 11815
rect 16957 11781 16991 11815
rect 17417 11781 17451 11815
rect 24777 11781 24811 11815
rect 8539 11713 8573 11747
rect 11345 11713 11379 11747
rect 15209 11713 15243 11747
rect 18797 11713 18831 11747
rect 25513 11713 25547 11747
rect 8436 11645 8470 11679
rect 9505 11645 9539 11679
rect 10241 11645 10275 11679
rect 10517 11645 10551 11679
rect 10701 11645 10735 11679
rect 12909 11645 12943 11679
rect 13553 11645 13587 11679
rect 13829 11645 13863 11679
rect 14105 11645 14139 11679
rect 20361 11645 20395 11679
rect 21189 11645 21223 11679
rect 21373 11645 21407 11679
rect 24593 11645 24627 11679
rect 25145 11645 25179 11679
rect 8309 11577 8343 11611
rect 10977 11577 11011 11611
rect 14381 11577 14415 11611
rect 16405 11577 16439 11611
rect 16497 11577 16531 11611
rect 18153 11577 18187 11611
rect 18245 11577 18279 11611
rect 21281 11577 21315 11611
rect 3433 11509 3467 11543
rect 4813 11509 4847 11543
rect 8125 11509 8159 11543
rect 9413 11509 9447 11543
rect 11805 11509 11839 11543
rect 16221 11509 16255 11543
rect 17877 11509 17911 11543
rect 20177 11509 20211 11543
rect 22293 11509 22327 11543
rect 23029 11509 23063 11543
rect 1685 11305 1719 11339
rect 2145 11305 2179 11339
rect 3525 11305 3559 11339
rect 3893 11305 3927 11339
rect 5181 11305 5215 11339
rect 6745 11305 6779 11339
rect 7849 11305 7883 11339
rect 11391 11305 11425 11339
rect 12173 11305 12207 11339
rect 12541 11305 12575 11339
rect 15485 11305 15519 11339
rect 17555 11305 17589 11339
rect 19625 11305 19659 11339
rect 4077 11237 4111 11271
rect 5963 11237 5997 11271
rect 9873 11237 9907 11271
rect 11069 11237 11103 11271
rect 15990 11237 16024 11271
rect 19026 11237 19060 11271
rect 21097 11237 21131 11271
rect 2421 11169 2455 11203
rect 2513 11169 2547 11203
rect 2697 11169 2731 11203
rect 4261 11169 4295 11203
rect 5876 11169 5910 11203
rect 7481 11169 7515 11203
rect 8585 11169 8619 11203
rect 11253 11169 11287 11203
rect 12725 11169 12759 11203
rect 13185 11169 13219 11203
rect 13553 11169 13587 11203
rect 14105 11169 14139 11203
rect 15669 11169 15703 11203
rect 16589 11169 16623 11203
rect 17484 11169 17518 11203
rect 22544 11169 22578 11203
rect 3157 11101 3191 11135
rect 8723 11101 8757 11135
rect 9781 11101 9815 11135
rect 10057 11101 10091 11135
rect 14197 11101 14231 11135
rect 18705 11101 18739 11135
rect 21005 11101 21039 11135
rect 21557 11033 21591 11067
rect 5549 10965 5583 10999
rect 7113 10965 7147 10999
rect 9321 10965 9355 10999
rect 10793 10965 10827 10999
rect 11805 10965 11839 10999
rect 17141 10965 17175 10999
rect 18061 10965 18095 10999
rect 22615 10965 22649 10999
rect 2237 10761 2271 10795
rect 3433 10761 3467 10795
rect 5457 10761 5491 10795
rect 5917 10761 5951 10795
rect 9137 10761 9171 10795
rect 10241 10761 10275 10795
rect 10609 10761 10643 10795
rect 14473 10761 14507 10795
rect 14841 10761 14875 10795
rect 20269 10761 20303 10795
rect 21465 10761 21499 10795
rect 22845 10761 22879 10795
rect 8677 10693 8711 10727
rect 14105 10693 14139 10727
rect 17785 10693 17819 10727
rect 21097 10693 21131 10727
rect 22155 10693 22189 10727
rect 2513 10625 2547 10659
rect 3157 10625 3191 10659
rect 6653 10625 6687 10659
rect 9965 10625 9999 10659
rect 10885 10625 10919 10659
rect 11161 10625 11195 10659
rect 16957 10625 16991 10659
rect 18613 10625 18647 10659
rect 20545 10625 20579 10659
rect 2421 10557 2455 10591
rect 2697 10557 2731 10591
rect 4077 10557 4111 10591
rect 5089 10557 5123 10591
rect 6837 10557 6871 10591
rect 8033 10557 8067 10591
rect 12725 10557 12759 10591
rect 13185 10557 13219 10591
rect 13645 10557 13679 10591
rect 13921 10557 13955 10591
rect 15025 10557 15059 10591
rect 15945 10557 15979 10591
rect 17509 10557 17543 10591
rect 22084 10557 22118 10591
rect 22477 10557 22511 10591
rect 1961 10489 1995 10523
rect 4445 10489 4479 10523
rect 6285 10489 6319 10523
rect 7199 10489 7233 10523
rect 9321 10489 9355 10523
rect 9422 10489 9456 10523
rect 10977 10489 11011 10523
rect 11897 10489 11931 10523
rect 12265 10489 12299 10523
rect 15346 10489 15380 10523
rect 16221 10489 16255 10523
rect 18429 10489 18463 10523
rect 18934 10489 18968 10523
rect 20637 10489 20671 10523
rect 21833 10489 21867 10523
rect 7757 10421 7791 10455
rect 19533 10421 19567 10455
rect 2789 10217 2823 10251
rect 3249 10217 3283 10251
rect 4537 10217 4571 10251
rect 6929 10217 6963 10251
rect 9137 10217 9171 10251
rect 11575 10217 11609 10251
rect 12081 10217 12115 10251
rect 12449 10217 12483 10251
rect 15669 10217 15703 10251
rect 16037 10217 16071 10251
rect 18797 10217 18831 10251
rect 19165 10217 19199 10251
rect 20545 10217 20579 10251
rect 23719 10217 23753 10251
rect 24777 10217 24811 10251
rect 2145 10149 2179 10183
rect 3801 10149 3835 10183
rect 8033 10149 8067 10183
rect 9505 10149 9539 10183
rect 10057 10149 10091 10183
rect 10609 10149 10643 10183
rect 14381 10149 14415 10183
rect 15025 10149 15059 10183
rect 16405 10149 16439 10183
rect 16957 10149 16991 10183
rect 17785 10149 17819 10183
rect 21097 10149 21131 10183
rect 1501 10081 1535 10115
rect 5825 10081 5859 10115
rect 6285 10081 6319 10115
rect 6377 10081 6411 10115
rect 6929 10081 6963 10115
rect 7481 10081 7515 10115
rect 10885 10081 10919 10115
rect 11504 10081 11538 10115
rect 12909 10081 12943 10115
rect 13645 10081 13679 10115
rect 13829 10081 13863 10115
rect 14105 10081 14139 10115
rect 17877 10081 17911 10115
rect 19660 10081 19694 10115
rect 23616 10081 23650 10115
rect 24593 10081 24627 10115
rect 7941 10013 7975 10047
rect 8217 10013 8251 10047
rect 9965 10013 9999 10047
rect 16313 10013 16347 10047
rect 21005 10013 21039 10047
rect 21281 10013 21315 10047
rect 7665 9945 7699 9979
rect 2421 9877 2455 9911
rect 7389 9877 7423 9911
rect 7481 9877 7515 9911
rect 11345 9877 11379 9911
rect 12725 9877 12759 9911
rect 19763 9877 19797 9911
rect 1869 9673 1903 9707
rect 2421 9673 2455 9707
rect 3249 9673 3283 9707
rect 5641 9673 5675 9707
rect 13277 9673 13311 9707
rect 13645 9673 13679 9707
rect 16589 9673 16623 9707
rect 17509 9673 17543 9707
rect 23857 9673 23891 9707
rect 24777 9673 24811 9707
rect 25145 9673 25179 9707
rect 6009 9605 6043 9639
rect 6653 9605 6687 9639
rect 16957 9605 16991 9639
rect 20545 9605 20579 9639
rect 9597 9537 9631 9571
rect 12909 9537 12943 9571
rect 14657 9537 14691 9571
rect 15577 9537 15611 9571
rect 19349 9537 19383 9571
rect 19993 9537 20027 9571
rect 21005 9537 21039 9571
rect 21465 9537 21499 9571
rect 2053 9469 2087 9503
rect 3617 9469 3651 9503
rect 3985 9469 4019 9503
rect 4445 9469 4479 9503
rect 4721 9469 4755 9503
rect 5089 9469 5123 9503
rect 7113 9469 7147 9503
rect 7573 9469 7607 9503
rect 7849 9469 7883 9503
rect 8217 9469 8251 9503
rect 9229 9469 9263 9503
rect 10333 9469 10367 9503
rect 10609 9469 10643 9503
rect 10885 9469 10919 9503
rect 11437 9469 11471 9503
rect 11897 9469 11931 9503
rect 14565 9469 14599 9503
rect 14933 9469 14967 9503
rect 21557 9469 21591 9503
rect 24593 9469 24627 9503
rect 8585 9401 8619 9435
rect 12173 9401 12207 9435
rect 15669 9401 15703 9435
rect 16221 9401 16255 9435
rect 18153 9401 18187 9435
rect 18245 9401 18279 9435
rect 18797 9401 18831 9435
rect 20085 9401 20119 9435
rect 21281 9401 21315 9435
rect 3801 9333 3835 9367
rect 6929 9333 6963 9367
rect 9965 9333 9999 9367
rect 11253 9333 11287 9367
rect 12449 9333 12483 9367
rect 15393 9333 15427 9367
rect 17785 9333 17819 9367
rect 19625 9333 19659 9367
rect 24409 9333 24443 9367
rect 2329 9129 2363 9163
rect 3801 9129 3835 9163
rect 4169 9129 4203 9163
rect 6285 9129 6319 9163
rect 8401 9129 8435 9163
rect 8723 9129 8757 9163
rect 9413 9129 9447 9163
rect 9781 9129 9815 9163
rect 12357 9129 12391 9163
rect 12817 9129 12851 9163
rect 15669 9129 15703 9163
rect 16221 9129 16255 9163
rect 19993 9129 20027 9163
rect 23719 9129 23753 9163
rect 3157 9061 3191 9095
rect 7158 9061 7192 9095
rect 8033 9061 8067 9095
rect 17233 9061 17267 9095
rect 18705 9061 18739 9095
rect 18797 9061 18831 9095
rect 1476 8993 1510 9027
rect 3065 8993 3099 9027
rect 4261 8993 4295 9027
rect 4629 8993 4663 9027
rect 4905 8993 4939 9027
rect 5273 8993 5307 9027
rect 6837 8993 6871 9027
rect 8652 8993 8686 9027
rect 9965 8993 9999 9027
rect 10149 8993 10183 9027
rect 10701 8993 10735 9027
rect 10977 8993 11011 9027
rect 12909 8993 12943 9027
rect 13369 8993 13403 9027
rect 13737 8993 13771 9027
rect 14197 8993 14231 9027
rect 23648 8993 23682 9027
rect 24593 8993 24627 9027
rect 5917 8925 5951 8959
rect 14381 8925 14415 8959
rect 15301 8925 15335 8959
rect 17141 8925 17175 8959
rect 17417 8925 17451 8959
rect 18429 8925 18463 8959
rect 18981 8925 19015 8959
rect 1869 8857 1903 8891
rect 21189 8857 21223 8891
rect 24731 8857 24765 8891
rect 1547 8789 1581 8823
rect 7757 8789 7791 8823
rect 11437 8789 11471 8823
rect 18061 8789 18095 8823
rect 1593 8585 1627 8619
rect 1961 8585 1995 8619
rect 3249 8585 3283 8619
rect 3801 8585 3835 8619
rect 5825 8585 5859 8619
rect 8677 8585 8711 8619
rect 9229 8585 9263 8619
rect 10885 8585 10919 8619
rect 12265 8585 12299 8619
rect 15117 8585 15151 8619
rect 16129 8585 16163 8619
rect 24685 8585 24719 8619
rect 7481 8517 7515 8551
rect 10517 8517 10551 8551
rect 12725 8517 12759 8551
rect 14657 8517 14691 8551
rect 16405 8517 16439 8551
rect 18889 8517 18923 8551
rect 2881 8449 2915 8483
rect 4261 8449 4295 8483
rect 6929 8449 6963 8483
rect 7849 8449 7883 8483
rect 9321 8449 9355 8483
rect 18153 8449 18187 8483
rect 18429 8449 18463 8483
rect 2145 8381 2179 8415
rect 2237 8381 2271 8415
rect 2421 8381 2455 8415
rect 11136 8381 11170 8415
rect 12909 8381 12943 8415
rect 13369 8381 13403 8415
rect 13737 8381 13771 8415
rect 14105 8381 14139 8415
rect 14381 8381 14415 8415
rect 15209 8381 15243 8415
rect 16957 8381 16991 8415
rect 17325 8381 17359 8415
rect 17785 8381 17819 8415
rect 5457 8313 5491 8347
rect 6285 8313 6319 8347
rect 7021 8313 7055 8347
rect 9597 8313 9631 8347
rect 17095 8313 17129 8347
rect 18245 8313 18279 8347
rect 19441 8449 19475 8483
rect 4077 8245 4111 8279
rect 4629 8245 4663 8279
rect 5181 8245 5215 8279
rect 6561 8245 6595 8279
rect 10241 8245 10275 8279
rect 11207 8245 11241 8279
rect 11621 8245 11655 8279
rect 15577 8245 15611 8279
rect 16773 8245 16807 8279
rect 17325 8245 17359 8279
rect 17417 8245 17451 8279
rect 18889 8245 18923 8279
rect 19073 8245 19107 8279
rect 23857 8245 23891 8279
rect 1593 8041 1627 8075
rect 2237 8041 2271 8075
rect 3525 8041 3559 8075
rect 4629 8041 4663 8075
rect 7297 8041 7331 8075
rect 9321 8041 9355 8075
rect 10149 8041 10183 8075
rect 10609 8041 10643 8075
rect 11161 8041 11195 8075
rect 12357 8041 12391 8075
rect 13553 8041 13587 8075
rect 15025 8041 15059 8075
rect 15945 8041 15979 8075
rect 17509 8041 17543 8075
rect 3801 7973 3835 8007
rect 8033 7973 8067 8007
rect 12633 7973 12667 8007
rect 12725 7973 12759 8007
rect 15485 7973 15519 8007
rect 16681 7973 16715 8007
rect 17233 7973 17267 8007
rect 18797 7973 18831 8007
rect 1409 7905 1443 7939
rect 2421 7905 2455 7939
rect 4261 7905 4295 7939
rect 6929 7905 6963 7939
rect 9724 7905 9758 7939
rect 9827 7905 9861 7939
rect 12081 7905 12115 7939
rect 18153 7905 18187 7939
rect 24593 7905 24627 7939
rect 7021 7837 7055 7871
rect 7941 7837 7975 7871
rect 10793 7837 10827 7871
rect 16589 7837 16623 7871
rect 8493 7769 8527 7803
rect 13185 7769 13219 7803
rect 2651 7701 2685 7735
rect 5181 7701 5215 7735
rect 5457 7701 5491 7735
rect 11713 7701 11747 7735
rect 24777 7701 24811 7735
rect 1685 7497 1719 7531
rect 7849 7497 7883 7531
rect 10057 7497 10091 7531
rect 11161 7497 11195 7531
rect 15761 7497 15795 7531
rect 16865 7497 16899 7531
rect 18245 7497 18279 7531
rect 24685 7497 24719 7531
rect 2605 7429 2639 7463
rect 6377 7429 6411 7463
rect 7573 7429 7607 7463
rect 5181 7361 5215 7395
rect 5457 7361 5491 7395
rect 8493 7361 8527 7395
rect 9597 7361 9631 7395
rect 10241 7361 10275 7395
rect 12265 7361 12299 7395
rect 12449 7361 12483 7395
rect 16589 7361 16623 7395
rect 3433 7293 3467 7327
rect 4169 7293 4203 7327
rect 11897 7293 11931 7327
rect 12541 7293 12575 7327
rect 16129 7293 16163 7327
rect 4261 7225 4295 7259
rect 5273 7225 5307 7259
rect 7021 7225 7055 7259
rect 8125 7225 8159 7259
rect 8217 7225 8251 7259
rect 10333 7225 10367 7259
rect 10885 7225 10919 7259
rect 4537 7157 4571 7191
rect 4905 7157 4939 7191
rect 17325 7157 17359 7191
rect 4261 6953 4295 6987
rect 8125 6953 8159 6987
rect 8401 6953 8435 6987
rect 10793 6953 10827 6987
rect 12541 6953 12575 6987
rect 5181 6885 5215 6919
rect 6745 6885 6779 6919
rect 9965 6885 9999 6919
rect 11621 6885 11655 6919
rect 12173 6885 12207 6919
rect 24593 6817 24627 6851
rect 5089 6749 5123 6783
rect 5549 6749 5583 6783
rect 6653 6749 6687 6783
rect 9873 6749 9907 6783
rect 10517 6749 10551 6783
rect 11529 6749 11563 6783
rect 7205 6681 7239 6715
rect 2881 6613 2915 6647
rect 3111 6613 3145 6647
rect 24777 6613 24811 6647
rect 6561 6409 6595 6443
rect 11805 6409 11839 6443
rect 24685 6409 24719 6443
rect 19901 6341 19935 6375
rect 4169 6273 4203 6307
rect 5457 6273 5491 6307
rect 9597 6273 9631 6307
rect 9689 6273 9723 6307
rect 11529 6273 11563 6307
rect 4077 6205 4111 6239
rect 9229 6205 9263 6239
rect 10057 6205 10091 6239
rect 19717 6205 19751 6239
rect 20269 6205 20303 6239
rect 5089 6137 5123 6171
rect 5181 6137 5215 6171
rect 2973 6069 3007 6103
rect 4537 6069 4571 6103
rect 4905 6069 4939 6103
rect 6009 6069 6043 6103
rect 7021 6069 7055 6103
rect 4261 5865 4295 5899
rect 24731 5865 24765 5899
rect 3525 5797 3559 5831
rect 5089 5797 5123 5831
rect 5457 5797 5491 5831
rect 24660 5729 24694 5763
rect 5365 5661 5399 5695
rect 5641 5661 5675 5695
rect 9873 5525 9907 5559
rect 4629 5321 4663 5355
rect 5825 5321 5859 5355
rect 24777 5321 24811 5355
rect 4905 5185 4939 5219
rect 5181 5185 5215 5219
rect 24409 5117 24443 5151
rect 24593 5117 24627 5151
rect 4997 5049 5031 5083
rect 25237 4981 25271 5015
rect 1593 4777 1627 4811
rect 4905 4777 4939 4811
rect 5365 4777 5399 4811
rect 1409 4641 1443 4675
rect 24041 4165 24075 4199
rect 1685 4029 1719 4063
rect 23857 4029 23891 4063
rect 24409 4029 24443 4063
rect 10471 3145 10505 3179
rect 24731 3145 24765 3179
rect 10400 2941 10434 2975
rect 24660 2941 24694 2975
rect 10885 2805 10919 2839
rect 25145 2805 25179 2839
rect 5043 2601 5077 2635
rect 8815 2601 8849 2635
rect 11253 2601 11287 2635
rect 23075 2601 23109 2635
rect 24731 2601 24765 2635
rect 4972 2465 5006 2499
rect 8744 2465 8778 2499
rect 10609 2465 10643 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 15485 2465 15519 2499
rect 16037 2465 16071 2499
rect 23004 2465 23038 2499
rect 23489 2465 23523 2499
rect 24660 2465 24694 2499
rect 10793 2329 10827 2363
rect 15669 2329 15703 2363
rect 5457 2261 5491 2295
rect 9137 2261 9171 2295
rect 12817 2261 12851 2295
rect 25145 2261 25179 2295
<< metal1 >>
rect 3234 27480 3240 27532
rect 3292 27520 3298 27532
rect 3970 27520 3976 27532
rect 3292 27492 3976 27520
rect 3292 27480 3298 27492
rect 3970 27480 3976 27492
rect 4028 27480 4034 27532
rect 11238 27480 11244 27532
rect 11296 27520 11302 27532
rect 12250 27520 12256 27532
rect 11296 27492 12256 27520
rect 11296 27480 11302 27492
rect 12250 27480 12256 27492
rect 12308 27480 12314 27532
rect 26234 27480 26240 27532
rect 26292 27520 26298 27532
rect 27062 27520 27068 27532
rect 26292 27492 27068 27520
rect 26292 27480 26298 27492
rect 27062 27480 27068 27492
rect 27120 27480 27126 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 13541 24395 13599 24401
rect 13541 24361 13553 24395
rect 13587 24392 13599 24395
rect 13906 24392 13912 24404
rect 13587 24364 13912 24392
rect 13587 24361 13599 24364
rect 13541 24355 13599 24361
rect 13906 24352 13912 24364
rect 13964 24352 13970 24404
rect 5420 24259 5478 24265
rect 5420 24225 5432 24259
rect 5466 24256 5478 24259
rect 5534 24256 5540 24268
rect 5466 24228 5540 24256
rect 5466 24225 5478 24228
rect 5420 24219 5478 24225
rect 5534 24216 5540 24228
rect 5592 24216 5598 24268
rect 13354 24256 13360 24268
rect 13315 24228 13360 24256
rect 13354 24216 13360 24228
rect 13412 24216 13418 24268
rect 4614 24012 4620 24064
rect 4672 24052 4678 24064
rect 5491 24055 5549 24061
rect 5491 24052 5503 24055
rect 4672 24024 5503 24052
rect 4672 24012 4678 24024
rect 5491 24021 5503 24024
rect 5537 24021 5549 24055
rect 5491 24015 5549 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 5813 23851 5871 23857
rect 5813 23848 5825 23851
rect 5592 23820 5825 23848
rect 5592 23808 5598 23820
rect 5813 23817 5825 23820
rect 5859 23817 5871 23851
rect 13354 23848 13360 23860
rect 13315 23820 13360 23848
rect 5813 23811 5871 23817
rect 13354 23808 13360 23820
rect 13412 23808 13418 23860
rect 13633 23851 13691 23857
rect 13633 23817 13645 23851
rect 13679 23848 13691 23851
rect 15470 23848 15476 23860
rect 13679 23820 15476 23848
rect 13679 23817 13691 23820
rect 13633 23811 13691 23817
rect 15470 23808 15476 23820
rect 15528 23808 15534 23860
rect 18233 23851 18291 23857
rect 18233 23817 18245 23851
rect 18279 23848 18291 23851
rect 20438 23848 20444 23860
rect 18279 23820 20444 23848
rect 18279 23817 18291 23820
rect 18233 23811 18291 23817
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 21453 23851 21511 23857
rect 21453 23817 21465 23851
rect 21499 23848 21511 23851
rect 22094 23848 22100 23860
rect 21499 23820 22100 23848
rect 21499 23817 21511 23820
rect 21453 23811 21511 23817
rect 22094 23808 22100 23820
rect 22152 23808 22158 23860
rect 5258 23604 5264 23656
rect 5316 23644 5322 23656
rect 5388 23647 5446 23653
rect 5388 23644 5400 23647
rect 5316 23616 5400 23644
rect 5316 23604 5322 23616
rect 5388 23613 5400 23616
rect 5434 23644 5446 23647
rect 6181 23647 6239 23653
rect 6181 23644 6193 23647
rect 5434 23616 6193 23644
rect 5434 23613 5446 23616
rect 5388 23607 5446 23613
rect 6181 23613 6193 23616
rect 6227 23613 6239 23647
rect 6181 23607 6239 23613
rect 13449 23647 13507 23653
rect 13449 23613 13461 23647
rect 13495 23644 13507 23647
rect 18046 23644 18052 23656
rect 13495 23616 13814 23644
rect 17959 23616 18052 23644
rect 13495 23613 13507 23616
rect 13449 23607 13507 23613
rect 5491 23511 5549 23517
rect 5491 23477 5503 23511
rect 5537 23508 5549 23511
rect 5718 23508 5724 23520
rect 5537 23480 5724 23508
rect 5537 23477 5549 23480
rect 5491 23471 5549 23477
rect 5718 23468 5724 23480
rect 5776 23468 5782 23520
rect 13786 23508 13814 23616
rect 18046 23604 18052 23616
rect 18104 23644 18110 23656
rect 18601 23647 18659 23653
rect 18601 23644 18613 23647
rect 18104 23616 18613 23644
rect 18104 23604 18110 23616
rect 18601 23613 18613 23616
rect 18647 23613 18659 23647
rect 21266 23644 21272 23656
rect 21179 23616 21272 23644
rect 18601 23607 18659 23613
rect 21266 23604 21272 23616
rect 21324 23644 21330 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21324 23616 21833 23644
rect 21324 23604 21330 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 14093 23511 14151 23517
rect 14093 23508 14105 23511
rect 13786 23480 14105 23508
rect 14093 23477 14105 23480
rect 14139 23508 14151 23511
rect 14642 23508 14648 23520
rect 14139 23480 14648 23508
rect 14139 23477 14151 23480
rect 14093 23471 14151 23477
rect 14642 23468 14648 23480
rect 14700 23468 14706 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 5718 23264 5724 23316
rect 5776 23304 5782 23316
rect 6825 23307 6883 23313
rect 6825 23304 6837 23307
rect 5776 23276 6837 23304
rect 5776 23264 5782 23276
rect 6825 23273 6837 23276
rect 6871 23304 6883 23307
rect 6914 23304 6920 23316
rect 6871 23276 6920 23304
rect 6871 23273 6883 23276
rect 6825 23267 6883 23273
rect 6914 23264 6920 23276
rect 6972 23264 6978 23316
rect 13354 23264 13360 23316
rect 13412 23304 13418 23316
rect 13955 23307 14013 23313
rect 13955 23304 13967 23307
rect 13412 23276 13967 23304
rect 13412 23264 13418 23276
rect 13955 23273 13967 23276
rect 14001 23273 14013 23307
rect 13955 23267 14013 23273
rect 16347 23307 16405 23313
rect 16347 23273 16359 23307
rect 16393 23304 16405 23307
rect 18046 23304 18052 23316
rect 16393 23276 18052 23304
rect 16393 23273 16405 23276
rect 16347 23267 16405 23273
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 13884 23171 13942 23177
rect 13884 23137 13896 23171
rect 13930 23168 13942 23171
rect 14550 23168 14556 23180
rect 13930 23140 14556 23168
rect 13930 23137 13942 23140
rect 13884 23131 13942 23137
rect 14550 23128 14556 23140
rect 14608 23128 14614 23180
rect 16114 23168 16120 23180
rect 16075 23140 16120 23168
rect 16114 23128 16120 23140
rect 16172 23128 16178 23180
rect 24648 23171 24706 23177
rect 24648 23137 24660 23171
rect 24694 23168 24706 23171
rect 25130 23168 25136 23180
rect 24694 23140 25136 23168
rect 24694 23137 24706 23140
rect 24648 23131 24706 23137
rect 25130 23128 25136 23140
rect 25188 23128 25194 23180
rect 13170 22924 13176 22976
rect 13228 22964 13234 22976
rect 13633 22967 13691 22973
rect 13633 22964 13645 22967
rect 13228 22936 13645 22964
rect 13228 22924 13234 22936
rect 13633 22933 13645 22936
rect 13679 22964 13691 22967
rect 13814 22964 13820 22976
rect 13679 22936 13820 22964
rect 13679 22933 13691 22936
rect 13633 22927 13691 22933
rect 13814 22924 13820 22936
rect 13872 22924 13878 22976
rect 21450 22924 21456 22976
rect 21508 22964 21514 22976
rect 24719 22967 24777 22973
rect 24719 22964 24731 22967
rect 21508 22936 24731 22964
rect 21508 22924 21514 22936
rect 24719 22933 24731 22936
rect 24765 22933 24777 22967
rect 24719 22927 24777 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1854 22760 1860 22772
rect 1815 22732 1860 22760
rect 1854 22720 1860 22732
rect 1912 22720 1918 22772
rect 14550 22760 14556 22772
rect 14511 22732 14556 22760
rect 14550 22720 14556 22732
rect 14608 22760 14614 22772
rect 15378 22760 15384 22772
rect 14608 22732 15384 22760
rect 14608 22720 14614 22732
rect 15378 22720 15384 22732
rect 15436 22720 15442 22772
rect 20119 22763 20177 22769
rect 20119 22729 20131 22763
rect 20165 22760 20177 22763
rect 21266 22760 21272 22772
rect 20165 22732 21272 22760
rect 20165 22729 20177 22732
rect 20119 22723 20177 22729
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 25498 22760 25504 22772
rect 25459 22732 25504 22760
rect 25498 22720 25504 22732
rect 25556 22720 25562 22772
rect 6641 22695 6699 22701
rect 6641 22661 6653 22695
rect 6687 22692 6699 22695
rect 7006 22692 7012 22704
rect 6687 22664 7012 22692
rect 6687 22661 6699 22664
rect 6641 22655 6699 22661
rect 7006 22652 7012 22664
rect 7064 22652 7070 22704
rect 25130 22692 25136 22704
rect 25043 22664 25136 22692
rect 25130 22652 25136 22664
rect 25188 22692 25194 22704
rect 27614 22692 27620 22704
rect 25188 22664 27620 22692
rect 25188 22652 25194 22664
rect 27614 22652 27620 22664
rect 27672 22652 27678 22704
rect 6914 22624 6920 22636
rect 6875 22596 6920 22624
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 1448 22559 1506 22565
rect 1448 22525 1460 22559
rect 1494 22556 1506 22559
rect 1854 22556 1860 22568
rect 1494 22528 1860 22556
rect 1494 22525 1506 22528
rect 1448 22519 1506 22525
rect 1854 22516 1860 22528
rect 1912 22516 1918 22568
rect 8732 22559 8790 22565
rect 8732 22525 8744 22559
rect 8778 22556 8790 22559
rect 13541 22559 13599 22565
rect 13541 22556 13553 22559
rect 8778 22528 9260 22556
rect 8778 22525 8790 22528
rect 8732 22519 8790 22525
rect 1535 22491 1593 22497
rect 1535 22457 1547 22491
rect 1581 22488 1593 22491
rect 1581 22460 6960 22488
rect 1581 22457 1593 22460
rect 1535 22451 1593 22457
rect 6932 22420 6960 22460
rect 7006 22448 7012 22500
rect 7064 22488 7070 22500
rect 7558 22488 7564 22500
rect 7064 22460 7109 22488
rect 7471 22460 7564 22488
rect 7064 22448 7070 22460
rect 7558 22448 7564 22460
rect 7616 22488 7622 22500
rect 8570 22488 8576 22500
rect 7616 22460 8576 22488
rect 7616 22448 7622 22460
rect 8570 22448 8576 22460
rect 8628 22448 8634 22500
rect 8662 22420 8668 22432
rect 6932 22392 8668 22420
rect 8662 22380 8668 22392
rect 8720 22380 8726 22432
rect 8803 22423 8861 22429
rect 8803 22389 8815 22423
rect 8849 22420 8861 22423
rect 8938 22420 8944 22432
rect 8849 22392 8944 22420
rect 8849 22389 8861 22392
rect 8803 22383 8861 22389
rect 8938 22380 8944 22392
rect 8996 22380 9002 22432
rect 9232 22429 9260 22528
rect 13372 22528 13553 22556
rect 9217 22423 9275 22429
rect 9217 22389 9229 22423
rect 9263 22420 9275 22423
rect 9766 22420 9772 22432
rect 9263 22392 9772 22420
rect 9263 22389 9275 22392
rect 9217 22383 9275 22389
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 13372 22429 13400 22528
rect 13541 22525 13553 22528
rect 13587 22525 13599 22559
rect 13541 22519 13599 22525
rect 13814 22516 13820 22568
rect 13872 22556 13878 22568
rect 14001 22559 14059 22565
rect 14001 22556 14013 22559
rect 13872 22528 14013 22556
rect 13872 22516 13878 22528
rect 14001 22525 14013 22528
rect 14047 22525 14059 22559
rect 14001 22519 14059 22525
rect 20048 22559 20106 22565
rect 20048 22525 20060 22559
rect 20094 22556 20106 22559
rect 24648 22559 24706 22565
rect 20094 22528 20392 22556
rect 20094 22525 20106 22528
rect 20048 22519 20106 22525
rect 14274 22488 14280 22500
rect 14235 22460 14280 22488
rect 14274 22448 14280 22460
rect 14332 22448 14338 22500
rect 20364 22432 20392 22528
rect 24648 22525 24660 22559
rect 24694 22556 24706 22559
rect 25498 22556 25504 22568
rect 24694 22528 25504 22556
rect 24694 22525 24706 22528
rect 24648 22519 24706 22525
rect 25498 22516 25504 22528
rect 25556 22516 25562 22568
rect 13357 22423 13415 22429
rect 13357 22420 13369 22423
rect 11112 22392 13369 22420
rect 11112 22380 11118 22392
rect 13357 22389 13369 22392
rect 13403 22389 13415 22423
rect 13357 22383 13415 22389
rect 14826 22380 14832 22432
rect 14884 22420 14890 22432
rect 16114 22420 16120 22432
rect 14884 22392 16120 22420
rect 14884 22380 14890 22392
rect 16114 22380 16120 22392
rect 16172 22420 16178 22432
rect 16209 22423 16267 22429
rect 16209 22420 16221 22423
rect 16172 22392 16221 22420
rect 16172 22380 16178 22392
rect 16209 22389 16221 22392
rect 16255 22389 16267 22423
rect 16209 22383 16267 22389
rect 20346 22380 20352 22432
rect 20404 22420 20410 22432
rect 20441 22423 20499 22429
rect 20441 22420 20453 22423
rect 20404 22392 20453 22420
rect 20404 22380 20410 22392
rect 20441 22389 20453 22392
rect 20487 22389 20499 22423
rect 20441 22383 20499 22389
rect 21634 22380 21640 22432
rect 21692 22420 21698 22432
rect 24719 22423 24777 22429
rect 24719 22420 24731 22423
rect 21692 22392 24731 22420
rect 21692 22380 21698 22392
rect 24719 22389 24731 22392
rect 24765 22389 24777 22423
rect 24719 22383 24777 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 8938 22216 8944 22228
rect 8899 22188 8944 22216
rect 8938 22176 8944 22188
rect 8996 22176 9002 22228
rect 18782 22216 18788 22228
rect 12636 22188 18788 22216
rect 6454 22148 6460 22160
rect 6415 22120 6460 22148
rect 6454 22108 6460 22120
rect 6512 22108 6518 22160
rect 7009 22151 7067 22157
rect 7009 22117 7021 22151
rect 7055 22148 7067 22151
rect 7558 22148 7564 22160
rect 7055 22120 7564 22148
rect 7055 22117 7067 22120
rect 7009 22111 7067 22117
rect 7558 22108 7564 22120
rect 7616 22108 7622 22160
rect 8018 22148 8024 22160
rect 7979 22120 8024 22148
rect 8018 22108 8024 22120
rect 8076 22108 8082 22160
rect 8662 22108 8668 22160
rect 8720 22148 8726 22160
rect 12437 22151 12495 22157
rect 12437 22148 12449 22151
rect 8720 22120 12449 22148
rect 8720 22108 8726 22120
rect 12437 22117 12449 22120
rect 12483 22148 12495 22151
rect 12526 22148 12532 22160
rect 12483 22120 12532 22148
rect 12483 22117 12495 22120
rect 12437 22111 12495 22117
rect 12526 22108 12532 22120
rect 12584 22108 12590 22160
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 1486 22080 1492 22092
rect 1443 22052 1492 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 1486 22040 1492 22052
rect 1544 22040 1550 22092
rect 9766 22089 9772 22092
rect 9744 22083 9772 22089
rect 9744 22080 9756 22083
rect 9679 22052 9756 22080
rect 9744 22049 9756 22052
rect 9824 22080 9830 22092
rect 12636 22080 12664 22188
rect 18782 22176 18788 22188
rect 18840 22176 18846 22228
rect 21450 22216 21456 22228
rect 21411 22188 21456 22216
rect 21450 22176 21456 22188
rect 21508 22176 21514 22228
rect 12986 22148 12992 22160
rect 12947 22120 12992 22148
rect 12986 22108 12992 22120
rect 13044 22108 13050 22160
rect 16853 22151 16911 22157
rect 16853 22117 16865 22151
rect 16899 22148 16911 22151
rect 17402 22148 17408 22160
rect 16899 22120 17408 22148
rect 16899 22117 16911 22120
rect 16853 22111 16911 22117
rect 17402 22108 17408 22120
rect 17460 22108 17466 22160
rect 23934 22148 23940 22160
rect 23559 22120 23940 22148
rect 9824 22052 12664 22080
rect 18300 22083 18358 22089
rect 9744 22043 9772 22049
rect 9766 22040 9772 22043
rect 9824 22040 9830 22052
rect 18300 22049 18312 22083
rect 18346 22080 18358 22083
rect 19150 22080 19156 22092
rect 18346 22052 19156 22080
rect 18346 22049 18358 22052
rect 18300 22043 18358 22049
rect 19150 22040 19156 22052
rect 19208 22040 19214 22092
rect 21980 22083 22038 22089
rect 21980 22049 21992 22083
rect 22026 22080 22038 22083
rect 22370 22080 22376 22092
rect 22026 22052 22376 22080
rect 22026 22049 22038 22052
rect 21980 22043 22038 22049
rect 22370 22040 22376 22052
rect 22428 22040 22434 22092
rect 23559 22089 23587 22120
rect 23934 22108 23940 22120
rect 23992 22148 23998 22160
rect 25406 22148 25412 22160
rect 23992 22120 25412 22148
rect 23992 22108 23998 22120
rect 25406 22108 25412 22120
rect 25464 22108 25470 22160
rect 24670 22089 24676 22092
rect 23544 22083 23602 22089
rect 23544 22049 23556 22083
rect 23590 22049 23602 22083
rect 24648 22083 24676 22089
rect 24648 22080 24660 22083
rect 24583 22052 24660 22080
rect 23544 22043 23602 22049
rect 24648 22049 24660 22052
rect 24728 22080 24734 22092
rect 25222 22080 25228 22092
rect 24728 22052 25228 22080
rect 24648 22043 24676 22049
rect 24670 22040 24676 22043
rect 24728 22040 24734 22052
rect 25222 22040 25228 22052
rect 25280 22040 25286 22092
rect 5534 21972 5540 22024
rect 5592 22012 5598 22024
rect 6365 22015 6423 22021
rect 6365 22012 6377 22015
rect 5592 21984 6377 22012
rect 5592 21972 5598 21984
rect 6365 21981 6377 21984
rect 6411 21981 6423 22015
rect 7926 22012 7932 22024
rect 7887 21984 7932 22012
rect 6365 21975 6423 21981
rect 7926 21972 7932 21984
rect 7984 21972 7990 22024
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 8662 22012 8668 22024
rect 8619 21984 8668 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 8662 21972 8668 21984
rect 8720 21972 8726 22024
rect 12894 22012 12900 22024
rect 12855 21984 12900 22012
rect 12894 21972 12900 21984
rect 12952 21972 12958 22024
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 13814 22012 13820 22024
rect 13587 21984 13820 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 15562 22012 15568 22024
rect 15523 21984 15568 22012
rect 15562 21972 15568 21984
rect 15620 21972 15626 22024
rect 16761 22015 16819 22021
rect 16761 21981 16773 22015
rect 16807 21981 16819 22015
rect 17034 22012 17040 22024
rect 16995 21984 17040 22012
rect 16761 21975 16819 21981
rect 10962 21904 10968 21956
rect 11020 21944 11026 21956
rect 15838 21944 15844 21956
rect 11020 21916 15844 21944
rect 11020 21904 11026 21916
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 15930 21904 15936 21956
rect 15988 21944 15994 21956
rect 16776 21944 16804 21975
rect 17034 21972 17040 21984
rect 17092 21972 17098 22024
rect 20898 22012 20904 22024
rect 20859 21984 20904 22012
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 23615 21947 23673 21953
rect 23615 21944 23627 21947
rect 15988 21916 23627 21944
rect 15988 21904 15994 21916
rect 23615 21913 23627 21916
rect 23661 21913 23673 21947
rect 23615 21907 23673 21913
rect 1535 21879 1593 21885
rect 1535 21845 1547 21879
rect 1581 21876 1593 21879
rect 5534 21876 5540 21888
rect 1581 21848 5540 21876
rect 1581 21845 1593 21848
rect 1535 21839 1593 21845
rect 5534 21836 5540 21848
rect 5592 21836 5598 21888
rect 9815 21879 9873 21885
rect 9815 21845 9827 21879
rect 9861 21876 9873 21879
rect 9950 21876 9956 21888
rect 9861 21848 9956 21876
rect 9861 21845 9873 21848
rect 9815 21839 9873 21845
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 14182 21836 14188 21888
rect 14240 21876 14246 21888
rect 14461 21879 14519 21885
rect 14461 21876 14473 21879
rect 14240 21848 14473 21876
rect 14240 21836 14246 21848
rect 14461 21845 14473 21848
rect 14507 21845 14519 21879
rect 14461 21839 14519 21845
rect 16482 21836 16488 21888
rect 16540 21876 16546 21888
rect 18371 21879 18429 21885
rect 18371 21876 18383 21879
rect 16540 21848 18383 21876
rect 16540 21836 16546 21848
rect 18371 21845 18383 21848
rect 18417 21845 18429 21879
rect 18371 21839 18429 21845
rect 22051 21879 22109 21885
rect 22051 21845 22063 21879
rect 22097 21876 22109 21879
rect 22186 21876 22192 21888
rect 22097 21848 22192 21876
rect 22097 21845 22109 21848
rect 22051 21839 22109 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 24026 21836 24032 21888
rect 24084 21876 24090 21888
rect 24719 21879 24777 21885
rect 24719 21876 24731 21879
rect 24084 21848 24731 21876
rect 24084 21836 24090 21848
rect 24719 21845 24731 21848
rect 24765 21845 24777 21879
rect 24719 21839 24777 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1486 21632 1492 21684
rect 1544 21672 1550 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1544 21644 1593 21672
rect 1544 21632 1550 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 5534 21672 5540 21684
rect 5495 21644 5540 21672
rect 1581 21635 1639 21641
rect 5534 21632 5540 21644
rect 5592 21632 5598 21684
rect 7006 21632 7012 21684
rect 7064 21672 7070 21684
rect 7742 21672 7748 21684
rect 7064 21644 7748 21672
rect 7064 21632 7070 21644
rect 7742 21632 7748 21644
rect 7800 21672 7806 21684
rect 8297 21675 8355 21681
rect 8297 21672 8309 21675
rect 7800 21644 8309 21672
rect 7800 21632 7806 21644
rect 8297 21641 8309 21644
rect 8343 21641 8355 21675
rect 8297 21635 8355 21641
rect 8018 21604 8024 21616
rect 7979 21576 8024 21604
rect 8018 21564 8024 21576
rect 8076 21564 8082 21616
rect 4154 21360 4160 21412
rect 4212 21400 4218 21412
rect 6549 21403 6607 21409
rect 6549 21400 6561 21403
rect 4212 21372 6561 21400
rect 4212 21360 4218 21372
rect 6549 21369 6561 21372
rect 6595 21400 6607 21403
rect 7009 21403 7067 21409
rect 7009 21400 7021 21403
rect 6595 21372 7021 21400
rect 6595 21369 6607 21372
rect 6549 21363 6607 21369
rect 7009 21369 7021 21372
rect 7055 21369 7067 21403
rect 7009 21363 7067 21369
rect 7098 21360 7104 21412
rect 7156 21400 7162 21412
rect 7653 21403 7711 21409
rect 7156 21372 7201 21400
rect 7156 21360 7162 21372
rect 7653 21369 7665 21403
rect 7699 21400 7711 21403
rect 7834 21400 7840 21412
rect 7699 21372 7840 21400
rect 7699 21369 7711 21372
rect 7653 21363 7711 21369
rect 7834 21360 7840 21372
rect 7892 21360 7898 21412
rect 8312 21400 8340 21635
rect 9030 21632 9036 21684
rect 9088 21672 9094 21684
rect 10229 21675 10287 21681
rect 10229 21672 10241 21675
rect 9088 21644 10241 21672
rect 9088 21632 9094 21644
rect 10229 21641 10241 21644
rect 10275 21641 10287 21675
rect 10229 21635 10287 21641
rect 12894 21632 12900 21684
rect 12952 21672 12958 21684
rect 15930 21672 15936 21684
rect 12952 21644 13814 21672
rect 15891 21644 15936 21672
rect 12952 21632 12958 21644
rect 9766 21604 9772 21616
rect 9727 21576 9772 21604
rect 9766 21564 9772 21576
rect 9824 21564 9830 21616
rect 13786 21604 13814 21644
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 22370 21672 22376 21684
rect 22331 21644 22376 21672
rect 22370 21632 22376 21644
rect 22428 21672 22434 21684
rect 23750 21672 23756 21684
rect 22428 21644 23756 21672
rect 22428 21632 22434 21644
rect 23750 21632 23756 21644
rect 23808 21632 23814 21684
rect 23934 21672 23940 21684
rect 23895 21644 23940 21672
rect 23934 21632 23940 21644
rect 23992 21632 23998 21684
rect 24670 21672 24676 21684
rect 24631 21644 24676 21672
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 17034 21604 17040 21616
rect 13786 21576 17040 21604
rect 8573 21539 8631 21545
rect 8573 21505 8585 21539
rect 8619 21536 8631 21539
rect 8938 21536 8944 21548
rect 8619 21508 8944 21536
rect 8619 21505 8631 21508
rect 8573 21499 8631 21505
rect 8938 21496 8944 21508
rect 8996 21496 9002 21548
rect 12526 21536 12532 21548
rect 12487 21508 12532 21536
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 12894 21536 12900 21548
rect 12855 21508 12900 21536
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 13630 21496 13636 21548
rect 13688 21536 13694 21548
rect 16482 21536 16488 21548
rect 13688 21508 13814 21536
rect 16443 21508 16488 21536
rect 13688 21496 13694 21508
rect 10042 21468 10048 21480
rect 10003 21440 10048 21468
rect 10042 21428 10048 21440
rect 10100 21468 10106 21480
rect 10597 21471 10655 21477
rect 10597 21468 10609 21471
rect 10100 21440 10609 21468
rect 10100 21428 10106 21440
rect 10597 21437 10609 21440
rect 10643 21437 10655 21471
rect 13786 21468 13814 21508
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 16776 21545 16804 21576
rect 17034 21564 17040 21576
rect 17092 21564 17098 21616
rect 16761 21539 16819 21545
rect 16761 21505 16773 21539
rect 16807 21505 16819 21539
rect 16761 21499 16819 21505
rect 17126 21496 17132 21548
rect 17184 21536 17190 21548
rect 19150 21536 19156 21548
rect 17184 21508 19057 21536
rect 19111 21508 19156 21536
rect 17184 21496 17190 21508
rect 14369 21471 14427 21477
rect 14369 21468 14381 21471
rect 13786 21440 14381 21468
rect 10597 21431 10655 21437
rect 14369 21437 14381 21440
rect 14415 21468 14427 21471
rect 14461 21471 14519 21477
rect 14461 21468 14473 21471
rect 14415 21440 14473 21468
rect 14415 21437 14427 21440
rect 14369 21431 14427 21437
rect 14461 21437 14473 21440
rect 14507 21437 14519 21471
rect 14461 21431 14519 21437
rect 14921 21471 14979 21477
rect 14921 21437 14933 21471
rect 14967 21437 14979 21471
rect 14921 21431 14979 21437
rect 17865 21471 17923 21477
rect 17865 21437 17877 21471
rect 17911 21468 17923 21471
rect 18049 21471 18107 21477
rect 18049 21468 18061 21471
rect 17911 21440 18061 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 18049 21437 18061 21440
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 8665 21403 8723 21409
rect 8665 21400 8677 21403
rect 8312 21372 8677 21400
rect 8665 21369 8677 21372
rect 8711 21369 8723 21403
rect 9214 21400 9220 21412
rect 9175 21372 9220 21400
rect 8665 21363 8723 21369
rect 9214 21360 9220 21372
rect 9272 21360 9278 21412
rect 12621 21403 12679 21409
rect 12621 21369 12633 21403
rect 12667 21369 12679 21403
rect 12621 21363 12679 21369
rect 5905 21335 5963 21341
rect 5905 21301 5917 21335
rect 5951 21332 5963 21335
rect 6273 21335 6331 21341
rect 6273 21332 6285 21335
rect 5951 21304 6285 21332
rect 5951 21301 5963 21304
rect 5905 21295 5963 21301
rect 6273 21301 6285 21304
rect 6319 21332 6331 21335
rect 6454 21332 6460 21344
rect 6319 21304 6460 21332
rect 6319 21301 6331 21304
rect 6273 21295 6331 21301
rect 6454 21292 6460 21304
rect 6512 21332 6518 21344
rect 7116 21332 7144 21360
rect 12250 21332 12256 21344
rect 6512 21304 7144 21332
rect 12211 21304 12256 21332
rect 6512 21292 6518 21304
rect 12250 21292 12256 21304
rect 12308 21332 12314 21344
rect 12636 21332 12664 21363
rect 14182 21360 14188 21412
rect 14240 21400 14246 21412
rect 14936 21400 14964 21431
rect 14240 21372 14964 21400
rect 15197 21403 15255 21409
rect 14240 21360 14246 21372
rect 15197 21369 15209 21403
rect 15243 21400 15255 21403
rect 15286 21400 15292 21412
rect 15243 21372 15292 21400
rect 15243 21369 15255 21372
rect 15197 21363 15255 21369
rect 15286 21360 15292 21372
rect 15344 21360 15350 21412
rect 16577 21403 16635 21409
rect 16577 21369 16589 21403
rect 16623 21369 16635 21403
rect 16577 21363 16635 21369
rect 12308 21304 12664 21332
rect 12308 21292 12314 21304
rect 12802 21292 12808 21344
rect 12860 21332 12866 21344
rect 12986 21332 12992 21344
rect 12860 21304 12992 21332
rect 12860 21292 12866 21304
rect 12986 21292 12992 21304
rect 13044 21332 13050 21344
rect 13449 21335 13507 21341
rect 13449 21332 13461 21335
rect 13044 21304 13461 21332
rect 13044 21292 13050 21304
rect 13449 21301 13461 21304
rect 13495 21301 13507 21335
rect 13449 21295 13507 21301
rect 15930 21292 15936 21344
rect 15988 21332 15994 21344
rect 16209 21335 16267 21341
rect 16209 21332 16221 21335
rect 15988 21304 16221 21332
rect 15988 21292 15994 21304
rect 16209 21301 16221 21304
rect 16255 21332 16267 21335
rect 16592 21332 16620 21363
rect 16850 21360 16856 21412
rect 16908 21400 16914 21412
rect 17880 21400 17908 21431
rect 18138 21428 18144 21480
rect 18196 21468 18202 21480
rect 18509 21471 18567 21477
rect 18509 21468 18521 21471
rect 18196 21440 18521 21468
rect 18196 21428 18202 21440
rect 18509 21437 18521 21440
rect 18555 21437 18567 21471
rect 19029 21468 19057 21508
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 21450 21536 21456 21548
rect 21411 21508 21456 21536
rect 21450 21496 21456 21508
rect 21508 21496 21514 21548
rect 21542 21496 21548 21548
rect 21600 21536 21606 21548
rect 21729 21539 21787 21545
rect 21729 21536 21741 21539
rect 21600 21508 21741 21536
rect 21600 21496 21606 21508
rect 21729 21505 21741 21508
rect 21775 21505 21787 21539
rect 21729 21499 21787 21505
rect 19648 21471 19706 21477
rect 19648 21468 19660 21471
rect 19029 21440 19660 21468
rect 18509 21431 18567 21437
rect 19648 21437 19660 21440
rect 19694 21468 19706 21471
rect 20073 21471 20131 21477
rect 20073 21468 20085 21471
rect 19694 21440 20085 21468
rect 19694 21437 19706 21440
rect 19648 21431 19706 21437
rect 20073 21437 20085 21440
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 18782 21400 18788 21412
rect 16908 21372 17908 21400
rect 18743 21372 18788 21400
rect 16908 21360 16914 21372
rect 18782 21360 18788 21372
rect 18840 21360 18846 21412
rect 21545 21403 21603 21409
rect 21545 21369 21557 21403
rect 21591 21369 21603 21403
rect 21545 21363 21603 21369
rect 17402 21332 17408 21344
rect 16255 21304 16620 21332
rect 17363 21304 17408 21332
rect 16255 21301 16267 21304
rect 16209 21295 16267 21301
rect 17402 21292 17408 21304
rect 17460 21292 17466 21344
rect 19751 21335 19809 21341
rect 19751 21301 19763 21335
rect 19797 21332 19809 21335
rect 19978 21332 19984 21344
rect 19797 21304 19984 21332
rect 19797 21301 19809 21304
rect 19751 21295 19809 21301
rect 19978 21292 19984 21304
rect 20036 21292 20042 21344
rect 20622 21292 20628 21344
rect 20680 21332 20686 21344
rect 21269 21335 21327 21341
rect 21269 21332 21281 21335
rect 20680 21304 21281 21332
rect 20680 21292 20686 21304
rect 21269 21301 21281 21304
rect 21315 21332 21327 21335
rect 21560 21332 21588 21363
rect 22830 21332 22836 21344
rect 21315 21304 22836 21332
rect 21315 21301 21327 21304
rect 21269 21295 21327 21301
rect 22830 21292 22836 21304
rect 22888 21292 22894 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 7006 21128 7012 21140
rect 6380 21100 7012 21128
rect 6380 21072 6408 21100
rect 7006 21088 7012 21100
rect 7064 21088 7070 21140
rect 8711 21131 8769 21137
rect 8711 21097 8723 21131
rect 8757 21128 8769 21131
rect 10042 21128 10048 21140
rect 8757 21100 10048 21128
rect 8757 21097 8769 21100
rect 8711 21091 8769 21097
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 15427 21131 15485 21137
rect 15427 21128 15439 21131
rect 12176 21100 15439 21128
rect 6362 21060 6368 21072
rect 5403 21032 6368 21060
rect 5403 21001 5431 21032
rect 6362 21020 6368 21032
rect 6420 21020 6426 21072
rect 6638 21060 6644 21072
rect 6599 21032 6644 21060
rect 6638 21020 6644 21032
rect 6696 21020 6702 21072
rect 12176 21069 12204 21100
rect 15427 21097 15439 21100
rect 15473 21097 15485 21131
rect 16482 21128 16488 21140
rect 16443 21100 16488 21128
rect 15427 21091 15485 21097
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 18782 21088 18788 21140
rect 18840 21128 18846 21140
rect 19061 21131 19119 21137
rect 19061 21128 19073 21131
rect 18840 21100 19073 21128
rect 18840 21088 18846 21100
rect 19061 21097 19073 21100
rect 19107 21097 19119 21131
rect 22186 21128 22192 21140
rect 22147 21100 22192 21128
rect 19061 21091 19119 21097
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 11977 21063 12035 21069
rect 11977 21029 11989 21063
rect 12023 21060 12035 21063
rect 12161 21063 12219 21069
rect 12161 21060 12173 21063
rect 12023 21032 12173 21060
rect 12023 21029 12035 21032
rect 11977 21023 12035 21029
rect 12161 21029 12173 21032
rect 12207 21029 12219 21063
rect 12161 21023 12219 21029
rect 12250 21020 12256 21072
rect 12308 21060 12314 21072
rect 12308 21032 12848 21060
rect 12308 21020 12314 21032
rect 5388 20995 5446 21001
rect 5388 20961 5400 20995
rect 5434 20961 5446 20995
rect 5388 20955 5446 20961
rect 5491 20995 5549 21001
rect 5491 20961 5503 20995
rect 5537 20992 5549 20995
rect 7374 20992 7380 21004
rect 5537 20964 7380 20992
rect 5537 20961 5549 20964
rect 5491 20955 5549 20961
rect 7374 20952 7380 20964
rect 7432 20952 7438 21004
rect 8478 20952 8484 21004
rect 8536 20992 8542 21004
rect 8608 20995 8666 21001
rect 8608 20992 8620 20995
rect 8536 20964 8620 20992
rect 8536 20952 8542 20964
rect 8608 20961 8620 20964
rect 8654 20961 8666 20995
rect 10686 20992 10692 21004
rect 10647 20964 10692 20992
rect 8608 20955 8666 20961
rect 10686 20952 10692 20964
rect 10744 20952 10750 21004
rect 11054 20992 11060 21004
rect 11015 20964 11060 20992
rect 11054 20952 11060 20964
rect 11112 20952 11118 21004
rect 12820 20992 12848 21032
rect 12894 21020 12900 21072
rect 12952 21060 12958 21072
rect 13081 21063 13139 21069
rect 13081 21060 13093 21063
rect 12952 21032 13093 21060
rect 12952 21020 12958 21032
rect 13081 21029 13093 21032
rect 13127 21029 13139 21063
rect 13354 21060 13360 21072
rect 13081 21023 13139 21029
rect 13188 21032 13360 21060
rect 13188 20992 13216 21032
rect 13354 21020 13360 21032
rect 13412 21060 13418 21072
rect 13817 21063 13875 21069
rect 13817 21060 13829 21063
rect 13412 21032 13829 21060
rect 13412 21020 13418 21032
rect 13817 21029 13829 21032
rect 13863 21029 13875 21063
rect 16758 21060 16764 21072
rect 16671 21032 16764 21060
rect 13817 21023 13875 21029
rect 16758 21020 16764 21032
rect 16816 21060 16822 21072
rect 17402 21060 17408 21072
rect 16816 21032 17408 21060
rect 16816 21020 16822 21032
rect 17402 21020 17408 21032
rect 17460 21020 17466 21072
rect 19429 21063 19487 21069
rect 19429 21029 19441 21063
rect 19475 21060 19487 21063
rect 19518 21060 19524 21072
rect 19475 21032 19524 21060
rect 19475 21029 19487 21032
rect 19429 21023 19487 21029
rect 19518 21020 19524 21032
rect 19576 21020 19582 21072
rect 20898 21020 20904 21072
rect 20956 21060 20962 21072
rect 21177 21063 21235 21069
rect 21177 21060 21189 21063
rect 20956 21032 21189 21060
rect 20956 21020 20962 21032
rect 21177 21029 21189 21032
rect 21223 21029 21235 21063
rect 21177 21023 21235 21029
rect 21269 21063 21327 21069
rect 21269 21029 21281 21063
rect 21315 21060 21327 21063
rect 21358 21060 21364 21072
rect 21315 21032 21364 21060
rect 21315 21029 21327 21032
rect 21269 21023 21327 21029
rect 21358 21020 21364 21032
rect 21416 21020 21422 21072
rect 22830 21060 22836 21072
rect 22791 21032 22836 21060
rect 22830 21020 22836 21032
rect 22888 21020 22894 21072
rect 12820 20964 13216 20992
rect 14642 20952 14648 21004
rect 14700 20992 14706 21004
rect 15324 20995 15382 21001
rect 15324 20992 15336 20995
rect 14700 20964 15336 20992
rect 14700 20952 14706 20964
rect 15324 20961 15336 20964
rect 15370 20961 15382 20995
rect 18230 20992 18236 21004
rect 18191 20964 18236 20992
rect 15324 20955 15382 20961
rect 18230 20952 18236 20964
rect 18288 20952 18294 21004
rect 24648 20995 24706 21001
rect 24648 20961 24660 20995
rect 24694 20992 24706 20995
rect 25498 20992 25504 21004
rect 24694 20964 25504 20992
rect 24694 20961 24706 20964
rect 24648 20955 24706 20961
rect 25498 20952 25504 20964
rect 25556 20952 25562 21004
rect 6365 20927 6423 20933
rect 6365 20924 6377 20927
rect 6196 20896 6377 20924
rect 6196 20800 6224 20896
rect 6365 20893 6377 20896
rect 6411 20893 6423 20927
rect 6365 20887 6423 20893
rect 11241 20927 11299 20933
rect 11241 20893 11253 20927
rect 11287 20924 11299 20927
rect 12342 20924 12348 20936
rect 11287 20896 12348 20924
rect 11287 20893 11299 20896
rect 11241 20887 11299 20893
rect 12342 20884 12348 20896
rect 12400 20884 12406 20936
rect 12805 20927 12863 20933
rect 12805 20893 12817 20927
rect 12851 20924 12863 20927
rect 13446 20924 13452 20936
rect 12851 20896 13452 20924
rect 12851 20893 12863 20896
rect 12805 20887 12863 20893
rect 13446 20884 13452 20896
rect 13504 20884 13510 20936
rect 13722 20924 13728 20936
rect 13683 20896 13728 20924
rect 13722 20884 13728 20896
rect 13780 20884 13786 20936
rect 16666 20924 16672 20936
rect 16627 20896 16672 20924
rect 16666 20884 16672 20896
rect 16724 20884 16730 20936
rect 17313 20927 17371 20933
rect 17313 20893 17325 20927
rect 17359 20924 17371 20927
rect 17586 20924 17592 20936
rect 17359 20896 17592 20924
rect 17359 20893 17371 20896
rect 17313 20887 17371 20893
rect 14090 20816 14096 20868
rect 14148 20856 14154 20868
rect 14277 20859 14335 20865
rect 14277 20856 14289 20859
rect 14148 20828 14289 20856
rect 14148 20816 14154 20828
rect 14277 20825 14289 20828
rect 14323 20856 14335 20859
rect 17328 20856 17356 20887
rect 17586 20884 17592 20896
rect 17644 20884 17650 20936
rect 19337 20927 19395 20933
rect 19337 20893 19349 20927
rect 19383 20924 19395 20927
rect 19978 20924 19984 20936
rect 19383 20896 19984 20924
rect 19383 20893 19395 20896
rect 19337 20887 19395 20893
rect 19978 20884 19984 20896
rect 20036 20884 20042 20936
rect 21450 20924 21456 20936
rect 21411 20896 21456 20924
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 22738 20924 22744 20936
rect 22699 20896 22744 20924
rect 22738 20884 22744 20896
rect 22796 20884 22802 20936
rect 23017 20927 23075 20933
rect 23017 20924 23029 20927
rect 22848 20896 23029 20924
rect 14323 20828 17356 20856
rect 18371 20859 18429 20865
rect 14323 20825 14335 20828
rect 14277 20819 14335 20825
rect 18371 20825 18383 20859
rect 18417 20856 18429 20859
rect 19794 20856 19800 20868
rect 18417 20828 19800 20856
rect 18417 20825 18429 20828
rect 18371 20819 18429 20825
rect 19794 20816 19800 20828
rect 19852 20816 19858 20868
rect 19889 20859 19947 20865
rect 19889 20825 19901 20859
rect 19935 20856 19947 20859
rect 20806 20856 20812 20868
rect 19935 20828 20812 20856
rect 19935 20825 19947 20828
rect 19889 20819 19947 20825
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 22002 20816 22008 20868
rect 22060 20856 22066 20868
rect 22848 20856 22876 20896
rect 23017 20893 23029 20896
rect 23063 20893 23075 20927
rect 23017 20887 23075 20893
rect 22060 20828 22876 20856
rect 22060 20816 22066 20828
rect 5261 20791 5319 20797
rect 5261 20757 5273 20791
rect 5307 20788 5319 20791
rect 5534 20788 5540 20800
rect 5307 20760 5540 20788
rect 5307 20757 5319 20760
rect 5261 20751 5319 20757
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 6178 20788 6184 20800
rect 6139 20760 6184 20788
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 7282 20788 7288 20800
rect 7243 20760 7288 20788
rect 7282 20748 7288 20760
rect 7340 20748 7346 20800
rect 7926 20788 7932 20800
rect 7887 20760 7932 20788
rect 7926 20748 7932 20760
rect 7984 20748 7990 20800
rect 15654 20748 15660 20800
rect 15712 20788 15718 20800
rect 15749 20791 15807 20797
rect 15749 20788 15761 20791
rect 15712 20760 15761 20788
rect 15712 20748 15718 20760
rect 15749 20757 15761 20760
rect 15795 20757 15807 20791
rect 18046 20788 18052 20800
rect 18007 20760 18052 20788
rect 15749 20751 15807 20757
rect 18046 20748 18052 20760
rect 18104 20748 18110 20800
rect 18690 20788 18696 20800
rect 18651 20760 18696 20788
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 18874 20748 18880 20800
rect 18932 20788 18938 20800
rect 24719 20791 24777 20797
rect 24719 20788 24731 20791
rect 18932 20760 24731 20788
rect 18932 20748 18938 20760
rect 24719 20757 24731 20760
rect 24765 20757 24777 20791
rect 24719 20751 24777 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 7282 20544 7288 20596
rect 7340 20584 7346 20596
rect 8389 20587 8447 20593
rect 8389 20584 8401 20587
rect 7340 20556 8401 20584
rect 7340 20544 7346 20556
rect 8389 20553 8401 20556
rect 8435 20584 8447 20587
rect 8754 20584 8760 20596
rect 8435 20556 8760 20584
rect 8435 20553 8447 20556
rect 8389 20547 8447 20553
rect 8754 20544 8760 20556
rect 8812 20544 8818 20596
rect 13354 20584 13360 20596
rect 13315 20556 13360 20584
rect 13354 20544 13360 20556
rect 13412 20584 13418 20596
rect 13633 20587 13691 20593
rect 13633 20584 13645 20587
rect 13412 20556 13645 20584
rect 13412 20544 13418 20556
rect 13633 20553 13645 20556
rect 13679 20584 13691 20587
rect 14001 20587 14059 20593
rect 14001 20584 14013 20587
rect 13679 20556 14013 20584
rect 13679 20553 13691 20556
rect 13633 20547 13691 20553
rect 14001 20553 14013 20556
rect 14047 20553 14059 20587
rect 14001 20547 14059 20553
rect 14642 20544 14648 20596
rect 14700 20584 14706 20596
rect 15013 20587 15071 20593
rect 15013 20584 15025 20587
rect 14700 20556 15025 20584
rect 14700 20544 14706 20556
rect 15013 20553 15025 20556
rect 15059 20553 15071 20587
rect 15013 20547 15071 20553
rect 16666 20544 16672 20596
rect 16724 20584 16730 20596
rect 17083 20587 17141 20593
rect 17083 20584 17095 20587
rect 16724 20556 17095 20584
rect 16724 20544 16730 20556
rect 17083 20553 17095 20556
rect 17129 20553 17141 20587
rect 17083 20547 17141 20553
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 20956 20556 21465 20584
rect 20956 20544 20962 20556
rect 21453 20553 21465 20556
rect 21499 20553 21511 20587
rect 21453 20547 21511 20553
rect 22738 20544 22744 20596
rect 22796 20584 22802 20596
rect 23382 20584 23388 20596
rect 22796 20556 23388 20584
rect 22796 20544 22802 20556
rect 23382 20544 23388 20556
rect 23440 20544 23446 20596
rect 25130 20584 25136 20596
rect 25091 20556 25136 20584
rect 25130 20544 25136 20556
rect 25188 20544 25194 20596
rect 25498 20584 25504 20596
rect 25459 20556 25504 20584
rect 25498 20544 25504 20556
rect 25556 20544 25562 20596
rect 7742 20516 7748 20528
rect 7703 20488 7748 20516
rect 7742 20476 7748 20488
rect 7800 20476 7806 20528
rect 4154 20408 4160 20460
rect 4212 20448 4218 20460
rect 5905 20451 5963 20457
rect 4212 20420 4257 20448
rect 4212 20408 4218 20420
rect 5905 20417 5917 20451
rect 5951 20448 5963 20451
rect 6178 20448 6184 20460
rect 5951 20420 6184 20448
rect 5951 20417 5963 20420
rect 5905 20411 5963 20417
rect 6178 20408 6184 20420
rect 6236 20408 6242 20460
rect 8846 20408 8852 20460
rect 8904 20448 8910 20460
rect 8941 20451 8999 20457
rect 8941 20448 8953 20451
rect 8904 20420 8953 20448
rect 8904 20408 8910 20420
rect 8941 20417 8953 20420
rect 8987 20417 8999 20451
rect 10686 20448 10692 20460
rect 8941 20411 8999 20417
rect 9646 20420 10692 20448
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 5077 20383 5135 20389
rect 5077 20380 5089 20383
rect 1443 20352 2084 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2056 20256 2084 20352
rect 4126 20352 5089 20380
rect 3878 20272 3884 20324
rect 3936 20312 3942 20324
rect 4126 20312 4154 20352
rect 5077 20349 5089 20352
rect 5123 20380 5135 20383
rect 5169 20383 5227 20389
rect 5169 20380 5181 20383
rect 5123 20352 5181 20380
rect 5123 20349 5135 20352
rect 5077 20343 5135 20349
rect 5169 20349 5181 20352
rect 5215 20349 5227 20383
rect 5169 20343 5227 20349
rect 5534 20340 5540 20392
rect 5592 20380 5598 20392
rect 5629 20383 5687 20389
rect 5629 20380 5641 20383
rect 5592 20352 5641 20380
rect 5592 20340 5598 20352
rect 5629 20349 5641 20352
rect 5675 20349 5687 20383
rect 5629 20343 5687 20349
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 7650 20380 7656 20392
rect 6871 20352 7656 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 7650 20340 7656 20352
rect 7708 20380 7714 20392
rect 8021 20383 8079 20389
rect 8021 20380 8033 20383
rect 7708 20352 8033 20380
rect 7708 20340 7714 20352
rect 8021 20349 8033 20352
rect 8067 20349 8079 20383
rect 8021 20343 8079 20349
rect 6638 20312 6644 20324
rect 3936 20284 4154 20312
rect 6551 20284 6644 20312
rect 3936 20272 3942 20284
rect 6638 20272 6644 20284
rect 6696 20312 6702 20324
rect 7187 20315 7245 20321
rect 7187 20312 7199 20315
rect 6696 20284 7199 20312
rect 6696 20272 6702 20284
rect 7187 20281 7199 20284
rect 7233 20312 7245 20315
rect 7282 20312 7288 20324
rect 7233 20284 7288 20312
rect 7233 20281 7245 20284
rect 7187 20275 7245 20281
rect 7282 20272 7288 20284
rect 7340 20272 7346 20324
rect 8662 20312 8668 20324
rect 8623 20284 8668 20312
rect 8662 20272 8668 20284
rect 8720 20272 8726 20324
rect 8754 20272 8760 20324
rect 8812 20312 8818 20324
rect 8812 20284 8857 20312
rect 8812 20272 8818 20284
rect 2038 20244 2044 20256
rect 1999 20216 2044 20244
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 6273 20247 6331 20253
rect 6273 20213 6285 20247
rect 6319 20244 6331 20247
rect 6362 20244 6368 20256
rect 6319 20216 6368 20244
rect 6319 20213 6331 20216
rect 6273 20207 6331 20213
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 9646 20244 9674 20420
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 12250 20408 12256 20460
rect 12308 20448 12314 20460
rect 12308 20420 12848 20448
rect 12308 20408 12314 20420
rect 9861 20383 9919 20389
rect 9861 20349 9873 20383
rect 9907 20380 9919 20383
rect 10229 20383 10287 20389
rect 10229 20380 10241 20383
rect 9907 20352 10241 20380
rect 9907 20349 9919 20352
rect 9861 20343 9919 20349
rect 10229 20349 10241 20352
rect 10275 20380 10287 20383
rect 11054 20380 11060 20392
rect 10275 20352 11060 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 11054 20340 11060 20352
rect 11112 20340 11118 20392
rect 11241 20383 11299 20389
rect 11241 20349 11253 20383
rect 11287 20380 11299 20383
rect 11793 20383 11851 20389
rect 11793 20380 11805 20383
rect 11287 20352 11805 20380
rect 11287 20349 11299 20352
rect 11241 20343 11299 20349
rect 11793 20349 11805 20352
rect 11839 20349 11851 20383
rect 12434 20380 12440 20392
rect 12395 20352 12440 20380
rect 11793 20343 11851 20349
rect 10778 20272 10784 20324
rect 10836 20312 10842 20324
rect 11256 20312 11284 20343
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 10836 20284 11284 20312
rect 11517 20315 11575 20321
rect 10836 20272 10842 20284
rect 11517 20281 11529 20315
rect 11563 20312 11575 20315
rect 12618 20312 12624 20324
rect 11563 20284 12624 20312
rect 11563 20281 11575 20284
rect 11517 20275 11575 20281
rect 12618 20272 12624 20284
rect 12676 20272 12682 20324
rect 12820 20321 12848 20420
rect 12894 20408 12900 20460
rect 12952 20448 12958 20460
rect 14660 20448 14688 20544
rect 16117 20519 16175 20525
rect 16117 20485 16129 20519
rect 16163 20516 16175 20519
rect 16163 20488 16712 20516
rect 16163 20485 16175 20488
rect 16117 20479 16175 20485
rect 12952 20420 14688 20448
rect 15197 20451 15255 20457
rect 12952 20408 12958 20420
rect 15197 20417 15209 20451
rect 15243 20448 15255 20451
rect 15286 20448 15292 20460
rect 15243 20420 15292 20448
rect 15243 20417 15255 20420
rect 15197 20411 15255 20417
rect 15286 20408 15292 20420
rect 15344 20408 15350 20460
rect 16684 20457 16712 20488
rect 21542 20476 21548 20528
rect 21600 20516 21606 20528
rect 21600 20488 22416 20516
rect 21600 20476 21606 20488
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 16758 20448 16764 20460
rect 16715 20420 16764 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 16758 20408 16764 20420
rect 16816 20408 16822 20460
rect 17126 20448 17132 20460
rect 16868 20420 17132 20448
rect 14236 20383 14294 20389
rect 14236 20349 14248 20383
rect 14282 20380 14294 20383
rect 14645 20383 14703 20389
rect 14645 20380 14657 20383
rect 14282 20352 14657 20380
rect 14282 20349 14294 20352
rect 14236 20343 14294 20349
rect 14645 20349 14657 20352
rect 14691 20380 14703 20383
rect 16868 20380 16896 20420
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20448 18751 20451
rect 18782 20448 18788 20460
rect 18739 20420 18788 20448
rect 18739 20417 18751 20420
rect 18693 20411 18751 20417
rect 18782 20408 18788 20420
rect 18840 20408 18846 20460
rect 19794 20408 19800 20460
rect 19852 20448 19858 20460
rect 20530 20448 20536 20460
rect 19852 20420 20536 20448
rect 19852 20408 19858 20420
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 20806 20448 20812 20460
rect 20767 20420 20812 20448
rect 20806 20408 20812 20420
rect 20864 20408 20870 20460
rect 22097 20451 22155 20457
rect 22097 20417 22109 20451
rect 22143 20448 22155 20451
rect 22186 20448 22192 20460
rect 22143 20420 22192 20448
rect 22143 20417 22155 20420
rect 22097 20411 22155 20417
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 22388 20457 22416 20488
rect 22830 20476 22836 20528
rect 22888 20516 22894 20528
rect 23017 20519 23075 20525
rect 23017 20516 23029 20519
rect 22888 20488 23029 20516
rect 22888 20476 22894 20488
rect 23017 20485 23029 20488
rect 23063 20485 23075 20519
rect 23017 20479 23075 20485
rect 22373 20451 22431 20457
rect 22373 20417 22385 20451
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 14691 20352 16896 20380
rect 17012 20383 17070 20389
rect 14691 20349 14703 20352
rect 14645 20343 14703 20349
rect 17012 20349 17024 20383
rect 17058 20380 17070 20383
rect 17402 20380 17408 20392
rect 17058 20352 17408 20380
rect 17058 20349 17070 20352
rect 17012 20343 17070 20349
rect 17402 20340 17408 20352
rect 17460 20340 17466 20392
rect 19613 20383 19671 20389
rect 19613 20349 19625 20383
rect 19659 20380 19671 20383
rect 24648 20383 24706 20389
rect 19659 20352 20392 20380
rect 19659 20349 19671 20352
rect 19613 20343 19671 20349
rect 12799 20315 12857 20321
rect 12799 20281 12811 20315
rect 12845 20281 12857 20315
rect 12799 20275 12857 20281
rect 7524 20216 9674 20244
rect 10597 20247 10655 20253
rect 7524 20204 7530 20216
rect 10597 20213 10609 20247
rect 10643 20244 10655 20247
rect 10686 20244 10692 20256
rect 10643 20216 10692 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 10686 20204 10692 20216
rect 10744 20244 10750 20256
rect 11974 20244 11980 20256
rect 10744 20216 11980 20244
rect 10744 20204 10750 20216
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 12250 20244 12256 20256
rect 12211 20216 12256 20244
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 12820 20244 12848 20275
rect 13722 20272 13728 20324
rect 13780 20312 13786 20324
rect 14323 20315 14381 20321
rect 14323 20312 14335 20315
rect 13780 20284 14335 20312
rect 13780 20272 13786 20284
rect 14323 20281 14335 20284
rect 14369 20281 14381 20315
rect 14323 20275 14381 20281
rect 15559 20315 15617 20321
rect 15559 20281 15571 20315
rect 15605 20312 15617 20315
rect 15654 20312 15660 20324
rect 15605 20284 15660 20312
rect 15605 20281 15617 20284
rect 15559 20275 15617 20281
rect 15654 20272 15660 20284
rect 15712 20272 15718 20324
rect 18690 20272 18696 20324
rect 18748 20312 18754 20324
rect 20364 20321 20392 20352
rect 24648 20349 24660 20383
rect 24694 20380 24706 20383
rect 25130 20380 25136 20392
rect 24694 20352 25136 20380
rect 24694 20349 24706 20352
rect 24648 20343 24706 20349
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 19014 20315 19072 20321
rect 19014 20312 19026 20315
rect 18748 20284 19026 20312
rect 18748 20272 18754 20284
rect 19014 20281 19026 20284
rect 19060 20281 19072 20315
rect 19014 20275 19072 20281
rect 20349 20315 20407 20321
rect 20349 20281 20361 20315
rect 20395 20312 20407 20315
rect 20622 20312 20628 20324
rect 20395 20284 20628 20312
rect 20395 20281 20407 20284
rect 20349 20275 20407 20281
rect 20622 20272 20628 20284
rect 20680 20272 20686 20324
rect 21913 20315 21971 20321
rect 21913 20281 21925 20315
rect 21959 20312 21971 20315
rect 22189 20315 22247 20321
rect 22189 20312 22201 20315
rect 21959 20284 22201 20312
rect 21959 20281 21971 20284
rect 21913 20275 21971 20281
rect 22189 20281 22201 20284
rect 22235 20312 22247 20315
rect 22278 20312 22284 20324
rect 22235 20284 22284 20312
rect 22235 20281 22247 20284
rect 22189 20275 22247 20281
rect 22278 20272 22284 20284
rect 22336 20272 22342 20324
rect 14458 20244 14464 20256
rect 12820 20216 14464 20244
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 15838 20204 15844 20256
rect 15896 20244 15902 20256
rect 17310 20244 17316 20256
rect 15896 20216 17316 20244
rect 15896 20204 15902 20216
rect 17310 20204 17316 20216
rect 17368 20244 17374 20256
rect 18230 20244 18236 20256
rect 17368 20216 18236 20244
rect 17368 20204 17374 20216
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19981 20247 20039 20253
rect 19981 20244 19993 20247
rect 19576 20216 19993 20244
rect 19576 20204 19582 20216
rect 19981 20213 19993 20216
rect 20027 20244 20039 20247
rect 21358 20244 21364 20256
rect 20027 20216 21364 20244
rect 20027 20213 20039 20216
rect 19981 20207 20039 20213
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 23106 20204 23112 20256
rect 23164 20244 23170 20256
rect 24719 20247 24777 20253
rect 24719 20244 24731 20247
rect 23164 20216 24731 20244
rect 23164 20204 23170 20216
rect 24719 20213 24731 20216
rect 24765 20213 24777 20247
rect 24719 20207 24777 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1578 20040 1584 20052
rect 1539 20012 1584 20040
rect 1578 20000 1584 20012
rect 1636 20000 1642 20052
rect 7650 20040 7656 20052
rect 7611 20012 7656 20040
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 8478 20000 8484 20052
rect 8536 20040 8542 20052
rect 8573 20043 8631 20049
rect 8573 20040 8585 20043
rect 8536 20012 8585 20040
rect 8536 20000 8542 20012
rect 8573 20009 8585 20012
rect 8619 20009 8631 20043
rect 8573 20003 8631 20009
rect 6175 19975 6233 19981
rect 6175 19941 6187 19975
rect 6221 19972 6233 19975
rect 7469 19975 7527 19981
rect 6221 19944 7144 19972
rect 6221 19941 6233 19944
rect 6175 19935 6233 19941
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 1946 19904 1952 19916
rect 1443 19876 1952 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 1946 19864 1952 19876
rect 2004 19864 2010 19916
rect 4868 19907 4926 19913
rect 4868 19873 4880 19907
rect 4914 19904 4926 19907
rect 4982 19904 4988 19916
rect 4914 19876 4988 19904
rect 4914 19873 4926 19876
rect 4868 19867 4926 19873
rect 4982 19864 4988 19876
rect 5040 19864 5046 19916
rect 7116 19913 7144 19944
rect 7469 19941 7481 19975
rect 7515 19972 7527 19975
rect 7742 19972 7748 19984
rect 7515 19944 7748 19972
rect 7515 19941 7527 19944
rect 7469 19935 7527 19941
rect 7742 19932 7748 19944
rect 7800 19932 7806 19984
rect 8588 19972 8616 20003
rect 8662 20000 8668 20052
rect 8720 20040 8726 20052
rect 8941 20043 8999 20049
rect 8941 20040 8953 20043
rect 8720 20012 8953 20040
rect 8720 20000 8726 20012
rect 8941 20009 8953 20012
rect 8987 20009 8999 20043
rect 8941 20003 8999 20009
rect 12158 20000 12164 20052
rect 12216 20040 12222 20052
rect 12253 20043 12311 20049
rect 12253 20040 12265 20043
rect 12216 20012 12265 20040
rect 12216 20000 12222 20012
rect 12253 20009 12265 20012
rect 12299 20009 12311 20043
rect 12802 20040 12808 20052
rect 12763 20012 12808 20040
rect 12253 20003 12311 20009
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 13541 20043 13599 20049
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 13722 20040 13728 20052
rect 13587 20012 13728 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 15105 20043 15163 20049
rect 15105 20009 15117 20043
rect 15151 20040 15163 20043
rect 15286 20040 15292 20052
rect 15151 20012 15292 20040
rect 15151 20009 15163 20012
rect 15105 20003 15163 20009
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 16666 20000 16672 20052
rect 16724 20040 16730 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 16724 20012 16865 20040
rect 16724 20000 16730 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 19518 20040 19524 20052
rect 19479 20012 19524 20040
rect 16853 20003 16911 20009
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 19889 20043 19947 20049
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 19978 20040 19984 20052
rect 19935 20012 19984 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 19978 20000 19984 20012
rect 20036 20000 20042 20052
rect 20530 20040 20536 20052
rect 20491 20012 20536 20040
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 23983 20043 24041 20049
rect 23983 20040 23995 20043
rect 23440 20012 23995 20040
rect 23440 20000 23446 20012
rect 23983 20009 23995 20012
rect 24029 20009 24041 20043
rect 23983 20003 24041 20009
rect 11974 19972 11980 19984
rect 8588 19944 11980 19972
rect 11974 19932 11980 19944
rect 12032 19932 12038 19984
rect 13817 19975 13875 19981
rect 13817 19972 13829 19975
rect 13556 19944 13829 19972
rect 13556 19916 13584 19944
rect 13817 19941 13829 19944
rect 13863 19941 13875 19975
rect 13817 19935 13875 19941
rect 13906 19932 13912 19984
rect 13964 19972 13970 19984
rect 14369 19975 14427 19981
rect 14369 19972 14381 19975
rect 13964 19944 14381 19972
rect 13964 19932 13970 19944
rect 14369 19941 14381 19944
rect 14415 19941 14427 19975
rect 14369 19935 14427 19941
rect 15470 19932 15476 19984
rect 15528 19972 15534 19984
rect 15654 19981 15660 19984
rect 15610 19975 15660 19981
rect 15610 19972 15622 19975
rect 15528 19944 15622 19972
rect 15528 19932 15534 19944
rect 15610 19941 15622 19944
rect 15656 19941 15660 19975
rect 15610 19935 15660 19941
rect 15654 19932 15660 19935
rect 15712 19932 15718 19984
rect 16022 19932 16028 19984
rect 16080 19972 16086 19984
rect 16577 19975 16635 19981
rect 16577 19972 16589 19975
rect 16080 19944 16589 19972
rect 16080 19932 16086 19944
rect 16577 19941 16589 19944
rect 16623 19972 16635 19975
rect 16758 19972 16764 19984
rect 16623 19944 16764 19972
rect 16623 19941 16635 19944
rect 16577 19935 16635 19941
rect 16758 19932 16764 19944
rect 16816 19932 16822 19984
rect 17218 19972 17224 19984
rect 17179 19944 17224 19972
rect 17218 19932 17224 19944
rect 17276 19932 17282 19984
rect 18690 19932 18696 19984
rect 18748 19972 18754 19984
rect 18922 19975 18980 19981
rect 18922 19972 18934 19975
rect 18748 19944 18934 19972
rect 18748 19932 18754 19944
rect 18922 19941 18934 19944
rect 18968 19941 18980 19975
rect 18922 19935 18980 19941
rect 21177 19975 21235 19981
rect 21177 19941 21189 19975
rect 21223 19972 21235 19975
rect 21358 19972 21364 19984
rect 21223 19944 21364 19972
rect 21223 19941 21235 19944
rect 21177 19935 21235 19941
rect 21358 19932 21364 19944
rect 21416 19972 21422 19984
rect 21453 19975 21511 19981
rect 21453 19972 21465 19975
rect 21416 19944 21465 19972
rect 21416 19932 21422 19944
rect 21453 19941 21465 19944
rect 21499 19972 21511 19975
rect 22094 19972 22100 19984
rect 21499 19944 22100 19972
rect 21499 19941 21511 19944
rect 21453 19935 21511 19941
rect 22094 19932 22100 19944
rect 22152 19932 22158 19984
rect 7101 19907 7159 19913
rect 7101 19873 7113 19907
rect 7147 19904 7159 19907
rect 7282 19904 7288 19916
rect 7147 19876 7288 19904
rect 7147 19873 7159 19876
rect 7101 19867 7159 19873
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 7837 19907 7895 19913
rect 7837 19873 7849 19907
rect 7883 19904 7895 19907
rect 7926 19904 7932 19916
rect 7883 19876 7932 19904
rect 7883 19873 7895 19876
rect 7837 19867 7895 19873
rect 7926 19864 7932 19876
rect 7984 19864 7990 19916
rect 8021 19907 8079 19913
rect 8021 19873 8033 19907
rect 8067 19873 8079 19907
rect 10318 19904 10324 19916
rect 10279 19876 10324 19904
rect 8021 19867 8079 19873
rect 5813 19839 5871 19845
rect 5813 19805 5825 19839
rect 5859 19836 5871 19839
rect 5994 19836 6000 19848
rect 5859 19808 6000 19836
rect 5859 19805 5871 19808
rect 5813 19799 5871 19805
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 7190 19796 7196 19848
rect 7248 19836 7254 19848
rect 8036 19836 8064 19867
rect 10318 19864 10324 19876
rect 10376 19904 10382 19916
rect 10778 19904 10784 19916
rect 10376 19876 10784 19904
rect 10376 19864 10382 19876
rect 10778 19864 10784 19876
rect 10836 19864 10842 19916
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19873 10931 19907
rect 10873 19867 10931 19873
rect 7248 19808 8064 19836
rect 7248 19796 7254 19808
rect 4062 19728 4068 19780
rect 4120 19768 4126 19780
rect 5261 19771 5319 19777
rect 5261 19768 5273 19771
rect 4120 19740 5273 19768
rect 4120 19728 4126 19740
rect 5261 19737 5273 19740
rect 5307 19737 5319 19771
rect 5261 19731 5319 19737
rect 6733 19771 6791 19777
rect 6733 19737 6745 19771
rect 6779 19768 6791 19771
rect 7098 19768 7104 19780
rect 6779 19740 7104 19768
rect 6779 19737 6791 19740
rect 6733 19731 6791 19737
rect 7098 19728 7104 19740
rect 7156 19768 7162 19780
rect 8386 19768 8392 19780
rect 7156 19740 8392 19768
rect 7156 19728 7162 19740
rect 8386 19728 8392 19740
rect 8444 19728 8450 19780
rect 10888 19768 10916 19867
rect 13538 19864 13544 19916
rect 13596 19864 13602 19916
rect 22002 19864 22008 19916
rect 22060 19904 22066 19916
rect 22830 19904 22836 19916
rect 22060 19876 22105 19904
rect 22791 19876 22836 19904
rect 22060 19864 22066 19876
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 23912 19907 23970 19913
rect 23912 19873 23924 19907
rect 23958 19904 23970 19907
rect 24210 19904 24216 19916
rect 23958 19876 24216 19904
rect 23958 19873 23970 19876
rect 23912 19867 23970 19873
rect 24210 19864 24216 19876
rect 24268 19864 24274 19916
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19836 11115 19839
rect 11882 19836 11888 19848
rect 11103 19808 11888 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 13725 19839 13783 19845
rect 13725 19836 13737 19839
rect 13504 19808 13737 19836
rect 13504 19796 13510 19808
rect 13725 19805 13737 19808
rect 13771 19836 13783 19839
rect 13998 19836 14004 19848
rect 13771 19808 14004 19836
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 13998 19796 14004 19808
rect 14056 19796 14062 19848
rect 15286 19836 15292 19848
rect 15247 19808 15292 19836
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 17129 19839 17187 19845
rect 17129 19805 17141 19839
rect 17175 19836 17187 19839
rect 17494 19836 17500 19848
rect 17175 19808 17500 19836
rect 17175 19805 17187 19808
rect 17129 19799 17187 19805
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 17586 19796 17592 19848
rect 17644 19836 17650 19848
rect 18598 19836 18604 19848
rect 17644 19808 17689 19836
rect 18559 19808 18604 19836
rect 17644 19796 17650 19808
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 20622 19796 20628 19848
rect 20680 19836 20686 19848
rect 21361 19839 21419 19845
rect 21361 19836 21373 19839
rect 20680 19808 21373 19836
rect 20680 19796 20686 19808
rect 21361 19805 21373 19808
rect 21407 19836 21419 19839
rect 23106 19836 23112 19848
rect 21407 19808 23112 19836
rect 21407 19805 21419 19808
rect 21361 19799 21419 19805
rect 23106 19796 23112 19808
rect 23164 19796 23170 19848
rect 11330 19768 11336 19780
rect 10888 19740 11336 19768
rect 11330 19728 11336 19740
rect 11388 19768 11394 19780
rect 11425 19771 11483 19777
rect 11425 19768 11437 19771
rect 11388 19740 11437 19768
rect 11388 19728 11394 19740
rect 11425 19737 11437 19740
rect 11471 19768 11483 19771
rect 14182 19768 14188 19780
rect 11471 19740 13216 19768
rect 11471 19737 11483 19740
rect 11425 19731 11483 19737
rect 3602 19700 3608 19712
rect 3563 19672 3608 19700
rect 3602 19660 3608 19672
rect 3660 19660 3666 19712
rect 4939 19703 4997 19709
rect 4939 19669 4951 19703
rect 4985 19700 4997 19703
rect 5442 19700 5448 19712
rect 4985 19672 5448 19700
rect 4985 19669 4997 19672
rect 4939 19663 4997 19669
rect 5442 19660 5448 19672
rect 5500 19660 5506 19712
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 5629 19703 5687 19709
rect 5629 19700 5641 19703
rect 5592 19672 5641 19700
rect 5592 19660 5598 19672
rect 5629 19669 5641 19672
rect 5675 19669 5687 19703
rect 5629 19663 5687 19669
rect 11514 19660 11520 19712
rect 11572 19700 11578 19712
rect 12434 19700 12440 19712
rect 11572 19672 12440 19700
rect 11572 19660 11578 19672
rect 12434 19660 12440 19672
rect 12492 19700 12498 19712
rect 13081 19703 13139 19709
rect 13081 19700 13093 19703
rect 12492 19672 13093 19700
rect 12492 19660 12498 19672
rect 13081 19669 13093 19672
rect 13127 19669 13139 19703
rect 13188 19700 13216 19740
rect 13786 19740 14188 19768
rect 13786 19712 13814 19740
rect 14182 19728 14188 19740
rect 14240 19728 14246 19780
rect 14734 19728 14740 19780
rect 14792 19768 14798 19780
rect 18874 19768 18880 19780
rect 14792 19740 18880 19768
rect 14792 19728 14798 19740
rect 18874 19728 18880 19740
rect 18932 19728 18938 19780
rect 13722 19700 13728 19712
rect 13188 19672 13728 19700
rect 13081 19663 13139 19669
rect 13722 19660 13728 19672
rect 13780 19672 13814 19712
rect 13780 19660 13786 19672
rect 15930 19660 15936 19712
rect 15988 19700 15994 19712
rect 16209 19703 16267 19709
rect 16209 19700 16221 19703
rect 15988 19672 16221 19700
rect 15988 19660 15994 19672
rect 16209 19669 16221 19672
rect 16255 19669 16267 19703
rect 16209 19663 16267 19669
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 22971 19703 23029 19709
rect 22971 19700 22983 19703
rect 19392 19672 22983 19700
rect 19392 19660 19398 19672
rect 22971 19669 22983 19672
rect 23017 19669 23029 19703
rect 22971 19663 23029 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2038 19456 2044 19508
rect 2096 19496 2102 19508
rect 2639 19499 2697 19505
rect 2639 19496 2651 19499
rect 2096 19468 2651 19496
rect 2096 19456 2102 19468
rect 2639 19465 2651 19468
rect 2685 19465 2697 19499
rect 4893 19499 4951 19505
rect 4893 19496 4905 19499
rect 2639 19459 2697 19465
rect 4126 19468 4905 19496
rect 3970 19320 3976 19372
rect 4028 19360 4034 19372
rect 4126 19360 4154 19468
rect 4893 19465 4905 19468
rect 4939 19496 4951 19499
rect 4982 19496 4988 19508
rect 4939 19468 4988 19496
rect 4939 19465 4951 19468
rect 4893 19459 4951 19465
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 8202 19456 8208 19508
rect 8260 19496 8266 19508
rect 10318 19496 10324 19508
rect 8260 19468 10324 19496
rect 8260 19456 8266 19468
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 13814 19496 13820 19508
rect 11756 19468 13820 19496
rect 11756 19456 11762 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 14458 19456 14464 19508
rect 14516 19496 14522 19508
rect 15289 19499 15347 19505
rect 15289 19496 15301 19499
rect 14516 19468 15301 19496
rect 14516 19456 14522 19468
rect 15289 19465 15301 19468
rect 15335 19496 15347 19499
rect 15470 19496 15476 19508
rect 15335 19468 15476 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 15562 19456 15568 19508
rect 15620 19496 15626 19508
rect 15657 19499 15715 19505
rect 15657 19496 15669 19499
rect 15620 19468 15669 19496
rect 15620 19456 15626 19468
rect 15657 19465 15669 19468
rect 15703 19465 15715 19499
rect 15657 19459 15715 19465
rect 6270 19388 6276 19440
rect 6328 19428 6334 19440
rect 9953 19431 10011 19437
rect 9953 19428 9965 19431
rect 6328 19400 9965 19428
rect 6328 19388 6334 19400
rect 9953 19397 9965 19400
rect 9999 19397 10011 19431
rect 9953 19391 10011 19397
rect 4028 19332 4154 19360
rect 5905 19363 5963 19369
rect 4028 19320 4034 19332
rect 5905 19329 5917 19363
rect 5951 19360 5963 19363
rect 5994 19360 6000 19372
rect 5951 19332 6000 19360
rect 5951 19329 5963 19332
rect 5905 19323 5963 19329
rect 5994 19320 6000 19332
rect 6052 19360 6058 19372
rect 6549 19363 6607 19369
rect 6549 19360 6561 19363
rect 6052 19332 6561 19360
rect 6052 19320 6058 19332
rect 6549 19329 6561 19332
rect 6595 19329 6607 19363
rect 7374 19360 7380 19372
rect 7335 19332 7380 19360
rect 6549 19323 6607 19329
rect 7374 19320 7380 19332
rect 7432 19320 7438 19372
rect 7834 19360 7840 19372
rect 7795 19332 7840 19360
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 8294 19320 8300 19372
rect 8352 19360 8358 19372
rect 9214 19360 9220 19372
rect 8352 19332 9220 19360
rect 8352 19320 8358 19332
rect 9214 19320 9220 19332
rect 9272 19320 9278 19372
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1670 19292 1676 19304
rect 1443 19264 1676 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 2568 19295 2626 19301
rect 2568 19261 2580 19295
rect 2614 19292 2626 19295
rect 2961 19295 3019 19301
rect 2961 19292 2973 19295
rect 2614 19264 2973 19292
rect 2614 19261 2626 19264
rect 2568 19255 2626 19261
rect 2961 19261 2973 19264
rect 3007 19292 3019 19295
rect 3418 19292 3424 19304
rect 3007 19264 3424 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 3418 19252 3424 19264
rect 3476 19252 3482 19304
rect 3602 19292 3608 19304
rect 3563 19264 3608 19292
rect 3602 19252 3608 19264
rect 3660 19252 3666 19304
rect 3694 19252 3700 19304
rect 3752 19292 3758 19304
rect 3881 19295 3939 19301
rect 3752 19264 3797 19292
rect 3752 19252 3758 19264
rect 3881 19261 3893 19295
rect 3927 19261 3939 19295
rect 3881 19255 3939 19261
rect 3896 19224 3924 19255
rect 4062 19252 4068 19304
rect 4120 19292 4126 19304
rect 5166 19292 5172 19304
rect 4120 19264 5172 19292
rect 4120 19252 4126 19264
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5258 19252 5264 19304
rect 5316 19292 5322 19304
rect 5534 19292 5540 19304
rect 5316 19264 5540 19292
rect 5316 19252 5322 19264
rect 5534 19252 5540 19264
rect 5592 19292 5598 19304
rect 5629 19295 5687 19301
rect 5629 19292 5641 19295
rect 5592 19264 5641 19292
rect 5592 19252 5598 19264
rect 5629 19261 5641 19264
rect 5675 19292 5687 19295
rect 7101 19295 7159 19301
rect 7101 19292 7113 19295
rect 5675 19264 7113 19292
rect 5675 19261 5687 19264
rect 5629 19255 5687 19261
rect 7101 19261 7113 19264
rect 7147 19292 7159 19295
rect 7190 19292 7196 19304
rect 7147 19264 7196 19292
rect 7147 19261 7159 19264
rect 7101 19255 7159 19261
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 9968 19292 9996 19391
rect 11514 19360 11520 19372
rect 11475 19332 11520 19360
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 13633 19363 13691 19369
rect 13633 19360 13645 19363
rect 12452 19332 13645 19360
rect 10781 19295 10839 19301
rect 10781 19292 10793 19295
rect 9968 19264 10793 19292
rect 10781 19261 10793 19264
rect 10827 19261 10839 19295
rect 11330 19292 11336 19304
rect 11291 19264 11336 19292
rect 10781 19255 10839 19261
rect 11330 19252 11336 19264
rect 11388 19252 11394 19304
rect 12250 19252 12256 19304
rect 12308 19292 12314 19304
rect 12452 19301 12480 19332
rect 13633 19329 13645 19332
rect 13679 19329 13691 19363
rect 13832 19360 13860 19456
rect 14553 19363 14611 19369
rect 14553 19360 14565 19363
rect 13832 19332 14565 19360
rect 13633 19323 13691 19329
rect 14553 19329 14565 19332
rect 14599 19329 14611 19363
rect 15672 19360 15700 19459
rect 15930 19456 15936 19508
rect 15988 19496 15994 19508
rect 17037 19499 17095 19505
rect 17037 19496 17049 19499
rect 15988 19468 17049 19496
rect 15988 19456 15994 19468
rect 17037 19465 17049 19468
rect 17083 19496 17095 19499
rect 17218 19496 17224 19508
rect 17083 19468 17224 19496
rect 17083 19465 17095 19468
rect 17037 19459 17095 19465
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 17865 19499 17923 19505
rect 17865 19465 17877 19499
rect 17911 19496 17923 19499
rect 18598 19496 18604 19508
rect 17911 19468 18604 19496
rect 17911 19465 17923 19468
rect 17865 19459 17923 19465
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 20622 19496 20628 19508
rect 20583 19468 20628 19496
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 22094 19496 22100 19508
rect 22055 19468 22100 19496
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 17402 19388 17408 19440
rect 17460 19428 17466 19440
rect 24210 19428 24216 19440
rect 17460 19400 24216 19428
rect 17460 19388 17466 19400
rect 24210 19388 24216 19400
rect 24268 19388 24274 19440
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15672 19332 15945 19360
rect 14553 19323 14611 19329
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 18601 19363 18659 19369
rect 18601 19360 18613 19363
rect 15933 19323 15991 19329
rect 17236 19332 18613 19360
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12308 19264 12449 19292
rect 12308 19252 12314 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 13357 19295 13415 19301
rect 13357 19261 13369 19295
rect 13403 19292 13415 19295
rect 14001 19295 14059 19301
rect 14001 19292 14013 19295
rect 13403 19264 14013 19292
rect 13403 19261 13415 19264
rect 13357 19255 13415 19261
rect 14001 19261 14013 19264
rect 14047 19261 14059 19295
rect 14001 19255 14059 19261
rect 4338 19224 4344 19236
rect 3436 19196 3924 19224
rect 4299 19196 4344 19224
rect 106 19116 112 19168
rect 164 19156 170 19168
rect 1581 19159 1639 19165
rect 1581 19156 1593 19159
rect 164 19128 1593 19156
rect 164 19116 170 19128
rect 1581 19125 1593 19128
rect 1627 19125 1639 19159
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1581 19119 1639 19125
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 3050 19116 3056 19168
rect 3108 19156 3114 19168
rect 3436 19165 3464 19196
rect 4338 19184 4344 19196
rect 4396 19184 4402 19236
rect 7469 19227 7527 19233
rect 7469 19193 7481 19227
rect 7515 19224 7527 19227
rect 7742 19224 7748 19236
rect 7515 19196 7748 19224
rect 7515 19193 7527 19196
rect 7469 19187 7527 19193
rect 7742 19184 7748 19196
rect 7800 19184 7806 19236
rect 8938 19224 8944 19236
rect 8899 19196 8944 19224
rect 8938 19184 8944 19196
rect 8996 19184 9002 19236
rect 9033 19227 9091 19233
rect 9033 19193 9045 19227
rect 9079 19193 9091 19227
rect 12710 19224 12716 19236
rect 12671 19196 12716 19224
rect 9033 19187 9091 19193
rect 3421 19159 3479 19165
rect 3421 19156 3433 19159
rect 3108 19128 3433 19156
rect 3108 19116 3114 19128
rect 3421 19125 3433 19128
rect 3467 19125 3479 19159
rect 3421 19119 3479 19125
rect 6273 19159 6331 19165
rect 6273 19125 6285 19159
rect 6319 19156 6331 19159
rect 6454 19156 6460 19168
rect 6319 19128 6460 19156
rect 6319 19125 6331 19128
rect 6273 19119 6331 19125
rect 6454 19116 6460 19128
rect 6512 19156 6518 19168
rect 7282 19156 7288 19168
rect 6512 19128 7288 19156
rect 6512 19116 6518 19128
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 7926 19116 7932 19168
rect 7984 19156 7990 19168
rect 8297 19159 8355 19165
rect 8297 19156 8309 19159
rect 7984 19128 8309 19156
rect 7984 19116 7990 19128
rect 8297 19125 8309 19128
rect 8343 19125 8355 19159
rect 8297 19119 8355 19125
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 8757 19159 8815 19165
rect 8757 19156 8769 19159
rect 8444 19128 8769 19156
rect 8444 19116 8450 19128
rect 8757 19125 8769 19128
rect 8803 19156 8815 19159
rect 9048 19156 9076 19187
rect 12710 19184 12716 19196
rect 12768 19184 12774 19236
rect 8803 19128 9076 19156
rect 11885 19159 11943 19165
rect 8803 19125 8815 19128
rect 8757 19119 8815 19125
rect 11885 19125 11897 19159
rect 11931 19156 11943 19159
rect 12158 19156 12164 19168
rect 11931 19128 12164 19156
rect 11931 19125 11943 19128
rect 11885 19119 11943 19125
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 14016 19156 14044 19255
rect 14090 19184 14096 19236
rect 14148 19224 14154 19236
rect 14277 19227 14335 19233
rect 14277 19224 14289 19227
rect 14148 19196 14289 19224
rect 14148 19184 14154 19196
rect 14277 19193 14289 19196
rect 14323 19193 14335 19227
rect 14277 19187 14335 19193
rect 14369 19227 14427 19233
rect 14369 19193 14381 19227
rect 14415 19193 14427 19227
rect 16022 19224 16028 19236
rect 15983 19196 16028 19224
rect 14369 19187 14427 19193
rect 14384 19156 14412 19187
rect 16022 19184 16028 19196
rect 16080 19184 16086 19236
rect 16574 19224 16580 19236
rect 16535 19196 16580 19224
rect 16574 19184 16580 19196
rect 16632 19184 16638 19236
rect 14016 19128 14412 19156
rect 15470 19116 15476 19168
rect 15528 19156 15534 19168
rect 17236 19156 17264 19332
rect 18601 19329 18613 19332
rect 18647 19360 18659 19363
rect 18690 19360 18696 19372
rect 18647 19332 18696 19360
rect 18647 19329 18659 19332
rect 18601 19323 18659 19329
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 19978 19320 19984 19372
rect 20036 19360 20042 19372
rect 20257 19363 20315 19369
rect 20257 19360 20269 19363
rect 20036 19332 20269 19360
rect 20036 19320 20042 19332
rect 20257 19329 20269 19332
rect 20303 19360 20315 19363
rect 21177 19363 21235 19369
rect 21177 19360 21189 19363
rect 20303 19332 21189 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 21177 19329 21189 19332
rect 21223 19360 21235 19363
rect 22002 19360 22008 19372
rect 21223 19332 22008 19360
rect 21223 19329 21235 19332
rect 21177 19323 21235 19329
rect 22002 19320 22008 19332
rect 22060 19320 22066 19372
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 18248 19264 18889 19292
rect 18248 19168 18276 19264
rect 18877 19261 18889 19264
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 18690 19184 18696 19236
rect 18748 19224 18754 19236
rect 19198 19227 19256 19233
rect 19198 19224 19210 19227
rect 18748 19196 19210 19224
rect 18748 19184 18754 19196
rect 19198 19193 19210 19196
rect 19244 19193 19256 19227
rect 19198 19187 19256 19193
rect 21266 19184 21272 19236
rect 21324 19224 21330 19236
rect 21821 19227 21879 19233
rect 21324 19196 21369 19224
rect 21324 19184 21330 19196
rect 21821 19193 21833 19227
rect 21867 19224 21879 19227
rect 22002 19224 22008 19236
rect 21867 19196 22008 19224
rect 21867 19193 21879 19196
rect 21821 19187 21879 19193
rect 22002 19184 22008 19196
rect 22060 19184 22066 19236
rect 17494 19156 17500 19168
rect 15528 19128 17264 19156
rect 17455 19128 17500 19156
rect 15528 19116 15534 19128
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 18230 19156 18236 19168
rect 18191 19128 18236 19156
rect 18230 19116 18236 19128
rect 18288 19116 18294 19168
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 19797 19159 19855 19165
rect 19797 19156 19809 19159
rect 19484 19128 19809 19156
rect 19484 19116 19490 19128
rect 19797 19125 19809 19128
rect 19843 19156 19855 19159
rect 20530 19156 20536 19168
rect 19843 19128 20536 19156
rect 19843 19125 19855 19128
rect 19797 19119 19855 19125
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 20993 19159 21051 19165
rect 20993 19125 21005 19159
rect 21039 19156 21051 19159
rect 21284 19156 21312 19184
rect 22830 19156 22836 19168
rect 21039 19128 21312 19156
rect 22791 19128 22836 19156
rect 21039 19125 21051 19128
rect 20993 19119 21051 19125
rect 22830 19116 22836 19128
rect 22888 19116 22894 19168
rect 23937 19159 23995 19165
rect 23937 19125 23949 19159
rect 23983 19156 23995 19159
rect 24210 19156 24216 19168
rect 23983 19128 24216 19156
rect 23983 19125 23995 19128
rect 23937 19119 23995 19125
rect 24210 19116 24216 19128
rect 24268 19116 24274 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1670 18952 1676 18964
rect 1631 18924 1676 18952
rect 1670 18912 1676 18924
rect 1728 18912 1734 18964
rect 7374 18912 7380 18964
rect 7432 18952 7438 18964
rect 7561 18955 7619 18961
rect 7561 18952 7573 18955
rect 7432 18924 7573 18952
rect 7432 18912 7438 18924
rect 7561 18921 7573 18924
rect 7607 18921 7619 18955
rect 8938 18952 8944 18964
rect 8899 18924 8944 18952
rect 7561 18915 7619 18921
rect 8938 18912 8944 18924
rect 8996 18912 9002 18964
rect 11882 18952 11888 18964
rect 11843 18924 11888 18952
rect 11882 18912 11888 18924
rect 11940 18912 11946 18964
rect 12158 18912 12164 18964
rect 12216 18952 12222 18964
rect 12710 18952 12716 18964
rect 12216 18924 12716 18952
rect 12216 18912 12222 18924
rect 6454 18844 6460 18896
rect 6512 18884 6518 18896
rect 6686 18887 6744 18893
rect 6686 18884 6698 18887
rect 6512 18856 6698 18884
rect 6512 18844 6518 18856
rect 6686 18853 6698 18856
rect 6732 18853 6744 18887
rect 6686 18847 6744 18853
rect 11241 18887 11299 18893
rect 11241 18853 11253 18887
rect 11287 18884 11299 18887
rect 12250 18884 12256 18896
rect 11287 18856 12256 18884
rect 11287 18853 11299 18856
rect 11241 18847 11299 18853
rect 12250 18844 12256 18856
rect 12308 18844 12314 18896
rect 12446 18893 12474 18924
rect 12710 18912 12716 18924
rect 12768 18912 12774 18964
rect 12989 18955 13047 18961
rect 12989 18921 13001 18955
rect 13035 18952 13047 18955
rect 13538 18952 13544 18964
rect 13035 18924 13544 18952
rect 13035 18921 13047 18924
rect 12989 18915 13047 18921
rect 13538 18912 13544 18924
rect 13596 18952 13602 18964
rect 13633 18955 13691 18961
rect 13633 18952 13645 18955
rect 13596 18924 13645 18952
rect 13596 18912 13602 18924
rect 13633 18921 13645 18924
rect 13679 18921 13691 18955
rect 13998 18952 14004 18964
rect 13959 18924 14004 18952
rect 13633 18915 13691 18921
rect 13998 18912 14004 18924
rect 14056 18952 14062 18964
rect 16574 18952 16580 18964
rect 14056 18924 16580 18952
rect 14056 18912 14062 18924
rect 12431 18887 12489 18893
rect 12431 18853 12443 18887
rect 12477 18853 12489 18887
rect 12431 18847 12489 18853
rect 14090 18844 14096 18896
rect 14148 18884 14154 18896
rect 14645 18887 14703 18893
rect 14645 18884 14657 18887
rect 14148 18856 14657 18884
rect 14148 18844 14154 18856
rect 14645 18853 14657 18856
rect 14691 18853 14703 18887
rect 15930 18884 15936 18896
rect 15891 18856 15936 18884
rect 14645 18847 14703 18853
rect 15930 18844 15936 18856
rect 15988 18844 15994 18896
rect 16500 18893 16528 18924
rect 16574 18912 16580 18924
rect 16632 18912 16638 18964
rect 18690 18912 18696 18964
rect 18748 18952 18754 18964
rect 18877 18955 18935 18961
rect 18877 18952 18889 18955
rect 18748 18924 18889 18952
rect 18748 18912 18754 18924
rect 18877 18921 18889 18924
rect 18923 18921 18935 18955
rect 18877 18915 18935 18921
rect 16485 18887 16543 18893
rect 16485 18853 16497 18887
rect 16531 18853 16543 18887
rect 16485 18847 16543 18853
rect 18417 18887 18475 18893
rect 18417 18853 18429 18887
rect 18463 18884 18475 18887
rect 18598 18884 18604 18896
rect 18463 18856 18604 18884
rect 18463 18853 18475 18856
rect 18417 18847 18475 18853
rect 18598 18844 18604 18856
rect 18656 18844 18662 18896
rect 19426 18884 19432 18896
rect 19387 18856 19432 18884
rect 19426 18844 19432 18856
rect 19484 18844 19490 18896
rect 19978 18884 19984 18896
rect 19939 18856 19984 18884
rect 19978 18844 19984 18856
rect 20036 18844 20042 18896
rect 21545 18887 21603 18893
rect 21545 18853 21557 18887
rect 21591 18884 21603 18887
rect 22186 18884 22192 18896
rect 21591 18856 22192 18884
rect 21591 18853 21603 18856
rect 21545 18847 21603 18853
rect 22186 18844 22192 18856
rect 22244 18844 22250 18896
rect 22278 18844 22284 18896
rect 22336 18884 22342 18896
rect 23106 18884 23112 18896
rect 22336 18856 23112 18884
rect 22336 18844 22342 18856
rect 23106 18844 23112 18856
rect 23164 18844 23170 18896
rect 2958 18816 2964 18828
rect 2919 18788 2964 18816
rect 2958 18776 2964 18788
rect 3016 18776 3022 18828
rect 4890 18816 4896 18828
rect 4851 18788 4896 18816
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 4982 18776 4988 18828
rect 5040 18816 5046 18828
rect 5258 18816 5264 18828
rect 5040 18788 5264 18816
rect 5040 18776 5046 18788
rect 5258 18776 5264 18788
rect 5316 18776 5322 18828
rect 5350 18776 5356 18828
rect 5408 18816 5414 18828
rect 7285 18819 7343 18825
rect 7285 18816 7297 18819
rect 5408 18788 7297 18816
rect 5408 18776 5414 18788
rect 7285 18785 7297 18788
rect 7331 18816 7343 18819
rect 8018 18816 8024 18828
rect 7331 18788 8024 18816
rect 7331 18785 7343 18788
rect 7285 18779 7343 18785
rect 8018 18776 8024 18788
rect 8076 18776 8082 18828
rect 8110 18776 8116 18828
rect 8168 18816 8174 18828
rect 10778 18816 10784 18828
rect 8168 18788 8213 18816
rect 10739 18788 10784 18816
rect 8168 18776 8174 18788
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 11057 18819 11115 18825
rect 11057 18785 11069 18819
rect 11103 18816 11115 18819
rect 11330 18816 11336 18828
rect 11103 18788 11336 18816
rect 11103 18785 11115 18788
rect 11057 18779 11115 18785
rect 5537 18751 5595 18757
rect 5537 18717 5549 18751
rect 5583 18748 5595 18751
rect 6181 18751 6239 18757
rect 6181 18748 6193 18751
rect 5583 18720 6193 18748
rect 5583 18717 5595 18720
rect 5537 18711 5595 18717
rect 6181 18717 6193 18720
rect 6227 18748 6239 18751
rect 6365 18751 6423 18757
rect 6365 18748 6377 18751
rect 6227 18720 6377 18748
rect 6227 18717 6239 18720
rect 6181 18711 6239 18717
rect 6365 18717 6377 18720
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 11072 18748 11100 18779
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 14252 18819 14310 18825
rect 14252 18785 14264 18819
rect 14298 18816 14310 18819
rect 14366 18816 14372 18828
rect 14298 18788 14372 18816
rect 14298 18785 14310 18788
rect 14252 18779 14310 18785
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 17678 18816 17684 18828
rect 17639 18788 17684 18816
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 18012 18788 18153 18816
rect 18012 18776 18018 18788
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 10459 18720 11100 18748
rect 12069 18751 12127 18757
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12526 18748 12532 18760
rect 12115 18720 12532 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18717 15899 18751
rect 19334 18748 19340 18760
rect 19295 18720 19340 18748
rect 15841 18711 15899 18717
rect 14323 18683 14381 18689
rect 14323 18649 14335 18683
rect 14369 18680 14381 18683
rect 15013 18683 15071 18689
rect 15013 18680 15025 18683
rect 14369 18652 15025 18680
rect 14369 18649 14381 18652
rect 14323 18643 14381 18649
rect 15013 18649 15025 18652
rect 15059 18680 15071 18683
rect 15856 18680 15884 18711
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 21450 18748 21456 18760
rect 20772 18720 21456 18748
rect 20772 18708 20778 18720
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 22646 18708 22652 18760
rect 22704 18748 22710 18760
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 22704 18720 23029 18748
rect 22704 18708 22710 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 23293 18751 23351 18757
rect 23293 18717 23305 18751
rect 23339 18717 23351 18751
rect 23293 18711 23351 18717
rect 15059 18652 15884 18680
rect 15059 18649 15071 18652
rect 15013 18643 15071 18649
rect 20806 18640 20812 18692
rect 20864 18680 20870 18692
rect 22002 18680 22008 18692
rect 20864 18652 21357 18680
rect 21963 18652 22008 18680
rect 20864 18640 20870 18652
rect 1762 18572 1768 18624
rect 1820 18612 1826 18624
rect 2222 18612 2228 18624
rect 1820 18584 2228 18612
rect 1820 18572 1826 18584
rect 2222 18572 2228 18584
rect 2280 18572 2286 18624
rect 2682 18612 2688 18624
rect 2643 18584 2688 18612
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 3694 18612 3700 18624
rect 3655 18584 3700 18612
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 7374 18572 7380 18624
rect 7432 18612 7438 18624
rect 8251 18615 8309 18621
rect 8251 18612 8263 18615
rect 7432 18584 8263 18612
rect 7432 18572 7438 18584
rect 8251 18581 8263 18584
rect 8297 18581 8309 18615
rect 8251 18575 8309 18581
rect 15286 18572 15292 18624
rect 15344 18612 15350 18624
rect 15565 18615 15623 18621
rect 15565 18612 15577 18615
rect 15344 18584 15577 18612
rect 15344 18572 15350 18584
rect 15565 18581 15577 18584
rect 15611 18612 15623 18615
rect 16482 18612 16488 18624
rect 15611 18584 16488 18612
rect 15611 18581 15623 18584
rect 15565 18575 15623 18581
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 21174 18612 21180 18624
rect 21135 18584 21180 18612
rect 21174 18572 21180 18584
rect 21232 18572 21238 18624
rect 21329 18612 21357 18652
rect 22002 18640 22008 18652
rect 22060 18640 22066 18692
rect 23308 18612 23336 18711
rect 21329 18584 23336 18612
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 3970 18408 3976 18420
rect 2832 18380 3976 18408
rect 2832 18368 2838 18380
rect 3970 18368 3976 18380
rect 4028 18408 4034 18420
rect 8389 18411 8447 18417
rect 8389 18408 8401 18411
rect 4028 18380 8401 18408
rect 4028 18368 4034 18380
rect 8389 18377 8401 18380
rect 8435 18377 8447 18411
rect 8389 18371 8447 18377
rect 8619 18411 8677 18417
rect 8619 18377 8631 18411
rect 8665 18408 8677 18411
rect 8938 18408 8944 18420
rect 8665 18380 8944 18408
rect 8665 18377 8677 18380
rect 8619 18371 8677 18377
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 11471 18411 11529 18417
rect 11471 18408 11483 18411
rect 10192 18380 11483 18408
rect 10192 18368 10198 18380
rect 11471 18377 11483 18380
rect 11517 18377 11529 18411
rect 11471 18371 11529 18377
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 14093 18411 14151 18417
rect 14093 18408 14105 18411
rect 13688 18380 14105 18408
rect 13688 18368 13694 18380
rect 14093 18377 14105 18380
rect 14139 18377 14151 18411
rect 14093 18371 14151 18377
rect 14277 18411 14335 18417
rect 14277 18377 14289 18411
rect 14323 18408 14335 18411
rect 14366 18408 14372 18420
rect 14323 18380 14372 18408
rect 14323 18377 14335 18380
rect 14277 18371 14335 18377
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 15930 18408 15936 18420
rect 15891 18380 15936 18408
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16301 18411 16359 18417
rect 16301 18377 16313 18411
rect 16347 18408 16359 18411
rect 16850 18408 16856 18420
rect 16347 18380 16856 18408
rect 16347 18377 16359 18380
rect 16301 18371 16359 18377
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 17494 18368 17500 18420
rect 17552 18408 17558 18420
rect 18187 18411 18245 18417
rect 18187 18408 18199 18411
rect 17552 18380 18199 18408
rect 17552 18368 17558 18380
rect 18187 18377 18199 18380
rect 18233 18377 18245 18411
rect 18187 18371 18245 18377
rect 18690 18368 18696 18420
rect 18748 18408 18754 18420
rect 19058 18408 19064 18420
rect 18748 18380 19064 18408
rect 18748 18368 18754 18380
rect 19058 18368 19064 18380
rect 19116 18368 19122 18420
rect 21266 18368 21272 18420
rect 21324 18408 21330 18420
rect 21913 18411 21971 18417
rect 21913 18408 21925 18411
rect 21324 18380 21925 18408
rect 21324 18368 21330 18380
rect 21913 18377 21925 18380
rect 21959 18377 21971 18411
rect 21913 18371 21971 18377
rect 23017 18411 23075 18417
rect 23017 18377 23029 18411
rect 23063 18408 23075 18411
rect 23106 18408 23112 18420
rect 23063 18380 23112 18408
rect 23063 18377 23075 18380
rect 23017 18371 23075 18377
rect 23106 18368 23112 18380
rect 23164 18368 23170 18420
rect 3142 18300 3148 18352
rect 3200 18340 3206 18352
rect 4065 18343 4123 18349
rect 4065 18340 4077 18343
rect 3200 18312 4077 18340
rect 3200 18300 3206 18312
rect 4065 18309 4077 18312
rect 4111 18340 4123 18343
rect 4430 18340 4436 18352
rect 4111 18312 4436 18340
rect 4111 18309 4123 18312
rect 4065 18303 4123 18309
rect 4430 18300 4436 18312
rect 4488 18300 4494 18352
rect 11149 18343 11207 18349
rect 5184 18312 7972 18340
rect 3418 18272 3424 18284
rect 3379 18244 3424 18272
rect 3418 18232 3424 18244
rect 3476 18232 3482 18284
rect 3510 18232 3516 18284
rect 3568 18272 3574 18284
rect 5184 18272 5212 18312
rect 3568 18244 5212 18272
rect 5261 18275 5319 18281
rect 3568 18232 3574 18244
rect 5261 18241 5273 18275
rect 5307 18272 5319 18275
rect 5534 18272 5540 18284
rect 5307 18244 5540 18272
rect 5307 18241 5319 18244
rect 5261 18235 5319 18241
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 5905 18275 5963 18281
rect 5905 18241 5917 18275
rect 5951 18272 5963 18275
rect 7009 18275 7067 18281
rect 7009 18272 7021 18275
rect 5951 18244 7021 18272
rect 5951 18241 5963 18244
rect 5905 18235 5963 18241
rect 7009 18241 7021 18244
rect 7055 18272 7067 18275
rect 7834 18272 7840 18284
rect 7055 18244 7840 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 3142 18136 3148 18148
rect 3103 18108 3148 18136
rect 3142 18096 3148 18108
rect 3200 18096 3206 18148
rect 3237 18139 3295 18145
rect 3237 18105 3249 18139
rect 3283 18136 3295 18139
rect 3786 18136 3792 18148
rect 3283 18108 3792 18136
rect 3283 18105 3295 18108
rect 3237 18099 3295 18105
rect 2038 18068 2044 18080
rect 1999 18040 2044 18068
rect 2038 18028 2044 18040
rect 2096 18028 2102 18080
rect 2593 18071 2651 18077
rect 2593 18037 2605 18071
rect 2639 18068 2651 18071
rect 2958 18068 2964 18080
rect 2639 18040 2964 18068
rect 2639 18037 2651 18040
rect 2593 18031 2651 18037
rect 2958 18028 2964 18040
rect 3016 18068 3022 18080
rect 3252 18068 3280 18099
rect 3786 18096 3792 18108
rect 3844 18096 3850 18148
rect 4525 18139 4583 18145
rect 4525 18105 4537 18139
rect 4571 18136 4583 18139
rect 4982 18136 4988 18148
rect 4571 18108 4988 18136
rect 4571 18105 4583 18108
rect 4525 18099 4583 18105
rect 4982 18096 4988 18108
rect 5040 18096 5046 18148
rect 5350 18136 5356 18148
rect 5311 18108 5356 18136
rect 5350 18096 5356 18108
rect 5408 18096 5414 18148
rect 7098 18096 7104 18148
rect 7156 18136 7162 18148
rect 7653 18139 7711 18145
rect 7156 18108 7201 18136
rect 7156 18096 7162 18108
rect 7653 18105 7665 18139
rect 7699 18136 7711 18139
rect 7944 18136 7972 18312
rect 11149 18309 11161 18343
rect 11195 18340 11207 18343
rect 11330 18340 11336 18352
rect 11195 18312 11336 18340
rect 11195 18309 11207 18312
rect 11149 18303 11207 18309
rect 11330 18300 11336 18312
rect 11388 18300 11394 18352
rect 13262 18300 13268 18352
rect 13320 18340 13326 18352
rect 13722 18340 13728 18352
rect 13320 18312 13728 18340
rect 13320 18300 13326 18312
rect 13722 18300 13728 18312
rect 13780 18340 13786 18352
rect 16390 18340 16396 18352
rect 13780 18312 16396 18340
rect 13780 18300 13786 18312
rect 16390 18300 16396 18312
rect 16448 18300 16454 18352
rect 20530 18340 20536 18352
rect 20443 18312 20536 18340
rect 20530 18300 20536 18312
rect 20588 18340 20594 18352
rect 22278 18340 22284 18352
rect 20588 18312 22284 18340
rect 20588 18300 20594 18312
rect 22278 18300 22284 18312
rect 22336 18300 22342 18352
rect 9769 18275 9827 18281
rect 9769 18241 9781 18275
rect 9815 18272 9827 18275
rect 9950 18272 9956 18284
rect 9815 18244 9956 18272
rect 9815 18241 9827 18244
rect 9769 18235 9827 18241
rect 9950 18232 9956 18244
rect 10008 18232 10014 18284
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 13817 18275 13875 18281
rect 13817 18272 13829 18275
rect 12584 18244 13829 18272
rect 12584 18232 12590 18244
rect 13817 18241 13829 18244
rect 13863 18241 13875 18275
rect 13817 18235 13875 18241
rect 14093 18275 14151 18281
rect 14093 18241 14105 18275
rect 14139 18272 14151 18275
rect 16408 18272 16436 18300
rect 14139 18244 16344 18272
rect 16408 18244 16896 18272
rect 14139 18241 14151 18244
rect 14093 18235 14151 18241
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18204 8447 18207
rect 8941 18207 8999 18213
rect 8941 18204 8953 18207
rect 8435 18176 8953 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 8941 18173 8953 18176
rect 8987 18173 8999 18207
rect 8941 18167 8999 18173
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18204 10471 18207
rect 10686 18204 10692 18216
rect 10459 18176 10692 18204
rect 10459 18173 10471 18176
rect 10413 18167 10471 18173
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 11400 18207 11458 18213
rect 11400 18173 11412 18207
rect 11446 18204 11458 18207
rect 11698 18204 11704 18216
rect 11446 18176 11704 18204
rect 11446 18173 11458 18176
rect 11400 18167 11458 18173
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12124 18176 12449 18204
rect 12124 18164 12130 18176
rect 12437 18173 12449 18176
rect 12483 18204 12495 18207
rect 12710 18204 12716 18216
rect 12483 18176 12716 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18204 13047 18207
rect 13035 18176 13308 18204
rect 13035 18173 13047 18176
rect 12989 18167 13047 18173
rect 8846 18136 8852 18148
rect 7699 18108 8852 18136
rect 7699 18105 7711 18108
rect 7653 18099 7711 18105
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 9582 18136 9588 18148
rect 9495 18108 9588 18136
rect 9582 18096 9588 18108
rect 9640 18136 9646 18148
rect 9861 18139 9919 18145
rect 9861 18136 9873 18139
rect 9640 18108 9873 18136
rect 9640 18096 9646 18108
rect 9861 18105 9873 18108
rect 9907 18105 9919 18139
rect 10778 18136 10784 18148
rect 10691 18108 10784 18136
rect 9861 18099 9919 18105
rect 10778 18096 10784 18108
rect 10836 18136 10842 18148
rect 13170 18136 13176 18148
rect 10836 18108 13176 18136
rect 10836 18096 10842 18108
rect 13170 18096 13176 18108
rect 13228 18096 13234 18148
rect 13280 18080 13308 18176
rect 14918 18136 14924 18148
rect 14879 18108 14924 18136
rect 14918 18096 14924 18108
rect 14976 18096 14982 18148
rect 15013 18139 15071 18145
rect 15013 18105 15025 18139
rect 15059 18105 15071 18139
rect 15013 18099 15071 18105
rect 4890 18068 4896 18080
rect 3016 18040 3280 18068
rect 4803 18040 4896 18068
rect 3016 18028 3022 18040
rect 4890 18028 4896 18040
rect 4948 18068 4954 18080
rect 6270 18068 6276 18080
rect 4948 18040 6276 18068
rect 4948 18028 4954 18040
rect 6270 18028 6276 18040
rect 6328 18028 6334 18080
rect 6454 18068 6460 18080
rect 6415 18040 6460 18068
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 7742 18028 7748 18080
rect 7800 18068 7806 18080
rect 8110 18068 8116 18080
rect 7800 18040 8116 18068
rect 7800 18028 7806 18040
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 12158 18068 12164 18080
rect 12119 18040 12164 18068
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 12526 18068 12532 18080
rect 12487 18040 12532 18068
rect 12526 18028 12532 18040
rect 12584 18028 12590 18080
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 13320 18040 13461 18068
rect 13320 18028 13326 18040
rect 13449 18037 13461 18040
rect 13495 18037 13507 18071
rect 13449 18031 13507 18037
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 14366 18068 14372 18080
rect 13596 18040 14372 18068
rect 13596 18028 13602 18040
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 14642 18068 14648 18080
rect 14603 18040 14648 18068
rect 14642 18028 14648 18040
rect 14700 18068 14706 18080
rect 15028 18068 15056 18099
rect 15378 18096 15384 18148
rect 15436 18136 15442 18148
rect 15565 18139 15623 18145
rect 15565 18136 15577 18139
rect 15436 18108 15577 18136
rect 15436 18096 15442 18108
rect 15565 18105 15577 18108
rect 15611 18136 15623 18139
rect 15654 18136 15660 18148
rect 15611 18108 15660 18136
rect 15611 18105 15623 18108
rect 15565 18099 15623 18105
rect 15654 18096 15660 18108
rect 15712 18096 15718 18148
rect 16316 18136 16344 18244
rect 16669 18207 16727 18213
rect 16669 18173 16681 18207
rect 16715 18204 16727 18207
rect 16758 18204 16764 18216
rect 16715 18176 16764 18204
rect 16715 18173 16727 18176
rect 16669 18167 16727 18173
rect 16758 18164 16764 18176
rect 16816 18164 16822 18216
rect 16868 18213 16896 18244
rect 17770 18232 17776 18284
rect 17828 18272 17834 18284
rect 17828 18244 23060 18272
rect 17828 18232 17834 18244
rect 16853 18207 16911 18213
rect 16853 18173 16865 18207
rect 16899 18173 16911 18207
rect 16853 18167 16911 18173
rect 18116 18207 18174 18213
rect 18116 18173 18128 18207
rect 18162 18204 18174 18207
rect 19242 18204 19248 18216
rect 18162 18176 18644 18204
rect 19203 18176 19248 18204
rect 18162 18173 18174 18176
rect 18116 18167 18174 18173
rect 17678 18136 17684 18148
rect 16316 18108 17684 18136
rect 17678 18096 17684 18108
rect 17736 18096 17742 18148
rect 16482 18068 16488 18080
rect 14700 18040 15056 18068
rect 16443 18040 16488 18068
rect 14700 18028 14706 18040
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 18616 18077 18644 18176
rect 19242 18164 19248 18176
rect 19300 18164 19306 18216
rect 20993 18207 21051 18213
rect 20993 18173 21005 18207
rect 21039 18204 21051 18207
rect 21174 18204 21180 18216
rect 21039 18176 21180 18204
rect 21039 18173 21051 18176
rect 20993 18167 21051 18173
rect 21174 18164 21180 18176
rect 21232 18204 21238 18216
rect 22554 18204 22560 18216
rect 21232 18176 22560 18204
rect 21232 18164 21238 18176
rect 22554 18164 22560 18176
rect 22612 18164 22618 18216
rect 23032 18204 23060 18244
rect 23385 18207 23443 18213
rect 23385 18204 23397 18207
rect 23032 18176 23397 18204
rect 23385 18173 23397 18176
rect 23431 18173 23443 18207
rect 23385 18167 23443 18173
rect 23661 18207 23719 18213
rect 23661 18173 23673 18207
rect 23707 18173 23719 18207
rect 23661 18167 23719 18173
rect 19058 18096 19064 18148
rect 19116 18136 19122 18148
rect 19566 18139 19624 18145
rect 19566 18136 19578 18139
rect 19116 18108 19578 18136
rect 19116 18096 19122 18108
rect 19566 18105 19578 18108
rect 19612 18136 19624 18139
rect 20809 18139 20867 18145
rect 20809 18136 20821 18139
rect 19612 18108 20821 18136
rect 19612 18105 19624 18108
rect 19566 18099 19624 18105
rect 20809 18105 20821 18108
rect 20855 18136 20867 18139
rect 21314 18139 21372 18145
rect 21314 18136 21326 18139
rect 20855 18108 21326 18136
rect 20855 18105 20867 18108
rect 20809 18099 20867 18105
rect 21314 18105 21326 18108
rect 21360 18105 21372 18139
rect 23400 18136 23428 18167
rect 23676 18136 23704 18167
rect 24026 18164 24032 18216
rect 24084 18204 24090 18216
rect 24121 18207 24179 18213
rect 24121 18204 24133 18207
rect 24084 18176 24133 18204
rect 24084 18164 24090 18176
rect 24121 18173 24133 18176
rect 24167 18173 24179 18207
rect 24121 18167 24179 18173
rect 23400 18108 23704 18136
rect 21314 18099 21372 18105
rect 18601 18071 18659 18077
rect 18601 18037 18613 18071
rect 18647 18068 18659 18071
rect 18690 18068 18696 18080
rect 18647 18040 18696 18068
rect 18647 18037 18659 18040
rect 18601 18031 18659 18037
rect 18690 18028 18696 18040
rect 18748 18028 18754 18080
rect 20165 18071 20223 18077
rect 20165 18037 20177 18071
rect 20211 18068 20223 18071
rect 21082 18068 21088 18080
rect 20211 18040 21088 18068
rect 20211 18037 20223 18040
rect 20165 18031 20223 18037
rect 21082 18028 21088 18040
rect 21140 18028 21146 18080
rect 22186 18068 22192 18080
rect 22147 18040 22192 18068
rect 22186 18028 22192 18040
rect 22244 18028 22250 18080
rect 22646 18068 22652 18080
rect 22607 18040 22652 18068
rect 22646 18028 22652 18040
rect 22704 18028 22710 18080
rect 23750 18068 23756 18080
rect 23711 18040 23756 18068
rect 23750 18028 23756 18040
rect 23808 18028 23814 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1535 17867 1593 17873
rect 1535 17833 1547 17867
rect 1581 17864 1593 17867
rect 1946 17864 1952 17876
rect 1581 17836 1952 17864
rect 1581 17833 1593 17836
rect 1535 17827 1593 17833
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 5261 17867 5319 17873
rect 5261 17833 5273 17867
rect 5307 17864 5319 17867
rect 5350 17864 5356 17876
rect 5307 17836 5356 17864
rect 5307 17833 5319 17836
rect 5261 17827 5319 17833
rect 5350 17824 5356 17836
rect 5408 17824 5414 17876
rect 6454 17864 6460 17876
rect 6415 17836 6460 17864
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 7009 17867 7067 17873
rect 7009 17833 7021 17867
rect 7055 17864 7067 17867
rect 7098 17864 7104 17876
rect 7055 17836 7104 17864
rect 7055 17833 7067 17836
rect 7009 17827 7067 17833
rect 7098 17824 7104 17836
rect 7156 17864 7162 17876
rect 7285 17867 7343 17873
rect 7285 17864 7297 17867
rect 7156 17836 7297 17864
rect 7156 17824 7162 17836
rect 7285 17833 7297 17836
rect 7331 17833 7343 17867
rect 7285 17827 7343 17833
rect 7745 17867 7803 17873
rect 7745 17833 7757 17867
rect 7791 17864 7803 17867
rect 7834 17864 7840 17876
rect 7791 17836 7840 17864
rect 7791 17833 7803 17836
rect 7745 17827 7803 17833
rect 7834 17824 7840 17836
rect 7892 17824 7898 17876
rect 9950 17864 9956 17876
rect 9911 17836 9956 17864
rect 9950 17824 9956 17836
rect 10008 17824 10014 17876
rect 11425 17867 11483 17873
rect 11425 17833 11437 17867
rect 11471 17864 11483 17867
rect 11698 17864 11704 17876
rect 11471 17836 11704 17864
rect 11471 17833 11483 17836
rect 11425 17827 11483 17833
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 12676 17836 13001 17864
rect 12676 17824 12682 17836
rect 12989 17833 13001 17836
rect 13035 17833 13047 17867
rect 12989 17827 13047 17833
rect 14369 17867 14427 17873
rect 14369 17833 14381 17867
rect 14415 17864 14427 17867
rect 14642 17864 14648 17876
rect 14415 17836 14648 17864
rect 14415 17833 14427 17836
rect 14369 17827 14427 17833
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 14918 17864 14924 17876
rect 14879 17836 14924 17864
rect 14918 17824 14924 17836
rect 14976 17864 14982 17876
rect 16206 17864 16212 17876
rect 14976 17836 16212 17864
rect 14976 17824 14982 17836
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 16390 17864 16396 17876
rect 16351 17836 16396 17864
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 18969 17867 19027 17873
rect 18969 17833 18981 17867
rect 19015 17864 19027 17867
rect 19334 17864 19340 17876
rect 19015 17836 19340 17864
rect 19015 17833 19027 17836
rect 18969 17827 19027 17833
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 20714 17864 20720 17876
rect 20675 17836 20720 17864
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 22554 17864 22560 17876
rect 22515 17836 22560 17864
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 22646 17824 22652 17876
rect 22704 17864 22710 17876
rect 25179 17867 25237 17873
rect 25179 17864 25191 17867
rect 22704 17836 25191 17864
rect 22704 17824 22710 17836
rect 25179 17833 25191 17836
rect 25225 17833 25237 17867
rect 25179 17827 25237 17833
rect 2038 17756 2044 17808
rect 2096 17796 2102 17808
rect 2501 17799 2559 17805
rect 2501 17796 2513 17799
rect 2096 17768 2513 17796
rect 2096 17756 2102 17768
rect 2501 17765 2513 17768
rect 2547 17765 2559 17799
rect 2501 17759 2559 17765
rect 2593 17799 2651 17805
rect 2593 17765 2605 17799
rect 2639 17796 2651 17799
rect 2682 17796 2688 17808
rect 2639 17768 2688 17796
rect 2639 17765 2651 17768
rect 2593 17759 2651 17765
rect 2682 17756 2688 17768
rect 2740 17756 2746 17808
rect 3145 17799 3203 17805
rect 3145 17765 3157 17799
rect 3191 17796 3203 17799
rect 3418 17796 3424 17808
rect 3191 17768 3424 17796
rect 3191 17765 3203 17768
rect 3145 17759 3203 17765
rect 3418 17756 3424 17768
rect 3476 17756 3482 17808
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 4249 17799 4307 17805
rect 4249 17796 4261 17799
rect 4212 17768 4261 17796
rect 4212 17756 4218 17768
rect 4249 17765 4261 17768
rect 4295 17765 4307 17799
rect 8018 17796 8024 17808
rect 7979 17768 8024 17796
rect 4249 17759 4307 17765
rect 8018 17756 8024 17768
rect 8076 17756 8082 17808
rect 8573 17799 8631 17805
rect 8573 17765 8585 17799
rect 8619 17796 8631 17799
rect 8846 17796 8852 17808
rect 8619 17768 8852 17796
rect 8619 17765 8631 17768
rect 8573 17759 8631 17765
rect 8846 17756 8852 17768
rect 8904 17756 8910 17808
rect 10229 17799 10287 17805
rect 10229 17765 10241 17799
rect 10275 17796 10287 17799
rect 10594 17796 10600 17808
rect 10275 17768 10600 17796
rect 10275 17765 10287 17768
rect 10229 17759 10287 17765
rect 10594 17756 10600 17768
rect 10652 17756 10658 17808
rect 11790 17796 11796 17808
rect 11751 17768 11796 17796
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 12710 17796 12716 17808
rect 12671 17768 12716 17796
rect 12710 17756 12716 17768
rect 12768 17796 12774 17808
rect 13811 17799 13869 17805
rect 12768 17768 13768 17796
rect 12768 17756 12774 17768
rect 1464 17731 1522 17737
rect 1464 17697 1476 17731
rect 1510 17728 1522 17731
rect 2314 17728 2320 17740
rect 1510 17700 2320 17728
rect 1510 17697 1522 17700
rect 1464 17691 1522 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 7742 17728 7748 17740
rect 6012 17700 7748 17728
rect 1578 17620 1584 17672
rect 1636 17660 1642 17672
rect 1949 17663 2007 17669
rect 1949 17660 1961 17663
rect 1636 17632 1961 17660
rect 1636 17620 1642 17632
rect 1949 17629 1961 17632
rect 1995 17660 2007 17663
rect 3510 17660 3516 17672
rect 1995 17632 3516 17660
rect 1995 17629 2007 17632
rect 1949 17623 2007 17629
rect 3510 17620 3516 17632
rect 3568 17620 3574 17672
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4430 17660 4436 17672
rect 4212 17632 4257 17660
rect 4391 17632 4436 17660
rect 4212 17620 4218 17632
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 14 17552 20 17604
rect 72 17592 78 17604
rect 6012 17592 6040 17700
rect 7742 17688 7748 17700
rect 7800 17688 7806 17740
rect 12342 17688 12348 17740
rect 12400 17728 12406 17740
rect 13449 17731 13507 17737
rect 13449 17728 13461 17731
rect 12400 17700 13461 17728
rect 12400 17688 12406 17700
rect 13449 17697 13461 17700
rect 13495 17728 13507 17731
rect 13538 17728 13544 17740
rect 13495 17700 13544 17728
rect 13495 17697 13507 17700
rect 13449 17691 13507 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 13740 17728 13768 17768
rect 13811 17765 13823 17799
rect 13857 17796 13869 17799
rect 14458 17796 14464 17808
rect 13857 17768 14464 17796
rect 13857 17765 13869 17768
rect 13811 17759 13869 17765
rect 14458 17756 14464 17768
rect 14516 17756 14522 17808
rect 15470 17796 15476 17808
rect 15431 17768 15476 17796
rect 15470 17756 15476 17768
rect 15528 17756 15534 17808
rect 18230 17796 18236 17808
rect 18191 17768 18236 17796
rect 18230 17756 18236 17768
rect 18288 17756 18294 17808
rect 21082 17796 21088 17808
rect 18524 17768 19564 17796
rect 21043 17768 21088 17796
rect 17494 17728 17500 17740
rect 13740 17700 13814 17728
rect 17407 17700 17500 17728
rect 6089 17663 6147 17669
rect 6089 17629 6101 17663
rect 6135 17629 6147 17663
rect 6089 17623 6147 17629
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17660 7987 17663
rect 8294 17660 8300 17672
rect 7975 17632 8300 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 72 17564 6040 17592
rect 72 17552 78 17564
rect 2958 17484 2964 17536
rect 3016 17524 3022 17536
rect 3421 17527 3479 17533
rect 3421 17524 3433 17527
rect 3016 17496 3433 17524
rect 3016 17484 3022 17496
rect 3421 17493 3433 17496
rect 3467 17493 3479 17527
rect 5534 17524 5540 17536
rect 5495 17496 5540 17524
rect 3421 17487 3479 17493
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 5994 17524 6000 17536
rect 5955 17496 6000 17524
rect 5994 17484 6000 17496
rect 6052 17524 6058 17536
rect 6104 17524 6132 17623
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 10134 17660 10140 17672
rect 10095 17632 10140 17660
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 10704 17632 11713 17660
rect 10704 17604 10732 17632
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11974 17660 11980 17672
rect 11935 17632 11980 17660
rect 11701 17623 11759 17629
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 10686 17592 10692 17604
rect 10647 17564 10692 17592
rect 10686 17552 10692 17564
rect 10744 17552 10750 17604
rect 11330 17552 11336 17604
rect 11388 17592 11394 17604
rect 13630 17592 13636 17604
rect 11388 17564 13636 17592
rect 11388 17552 11394 17564
rect 13630 17552 13636 17564
rect 13688 17552 13694 17604
rect 13786 17592 13814 17700
rect 17494 17688 17500 17700
rect 17552 17688 17558 17740
rect 17954 17728 17960 17740
rect 17915 17700 17960 17728
rect 17954 17688 17960 17700
rect 18012 17728 18018 17740
rect 18524 17737 18552 17768
rect 19536 17740 19564 17768
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 18509 17731 18567 17737
rect 18509 17728 18521 17731
rect 18012 17700 18521 17728
rect 18012 17688 18018 17700
rect 18509 17697 18521 17700
rect 18555 17697 18567 17731
rect 18509 17691 18567 17697
rect 19061 17731 19119 17737
rect 19061 17697 19073 17731
rect 19107 17697 19119 17731
rect 19518 17728 19524 17740
rect 19431 17700 19524 17728
rect 19061 17691 19119 17697
rect 15378 17660 15384 17672
rect 15339 17632 15384 17660
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 15654 17660 15660 17672
rect 15615 17632 15660 17660
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 19076 17604 19104 17691
rect 19518 17688 19524 17700
rect 19576 17688 19582 17740
rect 22462 17728 22468 17740
rect 22423 17700 22468 17728
rect 22462 17688 22468 17700
rect 22520 17688 22526 17740
rect 22922 17728 22928 17740
rect 22883 17700 22928 17728
rect 22922 17688 22928 17700
rect 22980 17728 22986 17740
rect 23661 17731 23719 17737
rect 23661 17728 23673 17731
rect 22980 17700 23673 17728
rect 22980 17688 22986 17700
rect 23661 17697 23673 17700
rect 23707 17728 23719 17731
rect 24026 17728 24032 17740
rect 23707 17700 24032 17728
rect 23707 17697 23719 17700
rect 23661 17691 23719 17697
rect 24026 17688 24032 17700
rect 24084 17688 24090 17740
rect 25108 17731 25166 17737
rect 25108 17697 25120 17731
rect 25154 17728 25166 17731
rect 25222 17728 25228 17740
rect 25154 17700 25228 17728
rect 25154 17697 25166 17700
rect 25108 17691 25166 17697
rect 25222 17688 25228 17700
rect 25280 17688 25286 17740
rect 19610 17660 19616 17672
rect 19571 17632 19616 17660
rect 19610 17620 19616 17632
rect 19668 17620 19674 17672
rect 20806 17620 20812 17672
rect 20864 17660 20870 17672
rect 20993 17663 21051 17669
rect 20993 17660 21005 17663
rect 20864 17632 21005 17660
rect 20864 17620 20870 17632
rect 20993 17629 21005 17632
rect 21039 17629 21051 17663
rect 23750 17660 23756 17672
rect 20993 17623 21051 17629
rect 21100 17632 23756 17660
rect 17402 17592 17408 17604
rect 13786 17564 17408 17592
rect 17402 17552 17408 17564
rect 17460 17592 17466 17604
rect 19058 17592 19064 17604
rect 17460 17564 19064 17592
rect 17460 17552 17466 17564
rect 19058 17552 19064 17564
rect 19116 17552 19122 17604
rect 19242 17552 19248 17604
rect 19300 17592 19306 17604
rect 20165 17595 20223 17601
rect 20165 17592 20177 17595
rect 19300 17564 20177 17592
rect 19300 17552 19306 17564
rect 20165 17561 20177 17564
rect 20211 17592 20223 17595
rect 21100 17592 21128 17632
rect 23750 17620 23756 17632
rect 23808 17620 23814 17672
rect 23842 17620 23848 17672
rect 23900 17660 23906 17672
rect 24167 17663 24225 17669
rect 24167 17660 24179 17663
rect 23900 17632 24179 17660
rect 23900 17620 23906 17632
rect 24167 17629 24179 17632
rect 24213 17629 24225 17663
rect 24167 17623 24225 17629
rect 20211 17564 21128 17592
rect 21545 17595 21603 17601
rect 20211 17561 20223 17564
rect 20165 17555 20223 17561
rect 21545 17561 21557 17595
rect 21591 17592 21603 17595
rect 22002 17592 22008 17604
rect 21591 17564 22008 17592
rect 21591 17561 21603 17564
rect 21545 17555 21603 17561
rect 22002 17552 22008 17564
rect 22060 17592 22066 17604
rect 22060 17564 23980 17592
rect 22060 17552 22066 17564
rect 16758 17524 16764 17536
rect 6052 17496 6132 17524
rect 16719 17496 16764 17524
rect 6052 17484 6058 17496
rect 16758 17484 16764 17496
rect 16816 17484 16822 17536
rect 21910 17524 21916 17536
rect 21871 17496 21916 17524
rect 21910 17484 21916 17496
rect 21968 17484 21974 17536
rect 23952 17533 23980 17564
rect 23937 17527 23995 17533
rect 23937 17493 23949 17527
rect 23983 17524 23995 17527
rect 24026 17524 24032 17536
rect 23983 17496 24032 17524
rect 23983 17493 23995 17496
rect 23937 17487 23995 17493
rect 24026 17484 24032 17496
rect 24084 17484 24090 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2409 17323 2467 17329
rect 2409 17289 2421 17323
rect 2455 17320 2467 17323
rect 2682 17320 2688 17332
rect 2455 17292 2688 17320
rect 2455 17289 2467 17292
rect 2409 17283 2467 17289
rect 2682 17280 2688 17292
rect 2740 17280 2746 17332
rect 3786 17320 3792 17332
rect 3747 17292 3792 17320
rect 3786 17280 3792 17292
rect 3844 17280 3850 17332
rect 4062 17320 4068 17332
rect 4023 17292 4068 17320
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 7745 17323 7803 17329
rect 7745 17289 7757 17323
rect 7791 17320 7803 17323
rect 8018 17320 8024 17332
rect 7791 17292 8024 17320
rect 7791 17289 7803 17292
rect 7745 17283 7803 17289
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 10134 17280 10140 17332
rect 10192 17320 10198 17332
rect 11057 17323 11115 17329
rect 11057 17320 11069 17323
rect 10192 17292 11069 17320
rect 10192 17280 10198 17292
rect 11057 17289 11069 17292
rect 11103 17320 11115 17323
rect 14734 17320 14740 17332
rect 11103 17292 14740 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 14734 17280 14740 17292
rect 14792 17280 14798 17332
rect 15470 17320 15476 17332
rect 15431 17292 15476 17320
rect 15470 17280 15476 17292
rect 15528 17320 15534 17332
rect 15749 17323 15807 17329
rect 15749 17320 15761 17323
rect 15528 17292 15761 17320
rect 15528 17280 15534 17292
rect 15749 17289 15761 17292
rect 15795 17289 15807 17323
rect 17494 17320 17500 17332
rect 17455 17292 17500 17320
rect 15749 17283 15807 17289
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 17678 17280 17684 17332
rect 17736 17320 17742 17332
rect 17773 17323 17831 17329
rect 17773 17320 17785 17323
rect 17736 17292 17785 17320
rect 17736 17280 17742 17292
rect 17773 17289 17785 17292
rect 17819 17289 17831 17323
rect 19058 17320 19064 17332
rect 19019 17292 19064 17320
rect 17773 17283 17831 17289
rect 1535 17255 1593 17261
rect 1535 17221 1547 17255
rect 1581 17252 1593 17255
rect 10042 17252 10048 17264
rect 1581 17224 10048 17252
rect 1581 17221 1593 17224
rect 1535 17215 1593 17221
rect 10042 17212 10048 17224
rect 10100 17212 10106 17264
rect 10321 17255 10379 17261
rect 10321 17221 10333 17255
rect 10367 17252 10379 17255
rect 11790 17252 11796 17264
rect 10367 17224 11796 17252
rect 10367 17221 10379 17224
rect 10321 17215 10379 17221
rect 11790 17212 11796 17224
rect 11848 17252 11854 17264
rect 11977 17255 12035 17261
rect 11977 17252 11989 17255
rect 11848 17224 11989 17252
rect 11848 17212 11854 17224
rect 11977 17221 11989 17224
rect 12023 17221 12035 17255
rect 11977 17215 12035 17221
rect 14093 17255 14151 17261
rect 14093 17221 14105 17255
rect 14139 17252 14151 17255
rect 14458 17252 14464 17264
rect 14139 17224 14464 17252
rect 14139 17221 14151 17224
rect 14093 17215 14151 17221
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 4525 17187 4583 17193
rect 4525 17184 4537 17187
rect 4212 17156 4537 17184
rect 4212 17144 4218 17156
rect 4525 17153 4537 17156
rect 4571 17184 4583 17187
rect 11425 17187 11483 17193
rect 11425 17184 11437 17187
rect 4571 17156 11437 17184
rect 4571 17153 4583 17156
rect 4525 17147 4583 17153
rect 11425 17153 11437 17156
rect 11471 17153 11483 17187
rect 11425 17147 11483 17153
rect 12618 17144 12624 17196
rect 12676 17184 12682 17196
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 12676 17156 12817 17184
rect 12676 17144 12682 17156
rect 12805 17153 12817 17156
rect 12851 17153 12863 17187
rect 12805 17147 12863 17153
rect 1026 17076 1032 17128
rect 1084 17116 1090 17128
rect 1432 17119 1490 17125
rect 1432 17116 1444 17119
rect 1084 17088 1444 17116
rect 1084 17076 1090 17088
rect 1432 17085 1444 17088
rect 1478 17116 1490 17119
rect 1857 17119 1915 17125
rect 1857 17116 1869 17119
rect 1478 17088 1869 17116
rect 1478 17085 1490 17088
rect 1432 17079 1490 17085
rect 1857 17085 1869 17088
rect 1903 17085 1915 17119
rect 1857 17079 1915 17085
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 2958 17116 2964 17128
rect 2915 17088 2964 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 5077 17119 5135 17125
rect 5077 17116 5089 17119
rect 3384 17088 5089 17116
rect 3384 17076 3390 17088
rect 5077 17085 5089 17088
rect 5123 17116 5135 17119
rect 5445 17119 5503 17125
rect 5445 17116 5457 17119
rect 5123 17088 5457 17116
rect 5123 17085 5135 17088
rect 5077 17079 5135 17085
rect 5445 17085 5457 17088
rect 5491 17116 5503 17119
rect 5626 17116 5632 17128
rect 5491 17088 5632 17116
rect 5491 17085 5503 17088
rect 5445 17079 5503 17085
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 5721 17119 5779 17125
rect 5721 17085 5733 17119
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 6822 17116 6828 17128
rect 5951 17088 6828 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 3190 17051 3248 17057
rect 3190 17048 3202 17051
rect 2792 17020 3202 17048
rect 2792 16992 2820 17020
rect 3190 17017 3202 17020
rect 3236 17048 3248 17051
rect 5736 17048 5764 17079
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 9398 17116 9404 17128
rect 9359 17088 9404 17116
rect 9398 17076 9404 17088
rect 9456 17076 9462 17128
rect 10594 17116 10600 17128
rect 10555 17088 10600 17116
rect 10594 17076 10600 17088
rect 10652 17116 10658 17128
rect 10778 17116 10784 17128
rect 10652 17088 10784 17116
rect 10652 17076 10658 17088
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 11238 17125 11244 17128
rect 11216 17119 11244 17125
rect 11216 17116 11228 17119
rect 11151 17088 11228 17116
rect 11216 17085 11228 17088
rect 11296 17116 11302 17128
rect 11609 17119 11667 17125
rect 11609 17116 11621 17119
rect 11296 17088 11621 17116
rect 11216 17079 11244 17085
rect 11238 17076 11244 17079
rect 11296 17076 11302 17088
rect 11609 17085 11621 17088
rect 11655 17085 11667 17119
rect 11609 17079 11667 17085
rect 6086 17048 6092 17060
rect 3236 17020 5672 17048
rect 5736 17020 6092 17048
rect 3236 17017 3248 17020
rect 3190 17011 3248 17017
rect 2774 16980 2780 16992
rect 2735 16952 2780 16980
rect 2774 16940 2780 16952
rect 2832 16940 2838 16992
rect 5644 16980 5672 17020
rect 6086 17008 6092 17020
rect 6144 17008 6150 17060
rect 7146 17051 7204 17057
rect 7146 17048 7158 17051
rect 6564 17020 7158 17048
rect 6181 16983 6239 16989
rect 6181 16980 6193 16983
rect 5644 16952 6193 16980
rect 6181 16949 6193 16952
rect 6227 16980 6239 16983
rect 6454 16980 6460 16992
rect 6227 16952 6460 16980
rect 6227 16949 6239 16952
rect 6181 16943 6239 16949
rect 6454 16940 6460 16952
rect 6512 16980 6518 16992
rect 6564 16989 6592 17020
rect 7146 17017 7158 17020
rect 7192 17048 7204 17051
rect 9217 17051 9275 17057
rect 9217 17048 9229 17051
rect 7192 17020 9229 17048
rect 7192 17017 7204 17020
rect 7146 17011 7204 17017
rect 9217 17017 9229 17020
rect 9263 17048 9275 17051
rect 9763 17051 9821 17057
rect 9763 17048 9775 17051
rect 9263 17020 9775 17048
rect 9263 17017 9275 17020
rect 9217 17011 9275 17017
rect 9763 17017 9775 17020
rect 9809 17048 9821 17051
rect 10134 17048 10140 17060
rect 9809 17020 10140 17048
rect 9809 17017 9821 17020
rect 9763 17011 9821 17017
rect 10134 17008 10140 17020
rect 10192 17008 10198 17060
rect 12158 17008 12164 17060
rect 12216 17048 12222 17060
rect 12713 17051 12771 17057
rect 12713 17048 12725 17051
rect 12216 17020 12725 17048
rect 12216 17008 12222 17020
rect 12713 17017 12725 17020
rect 12759 17048 12771 17051
rect 13167 17051 13225 17057
rect 13167 17048 13179 17051
rect 12759 17020 13179 17048
rect 12759 17017 12771 17020
rect 12713 17011 12771 17017
rect 13167 17017 13179 17020
rect 13213 17048 13225 17051
rect 13630 17048 13636 17060
rect 13213 17020 13636 17048
rect 13213 17017 13225 17020
rect 13167 17011 13225 17017
rect 13630 17008 13636 17020
rect 13688 17048 13694 17060
rect 14108 17048 14136 17215
rect 14458 17212 14464 17224
rect 14516 17212 14522 17264
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 14553 17187 14611 17193
rect 14553 17184 14565 17187
rect 14332 17156 14565 17184
rect 14332 17144 14338 17156
rect 14553 17153 14565 17156
rect 14599 17153 14611 17187
rect 14553 17147 14611 17153
rect 16393 17187 16451 17193
rect 16393 17153 16405 17187
rect 16439 17184 16451 17187
rect 16758 17184 16764 17196
rect 16439 17156 16764 17184
rect 16439 17153 16451 17156
rect 16393 17147 16451 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 17788 17116 17816 17283
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19518 17280 19524 17332
rect 19576 17320 19582 17332
rect 22833 17323 22891 17329
rect 22833 17320 22845 17323
rect 19576 17292 22845 17320
rect 19576 17280 19582 17292
rect 22833 17289 22845 17292
rect 22879 17320 22891 17323
rect 22922 17320 22928 17332
rect 22879 17292 22928 17320
rect 22879 17289 22891 17292
rect 22833 17283 22891 17289
rect 22922 17280 22928 17292
rect 22980 17280 22986 17332
rect 24026 17320 24032 17332
rect 23987 17292 24032 17320
rect 24026 17280 24032 17292
rect 24084 17280 24090 17332
rect 25501 17323 25559 17329
rect 25501 17289 25513 17323
rect 25547 17320 25559 17323
rect 26234 17320 26240 17332
rect 25547 17292 26240 17320
rect 25547 17289 25559 17292
rect 25501 17283 25559 17289
rect 20533 17255 20591 17261
rect 20533 17221 20545 17255
rect 20579 17252 20591 17255
rect 22186 17252 22192 17264
rect 20579 17224 22192 17252
rect 20579 17221 20591 17224
rect 20533 17215 20591 17221
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 19610 17184 19616 17196
rect 19571 17156 19616 17184
rect 19610 17144 19616 17156
rect 19668 17184 19674 17196
rect 20254 17184 20260 17196
rect 19668 17156 20260 17184
rect 19668 17144 19674 17156
rect 20254 17144 20260 17156
rect 20312 17144 20318 17196
rect 20438 17144 20444 17196
rect 20496 17184 20502 17196
rect 20990 17184 20996 17196
rect 20496 17156 20996 17184
rect 20496 17144 20502 17156
rect 20990 17144 20996 17156
rect 21048 17184 21054 17196
rect 21729 17187 21787 17193
rect 21729 17184 21741 17187
rect 21048 17156 21741 17184
rect 21048 17144 21054 17156
rect 21729 17153 21741 17156
rect 21775 17153 21787 17187
rect 21729 17147 21787 17153
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17788 17088 18061 17116
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 18230 17076 18236 17128
rect 18288 17116 18294 17128
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 18288 17088 18521 17116
rect 18288 17076 18294 17088
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 22462 17116 22468 17128
rect 22423 17088 22468 17116
rect 18509 17079 18567 17085
rect 22462 17076 22468 17088
rect 22520 17076 22526 17128
rect 24648 17119 24706 17125
rect 24648 17085 24660 17119
rect 24694 17116 24706 17119
rect 25516 17116 25544 17283
rect 26234 17280 26240 17292
rect 26292 17280 26298 17332
rect 24694 17088 25544 17116
rect 24694 17085 24706 17088
rect 24648 17079 24706 17085
rect 14874 17051 14932 17057
rect 14874 17048 14886 17051
rect 13688 17020 14886 17048
rect 13688 17008 13694 17020
rect 14874 17017 14886 17020
rect 14920 17017 14932 17051
rect 16462 17051 16520 17057
rect 16462 17048 16474 17051
rect 14874 17011 14932 17017
rect 16316 17020 16474 17048
rect 16316 16992 16344 17020
rect 16462 17017 16474 17020
rect 16508 17017 16520 17051
rect 16462 17011 16520 17017
rect 16574 17008 16580 17060
rect 16632 17048 16638 17060
rect 17037 17051 17095 17057
rect 17037 17048 17049 17051
rect 16632 17020 17049 17048
rect 16632 17008 16638 17020
rect 17037 17017 17049 17020
rect 17083 17017 17095 17051
rect 18782 17048 18788 17060
rect 18743 17020 18788 17048
rect 17037 17011 17095 17017
rect 18782 17008 18788 17020
rect 18840 17008 18846 17060
rect 19934 17051 19992 17057
rect 19934 17048 19946 17051
rect 19444 17020 19946 17048
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6512 16952 6561 16980
rect 6512 16940 6518 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 6549 16943 6607 16949
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 8389 16983 8447 16989
rect 8389 16980 8401 16983
rect 8352 16952 8401 16980
rect 8352 16940 8358 16952
rect 8389 16949 8401 16952
rect 8435 16949 8447 16983
rect 8389 16943 8447 16949
rect 13725 16983 13783 16989
rect 13725 16949 13737 16983
rect 13771 16980 13783 16983
rect 13814 16980 13820 16992
rect 13771 16952 13820 16980
rect 13771 16949 13783 16952
rect 13725 16943 13783 16949
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 16209 16983 16267 16989
rect 16209 16949 16221 16983
rect 16255 16980 16267 16983
rect 16298 16980 16304 16992
rect 16255 16952 16304 16980
rect 16255 16949 16267 16952
rect 16209 16943 16267 16949
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 18874 16940 18880 16992
rect 18932 16980 18938 16992
rect 19444 16989 19472 17020
rect 19934 17017 19946 17020
rect 19980 17017 19992 17051
rect 19934 17011 19992 17017
rect 20993 17051 21051 17057
rect 20993 17017 21005 17051
rect 21039 17048 21051 17051
rect 21082 17048 21088 17060
rect 21039 17020 21088 17048
rect 21039 17017 21051 17020
rect 20993 17011 21051 17017
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 21453 17051 21511 17057
rect 21453 17017 21465 17051
rect 21499 17017 21511 17051
rect 21453 17011 21511 17017
rect 21545 17051 21603 17057
rect 21545 17017 21557 17051
rect 21591 17048 21603 17051
rect 21910 17048 21916 17060
rect 21591 17020 21916 17048
rect 21591 17017 21603 17020
rect 21545 17011 21603 17017
rect 19429 16983 19487 16989
rect 19429 16980 19441 16983
rect 18932 16952 19441 16980
rect 18932 16940 18938 16952
rect 19429 16949 19441 16952
rect 19475 16949 19487 16983
rect 19429 16943 19487 16949
rect 20714 16940 20720 16992
rect 20772 16980 20778 16992
rect 21468 16980 21496 17011
rect 21910 17008 21916 17020
rect 21968 17008 21974 17060
rect 21634 16980 21640 16992
rect 20772 16952 21640 16980
rect 20772 16940 20778 16952
rect 21634 16940 21640 16952
rect 21692 16940 21698 16992
rect 24026 16940 24032 16992
rect 24084 16980 24090 16992
rect 24719 16983 24777 16989
rect 24719 16980 24731 16983
rect 24084 16952 24731 16980
rect 24084 16940 24090 16952
rect 24719 16949 24731 16952
rect 24765 16949 24777 16983
rect 24719 16943 24777 16949
rect 25133 16983 25191 16989
rect 25133 16949 25145 16983
rect 25179 16980 25191 16983
rect 25222 16980 25228 16992
rect 25179 16952 25228 16980
rect 25179 16949 25191 16952
rect 25133 16943 25191 16949
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2038 16736 2044 16788
rect 2096 16776 2102 16788
rect 2225 16779 2283 16785
rect 2225 16776 2237 16779
rect 2096 16748 2237 16776
rect 2096 16736 2102 16748
rect 2225 16745 2237 16748
rect 2271 16745 2283 16779
rect 2225 16739 2283 16745
rect 5626 16736 5632 16788
rect 5684 16736 5690 16788
rect 5905 16779 5963 16785
rect 5905 16745 5917 16779
rect 5951 16776 5963 16779
rect 5994 16776 6000 16788
rect 5951 16748 6000 16776
rect 5951 16745 5963 16748
rect 5905 16739 5963 16745
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 6822 16776 6828 16788
rect 6783 16748 6828 16776
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 10597 16779 10655 16785
rect 10597 16745 10609 16779
rect 10643 16776 10655 16779
rect 10778 16776 10784 16788
rect 10643 16748 10784 16776
rect 10643 16745 10655 16748
rect 10597 16739 10655 16745
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 14645 16779 14703 16785
rect 14645 16776 14657 16779
rect 14332 16748 14657 16776
rect 14332 16736 14338 16748
rect 14645 16745 14657 16748
rect 14691 16745 14703 16779
rect 17954 16776 17960 16788
rect 14645 16739 14703 16745
rect 16960 16748 17960 16776
rect 1670 16668 1676 16720
rect 1728 16708 1734 16720
rect 2593 16711 2651 16717
rect 2593 16708 2605 16711
rect 1728 16680 2605 16708
rect 1728 16668 1734 16680
rect 2593 16677 2605 16680
rect 2639 16708 2651 16711
rect 2866 16708 2872 16720
rect 2639 16680 2872 16708
rect 2639 16677 2651 16680
rect 2593 16671 2651 16677
rect 2866 16668 2872 16680
rect 2924 16668 2930 16720
rect 3142 16708 3148 16720
rect 3103 16680 3148 16708
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 4062 16708 4068 16720
rect 4023 16680 4068 16708
rect 4062 16668 4068 16680
rect 4120 16668 4126 16720
rect 5644 16708 5672 16736
rect 8386 16708 8392 16720
rect 5644 16680 8392 16708
rect 1464 16643 1522 16649
rect 1464 16609 1476 16643
rect 1510 16640 1522 16643
rect 1578 16640 1584 16652
rect 1510 16612 1584 16640
rect 1510 16609 1522 16612
rect 1464 16603 1522 16609
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4212 16612 4257 16640
rect 4212 16600 4218 16612
rect 4338 16600 4344 16652
rect 4396 16640 4402 16652
rect 5629 16643 5687 16649
rect 5629 16640 5641 16643
rect 4396 16612 5641 16640
rect 4396 16600 4402 16612
rect 5629 16609 5641 16612
rect 5675 16640 5687 16643
rect 5902 16640 5908 16652
rect 5675 16612 5908 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 6086 16640 6092 16652
rect 6047 16612 6092 16640
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 8312 16649 8340 16680
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 8757 16711 8815 16717
rect 8757 16677 8769 16711
rect 8803 16708 8815 16711
rect 9398 16708 9404 16720
rect 8803 16680 9404 16708
rect 8803 16677 8815 16680
rect 8757 16671 8815 16677
rect 9398 16668 9404 16680
rect 9456 16668 9462 16720
rect 10039 16711 10097 16717
rect 10039 16677 10051 16711
rect 10085 16708 10097 16711
rect 10134 16708 10140 16720
rect 10085 16680 10140 16708
rect 10085 16677 10097 16680
rect 10039 16671 10097 16677
rect 10134 16668 10140 16680
rect 10192 16668 10198 16720
rect 13538 16708 13544 16720
rect 13499 16680 13544 16708
rect 13538 16668 13544 16680
rect 13596 16668 13602 16720
rect 13814 16668 13820 16720
rect 13872 16708 13878 16720
rect 14369 16711 14427 16717
rect 13872 16680 13917 16708
rect 13872 16668 13878 16680
rect 14369 16677 14381 16711
rect 14415 16708 14427 16711
rect 15470 16708 15476 16720
rect 14415 16680 15476 16708
rect 14415 16677 14427 16680
rect 14369 16671 14427 16677
rect 15470 16668 15476 16680
rect 15528 16668 15534 16720
rect 15651 16711 15709 16717
rect 15651 16677 15663 16711
rect 15697 16708 15709 16711
rect 16114 16708 16120 16720
rect 15697 16680 16120 16708
rect 15697 16677 15709 16680
rect 15651 16671 15709 16677
rect 16114 16668 16120 16680
rect 16172 16668 16178 16720
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16609 8355 16643
rect 8478 16640 8484 16652
rect 8439 16612 8484 16640
rect 8297 16603 8355 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16609 12127 16643
rect 12342 16640 12348 16652
rect 12303 16612 12348 16640
rect 12069 16603 12127 16609
rect 2498 16572 2504 16584
rect 2459 16544 2504 16572
rect 2498 16532 2504 16544
rect 2556 16532 2562 16584
rect 5442 16532 5448 16584
rect 5500 16572 5506 16584
rect 9030 16572 9036 16584
rect 5500 16544 9036 16572
rect 5500 16532 5506 16544
rect 9030 16532 9036 16544
rect 9088 16532 9094 16584
rect 9674 16572 9680 16584
rect 9635 16544 9680 16572
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 12084 16572 12112 16603
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 16960 16640 16988 16748
rect 17954 16736 17960 16748
rect 18012 16776 18018 16788
rect 18049 16779 18107 16785
rect 18049 16776 18061 16779
rect 18012 16748 18061 16776
rect 18012 16736 18018 16748
rect 18049 16745 18061 16748
rect 18095 16776 18107 16779
rect 19061 16779 19119 16785
rect 19061 16776 19073 16779
rect 18095 16748 19073 16776
rect 18095 16745 18107 16748
rect 18049 16739 18107 16745
rect 19061 16745 19073 16748
rect 19107 16745 19119 16779
rect 20254 16776 20260 16788
rect 20215 16748 20260 16776
rect 19061 16739 19119 16745
rect 20254 16736 20260 16748
rect 20312 16736 20318 16788
rect 20714 16776 20720 16788
rect 20675 16748 20720 16776
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 24075 16779 24133 16785
rect 24075 16776 24087 16779
rect 20824 16748 24087 16776
rect 17221 16711 17279 16717
rect 17221 16677 17233 16711
rect 17267 16708 17279 16711
rect 17310 16708 17316 16720
rect 17267 16680 17316 16708
rect 17267 16677 17279 16680
rect 17221 16671 17279 16677
rect 17310 16668 17316 16680
rect 17368 16668 17374 16720
rect 19426 16708 19432 16720
rect 19387 16680 19432 16708
rect 19426 16668 19432 16680
rect 19484 16668 19490 16720
rect 19981 16711 20039 16717
rect 19981 16677 19993 16711
rect 20027 16708 20039 16711
rect 20438 16708 20444 16720
rect 20027 16680 20444 16708
rect 20027 16677 20039 16680
rect 19981 16671 20039 16677
rect 20438 16668 20444 16680
rect 20496 16668 20502 16720
rect 15028 16612 16988 16640
rect 12250 16572 12256 16584
rect 12084 16544 12256 16572
rect 12250 16532 12256 16544
rect 12308 16532 12314 16584
rect 12805 16575 12863 16581
rect 12805 16541 12817 16575
rect 12851 16541 12863 16575
rect 12805 16535 12863 16541
rect 13725 16575 13783 16581
rect 13725 16541 13737 16575
rect 13771 16572 13783 16575
rect 14182 16572 14188 16584
rect 13771 16544 14188 16572
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 1535 16507 1593 16513
rect 1535 16473 1547 16507
rect 1581 16504 1593 16507
rect 3878 16504 3884 16516
rect 1581 16476 3884 16504
rect 1581 16473 1593 16476
rect 1535 16467 1593 16473
rect 3878 16464 3884 16476
rect 3936 16464 3942 16516
rect 12161 16507 12219 16513
rect 12161 16473 12173 16507
rect 12207 16504 12219 16507
rect 12618 16504 12624 16516
rect 12207 16476 12624 16504
rect 12207 16473 12219 16476
rect 12161 16467 12219 16473
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 12820 16504 12848 16535
rect 14182 16532 14188 16544
rect 14240 16532 14246 16584
rect 15028 16504 15056 16612
rect 15286 16572 15292 16584
rect 15247 16544 15292 16572
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 17129 16575 17187 16581
rect 17129 16541 17141 16575
rect 17175 16572 17187 16575
rect 17770 16572 17776 16584
rect 17175 16544 17776 16572
rect 17175 16541 17187 16544
rect 17129 16535 17187 16541
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 19337 16575 19395 16581
rect 19337 16541 19349 16575
rect 19383 16572 19395 16575
rect 19978 16572 19984 16584
rect 19383 16544 19984 16572
rect 19383 16541 19395 16544
rect 19337 16535 19395 16541
rect 19978 16532 19984 16544
rect 20036 16572 20042 16584
rect 20824 16572 20852 16748
rect 24075 16745 24087 16748
rect 24121 16745 24133 16779
rect 24075 16739 24133 16745
rect 20898 16668 20904 16720
rect 20956 16708 20962 16720
rect 21085 16711 21143 16717
rect 21085 16708 21097 16711
rect 20956 16680 21097 16708
rect 20956 16668 20962 16680
rect 21085 16677 21097 16680
rect 21131 16677 21143 16711
rect 21085 16671 21143 16677
rect 21545 16711 21603 16717
rect 21545 16677 21557 16711
rect 21591 16708 21603 16711
rect 21634 16708 21640 16720
rect 21591 16680 21640 16708
rect 21591 16677 21603 16680
rect 21545 16671 21603 16677
rect 21634 16668 21640 16680
rect 21692 16668 21698 16720
rect 22925 16643 22983 16649
rect 22925 16609 22937 16643
rect 22971 16640 22983 16643
rect 23014 16640 23020 16652
rect 22971 16612 23020 16640
rect 22971 16609 22983 16612
rect 22925 16603 22983 16609
rect 23014 16600 23020 16612
rect 23072 16600 23078 16652
rect 23934 16640 23940 16652
rect 23895 16612 23940 16640
rect 23934 16600 23940 16612
rect 23992 16600 23998 16652
rect 20036 16544 20852 16572
rect 21453 16575 21511 16581
rect 20036 16532 20042 16544
rect 21453 16541 21465 16575
rect 21499 16572 21511 16575
rect 21499 16544 22416 16572
rect 21499 16541 21511 16544
rect 21453 16535 21511 16541
rect 12820 16476 15056 16504
rect 15105 16507 15163 16513
rect 15105 16473 15117 16507
rect 15151 16504 15163 16507
rect 15378 16504 15384 16516
rect 15151 16476 15384 16504
rect 15151 16473 15163 16476
rect 15105 16467 15163 16473
rect 15378 16464 15384 16476
rect 15436 16504 15442 16516
rect 16574 16504 16580 16516
rect 15436 16476 16580 16504
rect 15436 16464 15442 16476
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 17034 16464 17040 16516
rect 17092 16504 17098 16516
rect 17681 16507 17739 16513
rect 17681 16504 17693 16507
rect 17092 16476 17693 16504
rect 17092 16464 17098 16476
rect 17681 16473 17693 16476
rect 17727 16473 17739 16507
rect 17681 16467 17739 16473
rect 21542 16464 21548 16516
rect 21600 16504 21606 16516
rect 22005 16507 22063 16513
rect 22005 16504 22017 16507
rect 21600 16476 22017 16504
rect 21600 16464 21606 16476
rect 22005 16473 22017 16476
rect 22051 16473 22063 16507
rect 22005 16467 22063 16473
rect 22388 16448 22416 16544
rect 1949 16439 2007 16445
rect 1949 16405 1961 16439
rect 1995 16436 2007 16439
rect 2314 16436 2320 16448
rect 1995 16408 2320 16436
rect 1995 16405 2007 16408
rect 1949 16399 2007 16405
rect 2314 16396 2320 16408
rect 2372 16396 2378 16448
rect 2682 16396 2688 16448
rect 2740 16436 2746 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 2740 16408 3433 16436
rect 2740 16396 2746 16408
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 3421 16399 3479 16405
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 5169 16439 5227 16445
rect 5169 16436 5181 16439
rect 5040 16408 5181 16436
rect 5040 16396 5046 16408
rect 5169 16405 5181 16408
rect 5215 16436 5227 16439
rect 6086 16436 6092 16448
rect 5215 16408 6092 16436
rect 5215 16405 5227 16408
rect 5169 16399 5227 16405
rect 6086 16396 6092 16408
rect 6144 16396 6150 16448
rect 11330 16436 11336 16448
rect 11291 16408 11336 16436
rect 11330 16396 11336 16408
rect 11388 16396 11394 16448
rect 11422 16396 11428 16448
rect 11480 16436 11486 16448
rect 11609 16439 11667 16445
rect 11609 16436 11621 16439
rect 11480 16408 11621 16436
rect 11480 16396 11486 16408
rect 11609 16405 11621 16408
rect 11655 16405 11667 16439
rect 11609 16399 11667 16405
rect 16209 16439 16267 16445
rect 16209 16405 16221 16439
rect 16255 16436 16267 16439
rect 16298 16436 16304 16448
rect 16255 16408 16304 16436
rect 16255 16405 16267 16408
rect 16209 16399 16267 16405
rect 16298 16396 16304 16408
rect 16356 16436 16362 16448
rect 16485 16439 16543 16445
rect 16485 16436 16497 16439
rect 16356 16408 16497 16436
rect 16356 16396 16362 16408
rect 16485 16405 16497 16408
rect 16531 16405 16543 16439
rect 16485 16399 16543 16405
rect 18230 16396 18236 16448
rect 18288 16436 18294 16448
rect 18417 16439 18475 16445
rect 18417 16436 18429 16439
rect 18288 16408 18429 16436
rect 18288 16396 18294 16408
rect 18417 16405 18429 16408
rect 18463 16405 18475 16439
rect 18417 16399 18475 16405
rect 22370 16396 22376 16448
rect 22428 16436 22434 16448
rect 23063 16439 23121 16445
rect 23063 16436 23075 16439
rect 22428 16408 23075 16436
rect 22428 16396 22434 16408
rect 23063 16405 23075 16408
rect 23109 16405 23121 16439
rect 23063 16399 23121 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1670 16232 1676 16244
rect 1631 16204 1676 16232
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 1946 16241 1952 16244
rect 1903 16235 1952 16241
rect 1903 16232 1915 16235
rect 1859 16204 1915 16232
rect 1903 16201 1915 16204
rect 1949 16201 1952 16235
rect 1903 16195 1952 16201
rect 1946 16192 1952 16195
rect 2004 16232 2010 16244
rect 2498 16232 2504 16244
rect 2004 16204 2504 16232
rect 2004 16192 2010 16204
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 2866 16192 2872 16244
rect 2924 16232 2930 16244
rect 3697 16235 3755 16241
rect 3697 16232 3709 16235
rect 2924 16204 3709 16232
rect 2924 16192 2930 16204
rect 3697 16201 3709 16204
rect 3743 16232 3755 16235
rect 4065 16235 4123 16241
rect 4065 16232 4077 16235
rect 3743 16204 4077 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 4065 16201 4077 16204
rect 4111 16232 4123 16235
rect 4154 16232 4160 16244
rect 4111 16204 4160 16232
rect 4111 16201 4123 16204
rect 4065 16195 4123 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 5350 16232 5356 16244
rect 4755 16204 5356 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 6052 16204 6193 16232
rect 6052 16192 6058 16204
rect 6181 16201 6193 16204
rect 6227 16232 6239 16235
rect 7466 16232 7472 16244
rect 6227 16204 7472 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 7466 16192 7472 16204
rect 7524 16232 7530 16244
rect 7742 16232 7748 16244
rect 7524 16204 7748 16232
rect 7524 16192 7530 16204
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 8386 16192 8392 16244
rect 8444 16232 8450 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 8444 16204 8769 16232
rect 8444 16192 8450 16204
rect 8757 16201 8769 16204
rect 8803 16232 8815 16235
rect 10870 16232 10876 16244
rect 8803 16204 10876 16232
rect 8803 16201 8815 16204
rect 8757 16195 8815 16201
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 12161 16235 12219 16241
rect 12161 16201 12173 16235
rect 12207 16232 12219 16235
rect 12342 16232 12348 16244
rect 12207 16204 12348 16232
rect 12207 16201 12219 16204
rect 12161 16195 12219 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 15427 16235 15485 16241
rect 15427 16201 15439 16235
rect 15473 16232 15485 16235
rect 16758 16232 16764 16244
rect 15473 16204 16764 16232
rect 15473 16201 15485 16204
rect 15427 16195 15485 16201
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 18782 16192 18788 16244
rect 18840 16232 18846 16244
rect 20165 16235 20223 16241
rect 20165 16232 20177 16235
rect 18840 16204 20177 16232
rect 18840 16192 18846 16204
rect 20165 16201 20177 16204
rect 20211 16201 20223 16235
rect 20165 16195 20223 16201
rect 21637 16235 21695 16241
rect 21637 16201 21649 16235
rect 21683 16232 21695 16235
rect 21910 16232 21916 16244
rect 21683 16204 21916 16232
rect 21683 16201 21695 16204
rect 21637 16195 21695 16201
rect 5166 16124 5172 16176
rect 5224 16164 5230 16176
rect 7561 16167 7619 16173
rect 7561 16164 7573 16167
rect 5224 16136 7573 16164
rect 5224 16124 5230 16136
rect 7561 16133 7573 16136
rect 7607 16164 7619 16167
rect 7834 16164 7840 16176
rect 7607 16136 7840 16164
rect 7607 16133 7619 16136
rect 7561 16127 7619 16133
rect 7834 16124 7840 16136
rect 7892 16164 7898 16176
rect 11238 16164 11244 16176
rect 7892 16136 11244 16164
rect 7892 16124 7898 16136
rect 11238 16124 11244 16136
rect 11296 16124 11302 16176
rect 15105 16167 15163 16173
rect 15105 16164 15117 16167
rect 11532 16136 15117 16164
rect 5905 16099 5963 16105
rect 5905 16065 5917 16099
rect 5951 16096 5963 16099
rect 8294 16096 8300 16108
rect 5951 16068 8300 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 8389 16099 8447 16105
rect 8389 16065 8401 16099
rect 8435 16096 8447 16099
rect 9674 16096 9680 16108
rect 8435 16068 9680 16096
rect 8435 16065 8447 16068
rect 8389 16059 8447 16065
rect 9674 16056 9680 16068
rect 9732 16056 9738 16108
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16096 10011 16099
rect 10686 16096 10692 16108
rect 9999 16068 10692 16096
rect 9999 16065 10011 16068
rect 9953 16059 10011 16065
rect 10686 16056 10692 16068
rect 10744 16096 10750 16108
rect 11422 16096 11428 16108
rect 10744 16068 11428 16096
rect 10744 16056 10750 16068
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 11532 16105 11560 16136
rect 15105 16133 15117 16136
rect 15151 16164 15163 16167
rect 15286 16164 15292 16176
rect 15151 16136 15292 16164
rect 15151 16133 15163 16136
rect 15105 16127 15163 16133
rect 15286 16124 15292 16136
rect 15344 16124 15350 16176
rect 16114 16164 16120 16176
rect 16075 16136 16120 16164
rect 16114 16124 16120 16136
rect 16172 16164 16178 16176
rect 18874 16164 18880 16176
rect 16172 16136 18880 16164
rect 16172 16124 16178 16136
rect 18874 16124 18880 16136
rect 18932 16124 18938 16176
rect 11517 16099 11575 16105
rect 11517 16065 11529 16099
rect 11563 16065 11575 16099
rect 13633 16099 13691 16105
rect 13633 16096 13645 16099
rect 11517 16059 11575 16065
rect 11624 16068 13645 16096
rect 1210 15988 1216 16040
rect 1268 16028 1274 16040
rect 1800 16031 1858 16037
rect 1800 16028 1812 16031
rect 1268 16000 1812 16028
rect 1268 15988 1274 16000
rect 1800 15997 1812 16000
rect 1846 16028 1858 16031
rect 2225 16031 2283 16037
rect 2225 16028 2237 16031
rect 1846 16000 2237 16028
rect 1846 15997 1858 16000
rect 1800 15991 1858 15997
rect 2225 15997 2237 16000
rect 2271 15997 2283 16031
rect 2225 15991 2283 15997
rect 2682 15988 2688 16040
rect 2740 16028 2746 16040
rect 2777 16031 2835 16037
rect 2777 16028 2789 16031
rect 2740 16000 2789 16028
rect 2740 15988 2746 16000
rect 2777 15997 2789 16000
rect 2823 15997 2835 16031
rect 7834 16028 7840 16040
rect 7795 16000 7840 16028
rect 2777 15991 2835 15997
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 8478 16028 8484 16040
rect 8159 16000 8484 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 5258 15960 5264 15972
rect 5219 15932 5264 15960
rect 5258 15920 5264 15932
rect 5316 15920 5322 15972
rect 5350 15920 5356 15972
rect 5408 15960 5414 15972
rect 8128 15960 8156 15991
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 10597 16031 10655 16037
rect 10597 15997 10609 16031
rect 10643 16028 10655 16031
rect 11054 16028 11060 16040
rect 10643 16000 11060 16028
rect 10643 15997 10655 16000
rect 10597 15991 10655 15997
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 11238 16028 11244 16040
rect 11199 16000 11244 16028
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 5408 15932 5453 15960
rect 7208 15932 8156 15960
rect 5408 15920 5414 15932
rect 7208 15904 7236 15932
rect 9030 15920 9036 15972
rect 9088 15960 9094 15972
rect 9309 15963 9367 15969
rect 9309 15960 9321 15963
rect 9088 15932 9321 15960
rect 9088 15920 9094 15932
rect 9309 15929 9321 15932
rect 9355 15929 9367 15963
rect 9309 15923 9367 15929
rect 9398 15920 9404 15972
rect 9456 15960 9462 15972
rect 9456 15932 9501 15960
rect 9456 15920 9462 15932
rect 10042 15920 10048 15972
rect 10100 15960 10106 15972
rect 11624 15960 11652 16068
rect 13633 16065 13645 16068
rect 13679 16096 13691 16099
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 13679 16068 14565 16096
rect 13679 16065 13691 16068
rect 13633 16059 13691 16065
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 17034 16096 17040 16108
rect 14553 16059 14611 16065
rect 15212 16068 17040 16096
rect 14274 15988 14280 16040
rect 14332 16028 14338 16040
rect 15212 16028 15240 16068
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 17770 16096 17776 16108
rect 17731 16068 17776 16096
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16096 18567 16099
rect 20180 16096 20208 16195
rect 21910 16192 21916 16204
rect 21968 16192 21974 16244
rect 22370 16232 22376 16244
rect 22331 16204 22376 16232
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 23014 16232 23020 16244
rect 22975 16204 23020 16232
rect 23014 16192 23020 16204
rect 23072 16192 23078 16244
rect 23934 16232 23940 16244
rect 23895 16204 23940 16232
rect 23934 16192 23940 16204
rect 23992 16192 23998 16244
rect 20717 16099 20775 16105
rect 20717 16096 20729 16099
rect 18555 16068 19472 16096
rect 20180 16068 20729 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 19444 16040 19472 16068
rect 20717 16065 20729 16068
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 14332 16000 15240 16028
rect 15356 16031 15414 16037
rect 14332 15988 14338 16000
rect 15356 15997 15368 16031
rect 15402 16028 15414 16031
rect 15838 16028 15844 16040
rect 15402 16000 15844 16028
rect 15402 15997 15414 16000
rect 15356 15991 15414 15997
rect 15838 15988 15844 16000
rect 15896 15988 15902 16040
rect 18966 16028 18972 16040
rect 18927 16000 18972 16028
rect 18966 15988 18972 16000
rect 19024 15988 19030 16040
rect 19426 15988 19432 16040
rect 19484 16028 19490 16040
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 19484 16000 19901 16028
rect 19484 15988 19490 16000
rect 19889 15997 19901 16000
rect 19935 16028 19947 16031
rect 21634 16028 21640 16040
rect 19935 16000 21640 16028
rect 19935 15997 19947 16000
rect 19889 15991 19947 15997
rect 21634 15988 21640 16000
rect 21692 15988 21698 16040
rect 13722 15960 13728 15972
rect 10100 15932 11652 15960
rect 13683 15932 13728 15960
rect 10100 15920 10106 15932
rect 13722 15920 13728 15932
rect 13780 15920 13786 15972
rect 16390 15960 16396 15972
rect 16351 15932 16396 15960
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 16485 15963 16543 15969
rect 16485 15929 16497 15963
rect 16531 15929 16543 15963
rect 16485 15923 16543 15929
rect 2685 15895 2743 15901
rect 2685 15861 2697 15895
rect 2731 15892 2743 15895
rect 2774 15892 2780 15904
rect 2731 15864 2780 15892
rect 2731 15861 2743 15864
rect 2685 15855 2743 15861
rect 2774 15852 2780 15864
rect 2832 15892 2838 15904
rect 3145 15895 3203 15901
rect 3145 15892 3157 15895
rect 2832 15864 3157 15892
rect 2832 15852 2838 15864
rect 3145 15861 3157 15864
rect 3191 15861 3203 15895
rect 4982 15892 4988 15904
rect 4943 15864 4988 15892
rect 3145 15855 3203 15861
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 7190 15892 7196 15904
rect 7151 15864 7196 15892
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 9125 15895 9183 15901
rect 9125 15861 9137 15895
rect 9171 15892 9183 15895
rect 9416 15892 9444 15920
rect 9171 15864 9444 15892
rect 9171 15861 9183 15864
rect 9125 15855 9183 15861
rect 10134 15852 10140 15904
rect 10192 15892 10198 15904
rect 10229 15895 10287 15901
rect 10229 15892 10241 15895
rect 10192 15864 10241 15892
rect 10192 15852 10198 15864
rect 10229 15861 10241 15864
rect 10275 15861 10287 15895
rect 10229 15855 10287 15861
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 12437 15895 12495 15901
rect 12437 15892 12449 15895
rect 10744 15864 12449 15892
rect 10744 15852 10750 15864
rect 12437 15861 12449 15864
rect 12483 15861 12495 15895
rect 12437 15855 12495 15861
rect 12618 15852 12624 15904
rect 12676 15892 12682 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12676 15864 12909 15892
rect 12676 15852 12682 15864
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 12897 15855 12955 15861
rect 13449 15895 13507 15901
rect 13449 15861 13461 15895
rect 13495 15892 13507 15895
rect 13740 15892 13768 15920
rect 13495 15864 13768 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 16298 15892 16304 15904
rect 15712 15864 16304 15892
rect 15712 15852 15718 15864
rect 16298 15852 16304 15864
rect 16356 15892 16362 15904
rect 16500 15892 16528 15923
rect 18874 15920 18880 15972
rect 18932 15960 18938 15972
rect 19290 15963 19348 15969
rect 19290 15960 19302 15963
rect 18932 15932 19302 15960
rect 18932 15920 18938 15932
rect 19290 15929 19302 15932
rect 19336 15960 19348 15963
rect 20533 15963 20591 15969
rect 20533 15960 20545 15963
rect 19336 15932 20545 15960
rect 19336 15929 19348 15932
rect 19290 15923 19348 15929
rect 20533 15929 20545 15932
rect 20579 15960 20591 15963
rect 21038 15963 21096 15969
rect 21038 15960 21050 15963
rect 20579 15932 21050 15960
rect 20579 15929 20591 15932
rect 20533 15923 20591 15929
rect 21038 15929 21050 15932
rect 21084 15929 21096 15963
rect 21038 15923 21096 15929
rect 21174 15920 21180 15972
rect 21232 15960 21238 15972
rect 22465 15963 22523 15969
rect 22465 15960 22477 15963
rect 21232 15932 22477 15960
rect 21232 15920 21238 15932
rect 22465 15929 22477 15932
rect 22511 15929 22523 15963
rect 22465 15923 22523 15929
rect 17310 15892 17316 15904
rect 16356 15864 16528 15892
rect 17271 15864 17316 15892
rect 16356 15852 16362 15864
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 21634 15852 21640 15904
rect 21692 15892 21698 15904
rect 22005 15895 22063 15901
rect 22005 15892 22017 15895
rect 21692 15864 22017 15892
rect 21692 15852 21698 15864
rect 22005 15861 22017 15864
rect 22051 15892 22063 15895
rect 23014 15892 23020 15904
rect 22051 15864 23020 15892
rect 22051 15861 22063 15864
rect 22005 15855 22063 15861
rect 23014 15852 23020 15864
rect 23072 15852 23078 15904
rect 24026 15852 24032 15904
rect 24084 15892 24090 15904
rect 27614 15892 27620 15904
rect 24084 15864 27620 15892
rect 24084 15852 24090 15864
rect 27614 15852 27620 15864
rect 27672 15852 27678 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 5258 15648 5264 15700
rect 5316 15688 5322 15700
rect 5997 15691 6055 15697
rect 5997 15688 6009 15691
rect 5316 15660 6009 15688
rect 5316 15648 5322 15660
rect 5997 15657 6009 15660
rect 6043 15688 6055 15691
rect 7374 15688 7380 15700
rect 6043 15660 7380 15688
rect 6043 15657 6055 15660
rect 5997 15651 6055 15657
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 9674 15688 9680 15700
rect 9539 15660 9680 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10873 15691 10931 15697
rect 10873 15657 10885 15691
rect 10919 15688 10931 15691
rect 11238 15688 11244 15700
rect 10919 15660 11244 15688
rect 10919 15657 10931 15660
rect 10873 15651 10931 15657
rect 11238 15648 11244 15660
rect 11296 15648 11302 15700
rect 13262 15688 13268 15700
rect 13223 15660 13268 15688
rect 13262 15648 13268 15660
rect 13320 15648 13326 15700
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 14274 15688 14280 15700
rect 13872 15660 13917 15688
rect 14235 15660 14280 15688
rect 13872 15648 13878 15660
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 19889 15691 19947 15697
rect 19889 15657 19901 15691
rect 19935 15688 19947 15691
rect 19978 15688 19984 15700
rect 19935 15660 19984 15688
rect 19935 15657 19947 15660
rect 19889 15651 19947 15657
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 24762 15688 24768 15700
rect 24723 15660 24768 15688
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 3145 15623 3203 15629
rect 3145 15589 3157 15623
rect 3191 15620 3203 15623
rect 3326 15620 3332 15632
rect 3191 15592 3332 15620
rect 3191 15589 3203 15592
rect 3145 15583 3203 15589
rect 3326 15580 3332 15592
rect 3384 15580 3390 15632
rect 7190 15580 7196 15632
rect 7248 15620 7254 15632
rect 7653 15623 7711 15629
rect 7653 15620 7665 15623
rect 7248 15592 7665 15620
rect 7248 15580 7254 15592
rect 7653 15589 7665 15592
rect 7699 15620 7711 15623
rect 7699 15592 8524 15620
rect 7699 15589 7711 15592
rect 7653 15583 7711 15589
rect 8496 15564 8524 15592
rect 8846 15580 8852 15632
rect 8904 15620 8910 15632
rect 9769 15623 9827 15629
rect 9769 15620 9781 15623
rect 8904 15592 9781 15620
rect 8904 15580 8910 15592
rect 9769 15589 9781 15592
rect 9815 15589 9827 15623
rect 9769 15583 9827 15589
rect 9861 15623 9919 15629
rect 9861 15589 9873 15623
rect 9907 15620 9919 15623
rect 10778 15620 10784 15632
rect 9907 15592 10784 15620
rect 9907 15589 9919 15592
rect 9861 15583 9919 15589
rect 10778 15580 10784 15592
rect 10836 15580 10842 15632
rect 11422 15620 11428 15632
rect 11383 15592 11428 15620
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 11974 15620 11980 15632
rect 11935 15592 11980 15620
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 15654 15580 15660 15632
rect 15712 15620 15718 15632
rect 15749 15623 15807 15629
rect 15749 15620 15761 15623
rect 15712 15592 15761 15620
rect 15712 15580 15718 15592
rect 15749 15589 15761 15592
rect 15795 15589 15807 15623
rect 21174 15620 21180 15632
rect 21135 15592 21180 15620
rect 15749 15583 15807 15589
rect 21174 15580 21180 15592
rect 21232 15580 21238 15632
rect 21269 15623 21327 15629
rect 21269 15589 21281 15623
rect 21315 15620 21327 15623
rect 21910 15620 21916 15632
rect 21315 15592 21916 15620
rect 21315 15589 21327 15592
rect 21269 15583 21327 15589
rect 21910 15580 21916 15592
rect 21968 15580 21974 15632
rect 2406 15552 2412 15564
rect 2367 15524 2412 15552
rect 2406 15512 2412 15524
rect 2464 15512 2470 15564
rect 2590 15512 2596 15564
rect 2648 15552 2654 15564
rect 2685 15555 2743 15561
rect 2685 15552 2697 15555
rect 2648 15524 2697 15552
rect 2648 15512 2654 15524
rect 2685 15521 2697 15524
rect 2731 15552 2743 15555
rect 3050 15552 3056 15564
rect 2731 15524 3056 15552
rect 2731 15521 2743 15524
rect 2685 15515 2743 15521
rect 3050 15512 3056 15524
rect 3108 15552 3114 15564
rect 4062 15552 4068 15564
rect 3108 15524 4068 15552
rect 3108 15512 3114 15524
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 5442 15552 5448 15564
rect 5403 15524 5448 15552
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 6454 15552 6460 15564
rect 6415 15524 6460 15552
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15521 6791 15555
rect 8018 15552 8024 15564
rect 7979 15524 8024 15552
rect 6733 15515 6791 15521
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 3786 15484 3792 15496
rect 2363 15456 3792 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 4893 15487 4951 15493
rect 4893 15484 4905 15487
rect 4126 15456 4905 15484
rect 2498 15416 2504 15428
rect 2459 15388 2504 15416
rect 2498 15376 2504 15388
rect 2556 15416 2562 15428
rect 3694 15416 3700 15428
rect 2556 15388 3700 15416
rect 2556 15376 2562 15388
rect 3694 15376 3700 15388
rect 3752 15416 3758 15428
rect 4126 15416 4154 15456
rect 4893 15453 4905 15456
rect 4939 15453 4951 15487
rect 6748 15484 6776 15515
rect 8018 15512 8024 15524
rect 8076 15552 8082 15564
rect 8202 15552 8208 15564
rect 8076 15524 8208 15552
rect 8076 15512 8082 15524
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8478 15552 8484 15564
rect 8391 15524 8484 15552
rect 8478 15512 8484 15524
rect 8536 15512 8542 15564
rect 12526 15512 12532 15564
rect 12584 15552 12590 15564
rect 12713 15555 12771 15561
rect 12713 15552 12725 15555
rect 12584 15524 12725 15552
rect 12584 15512 12590 15524
rect 12713 15521 12725 15524
rect 12759 15552 12771 15555
rect 12805 15555 12863 15561
rect 12805 15552 12817 15555
rect 12759 15524 12817 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12805 15521 12817 15524
rect 12851 15521 12863 15555
rect 13078 15552 13084 15564
rect 13039 15524 13084 15552
rect 12805 15515 12863 15521
rect 13078 15512 13084 15524
rect 13136 15512 13142 15564
rect 17678 15512 17684 15564
rect 17736 15552 17742 15564
rect 17773 15555 17831 15561
rect 17773 15552 17785 15555
rect 17736 15524 17785 15552
rect 17736 15512 17742 15524
rect 17773 15521 17785 15524
rect 17819 15521 17831 15555
rect 18230 15552 18236 15564
rect 18191 15524 18236 15552
rect 17773 15515 17831 15521
rect 18230 15512 18236 15524
rect 18288 15512 18294 15564
rect 19337 15555 19395 15561
rect 19337 15552 19349 15555
rect 18340 15524 19349 15552
rect 4893 15447 4951 15453
rect 6288 15456 6776 15484
rect 7193 15487 7251 15493
rect 3752 15388 4154 15416
rect 3752 15376 3758 15388
rect 5074 15376 5080 15428
rect 5132 15416 5138 15428
rect 6288 15425 6316 15456
rect 7193 15453 7205 15487
rect 7239 15484 7251 15487
rect 7834 15484 7840 15496
rect 7239 15456 7840 15484
rect 7239 15453 7251 15456
rect 7193 15447 7251 15453
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 9398 15484 9404 15496
rect 8803 15456 9404 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 10042 15484 10048 15496
rect 10003 15456 10048 15484
rect 10042 15444 10048 15456
rect 10100 15484 10106 15496
rect 11330 15484 11336 15496
rect 10100 15456 11336 15484
rect 10100 15444 10106 15456
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15484 15715 15487
rect 15838 15484 15844 15496
rect 15703 15456 15844 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 15838 15444 15844 15456
rect 15896 15484 15902 15496
rect 18340 15484 18368 15524
rect 19337 15521 19349 15524
rect 19383 15521 19395 15555
rect 19337 15515 19395 15521
rect 21818 15512 21824 15564
rect 21876 15552 21882 15564
rect 22649 15555 22707 15561
rect 22649 15552 22661 15555
rect 21876 15524 22661 15552
rect 21876 15512 21882 15524
rect 22649 15521 22661 15524
rect 22695 15521 22707 15555
rect 22649 15515 22707 15521
rect 22925 15555 22983 15561
rect 22925 15521 22937 15555
rect 22971 15552 22983 15555
rect 23290 15552 23296 15564
rect 22971 15524 23296 15552
rect 22971 15521 22983 15524
rect 22925 15515 22983 15521
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 24118 15512 24124 15564
rect 24176 15552 24182 15564
rect 24581 15555 24639 15561
rect 24581 15552 24593 15555
rect 24176 15524 24593 15552
rect 24176 15512 24182 15524
rect 24581 15521 24593 15524
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 18506 15484 18512 15496
rect 15896 15456 18368 15484
rect 18467 15456 18512 15484
rect 15896 15444 15902 15456
rect 18506 15444 18512 15456
rect 18564 15444 18570 15496
rect 21542 15484 21548 15496
rect 21503 15456 21548 15484
rect 21542 15444 21548 15456
rect 21600 15444 21606 15496
rect 23106 15484 23112 15496
rect 23067 15456 23112 15484
rect 23106 15444 23112 15456
rect 23164 15444 23170 15496
rect 6273 15419 6331 15425
rect 6273 15416 6285 15419
rect 5132 15388 6285 15416
rect 5132 15376 5138 15388
rect 6273 15385 6285 15388
rect 6319 15385 6331 15419
rect 6546 15416 6552 15428
rect 6507 15388 6552 15416
rect 6273 15379 6331 15385
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 12897 15419 12955 15425
rect 12897 15385 12909 15419
rect 12943 15416 12955 15419
rect 12986 15416 12992 15428
rect 12943 15388 12992 15416
rect 12943 15385 12955 15388
rect 12897 15379 12955 15385
rect 12986 15376 12992 15388
rect 13044 15376 13050 15428
rect 16206 15416 16212 15428
rect 16167 15388 16212 15416
rect 16206 15376 16212 15388
rect 16264 15376 16270 15428
rect 22741 15419 22799 15425
rect 22741 15385 22753 15419
rect 22787 15416 22799 15419
rect 22922 15416 22928 15428
rect 22787 15388 22928 15416
rect 22787 15385 22799 15388
rect 22741 15379 22799 15385
rect 22922 15376 22928 15388
rect 22980 15376 22986 15428
rect 2866 15308 2872 15360
rect 2924 15348 2930 15360
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 2924 15320 3433 15348
rect 2924 15308 2930 15320
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 9030 15348 9036 15360
rect 8991 15320 9036 15348
rect 3421 15311 3479 15317
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 12250 15348 12256 15360
rect 12211 15320 12256 15348
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 16390 15308 16396 15360
rect 16448 15348 16454 15360
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 16448 15320 16681 15348
rect 16448 15308 16454 15320
rect 16669 15317 16681 15320
rect 16715 15348 16727 15351
rect 17678 15348 17684 15360
rect 16715 15320 17684 15348
rect 16715 15317 16727 15320
rect 16669 15311 16727 15317
rect 17678 15308 17684 15320
rect 17736 15308 17742 15360
rect 18966 15348 18972 15360
rect 18927 15320 18972 15348
rect 18966 15308 18972 15320
rect 19024 15308 19030 15360
rect 20438 15348 20444 15360
rect 20399 15320 20444 15348
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 22186 15348 22192 15360
rect 22147 15320 22192 15348
rect 22186 15308 22192 15320
rect 22244 15308 22250 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1765 15147 1823 15153
rect 1765 15113 1777 15147
rect 1811 15144 1823 15147
rect 2590 15144 2596 15156
rect 1811 15116 2596 15144
rect 1811 15113 1823 15116
rect 1765 15107 1823 15113
rect 2590 15104 2596 15116
rect 2648 15104 2654 15156
rect 8478 15104 8484 15156
rect 8536 15144 8542 15156
rect 9585 15147 9643 15153
rect 9585 15144 9597 15147
rect 8536 15116 9597 15144
rect 8536 15104 8542 15116
rect 9585 15113 9597 15116
rect 9631 15113 9643 15147
rect 9585 15107 9643 15113
rect 10778 15104 10784 15156
rect 10836 15144 10842 15156
rect 11333 15147 11391 15153
rect 11333 15144 11345 15147
rect 10836 15116 11345 15144
rect 10836 15104 10842 15116
rect 11333 15113 11345 15116
rect 11379 15113 11391 15147
rect 14185 15147 14243 15153
rect 14185 15144 14197 15147
rect 11333 15107 11391 15113
rect 13786 15116 14197 15144
rect 11057 15079 11115 15085
rect 11057 15045 11069 15079
rect 11103 15076 11115 15079
rect 11422 15076 11428 15088
rect 11103 15048 11428 15076
rect 11103 15045 11115 15048
rect 11057 15039 11115 15045
rect 11422 15036 11428 15048
rect 11480 15076 11486 15088
rect 11701 15079 11759 15085
rect 11701 15076 11713 15079
rect 11480 15048 11713 15076
rect 11480 15036 11486 15048
rect 11701 15045 11713 15048
rect 11747 15045 11759 15079
rect 11701 15039 11759 15045
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 15008 2191 15011
rect 2406 15008 2412 15020
rect 2179 14980 2412 15008
rect 2179 14977 2191 14980
rect 2133 14971 2191 14977
rect 2406 14968 2412 14980
rect 2464 15008 2470 15020
rect 2501 15011 2559 15017
rect 2501 15008 2513 15011
rect 2464 14980 2513 15008
rect 2464 14968 2470 14980
rect 2501 14977 2513 14980
rect 2547 15008 2559 15011
rect 8386 15008 8392 15020
rect 2547 14980 6132 15008
rect 8299 14980 8392 15008
rect 2547 14977 2559 14980
rect 2501 14971 2559 14977
rect 2866 14940 2872 14952
rect 2827 14912 2872 14940
rect 2866 14900 2872 14912
rect 2924 14900 2930 14952
rect 3329 14943 3387 14949
rect 3329 14909 3341 14943
rect 3375 14909 3387 14943
rect 3329 14903 3387 14909
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14940 3663 14943
rect 3694 14940 3700 14952
rect 3651 14912 3700 14940
rect 3651 14909 3663 14912
rect 3605 14903 3663 14909
rect 3344 14872 3372 14903
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 3988 14949 4016 14980
rect 6104 14952 6132 14980
rect 8386 14968 8392 14980
rect 8444 15008 8450 15020
rect 9030 15008 9036 15020
rect 8444 14980 9036 15008
rect 8444 14968 8450 14980
rect 9030 14968 9036 14980
rect 9088 14968 9094 15020
rect 13786 15008 13814 15116
rect 14185 15113 14197 15116
rect 14231 15144 14243 15147
rect 16301 15147 16359 15153
rect 16301 15144 16313 15147
rect 14231 15116 16313 15144
rect 14231 15113 14243 15116
rect 14185 15107 14243 15113
rect 16301 15113 16313 15116
rect 16347 15144 16359 15147
rect 16482 15144 16488 15156
rect 16347 15116 16488 15144
rect 16347 15113 16359 15116
rect 16301 15107 16359 15113
rect 16482 15104 16488 15116
rect 16540 15144 16546 15156
rect 16850 15144 16856 15156
rect 16540 15116 16856 15144
rect 16540 15104 16546 15116
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 17586 15104 17592 15156
rect 17644 15144 17650 15156
rect 17681 15147 17739 15153
rect 17681 15144 17693 15147
rect 17644 15116 17693 15144
rect 17644 15104 17650 15116
rect 17681 15113 17693 15116
rect 17727 15144 17739 15147
rect 17773 15147 17831 15153
rect 17773 15144 17785 15147
rect 17727 15116 17785 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 17773 15113 17785 15116
rect 17819 15113 17831 15147
rect 17773 15107 17831 15113
rect 21174 15104 21180 15156
rect 21232 15144 21238 15156
rect 21361 15147 21419 15153
rect 21361 15144 21373 15147
rect 21232 15116 21373 15144
rect 21232 15104 21238 15116
rect 21361 15113 21373 15116
rect 21407 15113 21419 15147
rect 21726 15144 21732 15156
rect 21687 15116 21732 15144
rect 21361 15107 21419 15113
rect 21726 15104 21732 15116
rect 21784 15104 21790 15156
rect 15565 15079 15623 15085
rect 15565 15045 15577 15079
rect 15611 15076 15623 15079
rect 16390 15076 16396 15088
rect 15611 15048 16396 15076
rect 15611 15045 15623 15048
rect 15565 15039 15623 15045
rect 16390 15036 16396 15048
rect 16448 15076 16454 15088
rect 17310 15076 17316 15088
rect 16448 15048 17316 15076
rect 16448 15036 16454 15048
rect 17310 15036 17316 15048
rect 17368 15036 17374 15088
rect 22557 15079 22615 15085
rect 22557 15076 22569 15079
rect 20456 15048 22569 15076
rect 20456 15020 20484 15048
rect 22557 15045 22569 15048
rect 22603 15076 22615 15079
rect 22830 15076 22836 15088
rect 22603 15048 22836 15076
rect 22603 15045 22615 15048
rect 22557 15039 22615 15045
rect 22830 15036 22836 15048
rect 22888 15036 22894 15088
rect 13556 14980 13814 15008
rect 17129 15011 17187 15017
rect 13556 14952 13584 14980
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 18966 15008 18972 15020
rect 17175 14980 18972 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 20438 15008 20444 15020
rect 20399 14980 20444 15008
rect 20438 14968 20444 14980
rect 20496 14968 20502 15020
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 15008 22063 15011
rect 22186 15008 22192 15020
rect 22051 14980 22192 15008
rect 22051 14977 22063 14980
rect 22005 14971 22063 14977
rect 22186 14968 22192 14980
rect 22244 15008 22250 15020
rect 23799 15011 23857 15017
rect 23799 15008 23811 15011
rect 22244 14980 23811 15008
rect 22244 14968 22250 14980
rect 23799 14977 23811 14980
rect 23845 14977 23857 15011
rect 23799 14971 23857 14977
rect 3973 14943 4031 14949
rect 3973 14909 3985 14943
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4985 14943 5043 14949
rect 4985 14940 4997 14943
rect 4120 14912 4997 14940
rect 4120 14900 4126 14912
rect 4985 14909 4997 14912
rect 5031 14940 5043 14943
rect 5629 14943 5687 14949
rect 5629 14940 5641 14943
rect 5031 14912 5641 14940
rect 5031 14909 5043 14912
rect 4985 14903 5043 14909
rect 5629 14909 5641 14912
rect 5675 14940 5687 14943
rect 5902 14940 5908 14952
rect 5675 14912 5908 14940
rect 5675 14909 5687 14912
rect 5629 14903 5687 14909
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 6086 14940 6092 14952
rect 6047 14912 6092 14940
rect 6086 14900 6092 14912
rect 6144 14940 6150 14952
rect 6454 14940 6460 14952
rect 6144 14912 6460 14940
rect 6144 14900 6150 14912
rect 6454 14900 6460 14912
rect 6512 14940 6518 14952
rect 6917 14943 6975 14949
rect 6917 14940 6929 14943
rect 6512 14912 6929 14940
rect 6512 14900 6518 14912
rect 6917 14909 6929 14912
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 9398 14900 9404 14952
rect 9456 14940 9462 14952
rect 10137 14943 10195 14949
rect 10137 14940 10149 14943
rect 9456 14912 10149 14940
rect 9456 14900 9462 14912
rect 10137 14909 10149 14912
rect 10183 14909 10195 14943
rect 10137 14903 10195 14909
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 12253 14943 12311 14949
rect 12253 14940 12265 14943
rect 11112 14912 12265 14940
rect 11112 14900 11118 14912
rect 12253 14909 12265 14912
rect 12299 14940 12311 14943
rect 13262 14940 13268 14952
rect 12299 14912 13268 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13538 14940 13544 14952
rect 13499 14912 13544 14940
rect 13538 14900 13544 14912
rect 13596 14900 13602 14952
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14940 13875 14943
rect 14642 14940 14648 14952
rect 13863 14912 14648 14940
rect 13863 14909 13875 14912
rect 13817 14903 13875 14909
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 16482 14940 16488 14952
rect 16443 14912 16488 14940
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 17681 14943 17739 14949
rect 17681 14909 17693 14943
rect 17727 14940 17739 14943
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17727 14912 18061 14940
rect 17727 14909 17739 14912
rect 17681 14903 17739 14909
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 18509 14943 18567 14949
rect 18509 14909 18521 14943
rect 18555 14940 18567 14943
rect 19061 14943 19119 14949
rect 19061 14940 19073 14943
rect 18555 14912 19073 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 19061 14909 19073 14912
rect 19107 14940 19119 14943
rect 19242 14940 19248 14952
rect 19107 14912 19248 14940
rect 19107 14909 19119 14912
rect 19061 14903 19119 14909
rect 3510 14872 3516 14884
rect 3344 14844 3516 14872
rect 3510 14832 3516 14844
rect 3568 14832 3574 14884
rect 5074 14872 5080 14884
rect 5035 14844 5080 14872
rect 5074 14832 5080 14844
rect 5132 14832 5138 14884
rect 5350 14832 5356 14884
rect 5408 14872 5414 14884
rect 6825 14875 6883 14881
rect 6825 14872 6837 14875
rect 5408 14844 6837 14872
rect 5408 14832 5414 14844
rect 6825 14841 6837 14844
rect 6871 14841 6883 14875
rect 8294 14872 8300 14884
rect 8207 14844 8300 14872
rect 6825 14835 6883 14841
rect 8294 14832 8300 14844
rect 8352 14872 8358 14884
rect 8751 14875 8809 14881
rect 8751 14872 8763 14875
rect 8352 14844 8763 14872
rect 8352 14832 8358 14844
rect 8751 14841 8763 14844
rect 8797 14872 8809 14875
rect 10045 14875 10103 14881
rect 10045 14872 10057 14875
rect 8797 14844 10057 14872
rect 8797 14841 8809 14844
rect 8751 14835 8809 14841
rect 10045 14841 10057 14844
rect 10091 14872 10103 14875
rect 10499 14875 10557 14881
rect 10499 14872 10511 14875
rect 10091 14844 10511 14872
rect 10091 14841 10103 14844
rect 10045 14835 10103 14841
rect 10152 14816 10180 14844
rect 10499 14841 10511 14844
rect 10545 14872 10557 14875
rect 14461 14875 14519 14881
rect 14461 14872 14473 14875
rect 10545 14844 13676 14872
rect 10545 14841 10557 14844
rect 10499 14835 10557 14841
rect 13648 14816 13676 14844
rect 14016 14844 14473 14872
rect 2682 14804 2688 14816
rect 2643 14776 2688 14804
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 4617 14807 4675 14813
rect 4617 14773 4629 14807
rect 4663 14804 4675 14807
rect 5442 14804 5448 14816
rect 4663 14776 5448 14804
rect 4663 14773 4675 14776
rect 4617 14767 4675 14773
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 5994 14764 6000 14816
rect 6052 14804 6058 14816
rect 7837 14807 7895 14813
rect 7837 14804 7849 14807
rect 6052 14776 7849 14804
rect 6052 14764 6058 14776
rect 7837 14773 7849 14776
rect 7883 14804 7895 14807
rect 8018 14804 8024 14816
rect 7883 14776 8024 14804
rect 7883 14773 7895 14776
rect 7837 14767 7895 14773
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 9306 14804 9312 14816
rect 9267 14776 9312 14804
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 10134 14764 10140 14816
rect 10192 14764 10198 14816
rect 12897 14807 12955 14813
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 12986 14804 12992 14816
rect 12943 14776 12992 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 13630 14764 13636 14816
rect 13688 14804 13694 14816
rect 14016 14804 14044 14844
rect 14461 14841 14473 14844
rect 14507 14872 14519 14875
rect 14966 14875 15024 14881
rect 14966 14872 14978 14875
rect 14507 14844 14978 14872
rect 14507 14841 14519 14844
rect 14461 14835 14519 14841
rect 14966 14841 14978 14844
rect 15012 14841 15024 14875
rect 16868 14872 16896 14903
rect 17586 14872 17592 14884
rect 14966 14835 15024 14841
rect 15856 14844 17592 14872
rect 13688 14776 14044 14804
rect 13688 14764 13694 14776
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 15856 14813 15884 14844
rect 17586 14832 17592 14844
rect 17644 14872 17650 14884
rect 18230 14872 18236 14884
rect 17644 14844 18236 14872
rect 17644 14832 17650 14844
rect 18230 14832 18236 14844
rect 18288 14872 18294 14884
rect 18524 14872 18552 14903
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 23712 14943 23770 14949
rect 23712 14909 23724 14943
rect 23758 14909 23770 14943
rect 23712 14903 23770 14909
rect 18782 14872 18788 14884
rect 18288 14844 18552 14872
rect 18743 14844 18788 14872
rect 18288 14832 18294 14844
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 20530 14832 20536 14884
rect 20588 14872 20594 14884
rect 21085 14875 21143 14881
rect 20588 14844 20633 14872
rect 20588 14832 20594 14844
rect 21085 14841 21097 14875
rect 21131 14872 21143 14875
rect 21266 14872 21272 14884
rect 21131 14844 21272 14872
rect 21131 14841 21143 14844
rect 21085 14835 21143 14841
rect 21266 14832 21272 14844
rect 21324 14832 21330 14884
rect 22002 14872 22008 14884
rect 21560 14844 22008 14872
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 14792 14776 15853 14804
rect 14792 14764 14798 14776
rect 15841 14773 15853 14776
rect 15887 14773 15899 14807
rect 15841 14767 15899 14773
rect 17497 14807 17555 14813
rect 17497 14773 17509 14807
rect 17543 14804 17555 14807
rect 17770 14804 17776 14816
rect 17543 14776 17776 14804
rect 17543 14773 17555 14776
rect 17497 14767 17555 14773
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 20257 14807 20315 14813
rect 20257 14773 20269 14807
rect 20303 14804 20315 14807
rect 21560 14804 21588 14844
rect 22002 14832 22008 14844
rect 22060 14872 22066 14884
rect 22097 14875 22155 14881
rect 22097 14872 22109 14875
rect 22060 14844 22109 14872
rect 22060 14832 22066 14844
rect 22097 14841 22109 14844
rect 22143 14841 22155 14875
rect 22097 14835 22155 14841
rect 22738 14832 22744 14884
rect 22796 14872 22802 14884
rect 23727 14872 23755 14903
rect 24118 14900 24124 14952
rect 24176 14940 24182 14952
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 24176 14912 24593 14940
rect 24176 14900 24182 14912
rect 24581 14909 24593 14912
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 22796 14844 24256 14872
rect 22796 14832 22802 14844
rect 22922 14804 22928 14816
rect 20303 14776 21588 14804
rect 22883 14776 22928 14804
rect 20303 14773 20315 14776
rect 20257 14767 20315 14773
rect 22922 14764 22928 14776
rect 22980 14764 22986 14816
rect 23290 14804 23296 14816
rect 23251 14776 23296 14804
rect 23290 14764 23296 14776
rect 23348 14764 23354 14816
rect 24228 14813 24256 14844
rect 24213 14807 24271 14813
rect 24213 14773 24225 14807
rect 24259 14804 24271 14807
rect 27614 14804 27620 14816
rect 24259 14776 27620 14804
rect 24259 14773 24271 14776
rect 24213 14767 24271 14773
rect 27614 14764 27620 14776
rect 27672 14764 27678 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2317 14603 2375 14609
rect 2317 14569 2329 14603
rect 2363 14600 2375 14603
rect 2498 14600 2504 14612
rect 2363 14572 2504 14600
rect 2363 14569 2375 14572
rect 2317 14563 2375 14569
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 3234 14560 3240 14612
rect 3292 14600 3298 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 3292 14572 5181 14600
rect 3292 14560 3298 14572
rect 5169 14569 5181 14572
rect 5215 14600 5227 14603
rect 5215 14572 5488 14600
rect 5215 14569 5227 14572
rect 5169 14563 5227 14569
rect 1949 14535 2007 14541
rect 1949 14501 1961 14535
rect 1995 14532 2007 14535
rect 5074 14532 5080 14544
rect 1995 14504 5080 14532
rect 1995 14501 2007 14504
rect 1949 14495 2007 14501
rect 2700 14473 2728 14504
rect 5074 14492 5080 14504
rect 5132 14492 5138 14544
rect 5460 14532 5488 14572
rect 5534 14560 5540 14612
rect 5592 14600 5598 14612
rect 7055 14603 7113 14609
rect 7055 14600 7067 14603
rect 5592 14572 7067 14600
rect 5592 14560 5598 14572
rect 7055 14569 7067 14572
rect 7101 14569 7113 14603
rect 9398 14600 9404 14612
rect 9359 14572 9404 14600
rect 7055 14563 7113 14569
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10045 14603 10103 14609
rect 10045 14600 10057 14603
rect 10008 14572 10057 14600
rect 10008 14560 10014 14572
rect 10045 14569 10057 14572
rect 10091 14569 10103 14603
rect 10045 14563 10103 14569
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 11422 14600 11428 14612
rect 10643 14572 11428 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 11422 14560 11428 14572
rect 11480 14600 11486 14612
rect 12897 14603 12955 14609
rect 11480 14572 11652 14600
rect 11480 14560 11486 14572
rect 5460 14504 5580 14532
rect 5552 14476 5580 14504
rect 10778 14492 10784 14544
rect 10836 14532 10842 14544
rect 11624 14541 11652 14572
rect 12897 14569 12909 14603
rect 12943 14600 12955 14603
rect 13078 14600 13084 14612
rect 12943 14572 13084 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 13630 14600 13636 14612
rect 13591 14572 13636 14600
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 14366 14600 14372 14612
rect 13780 14572 14372 14600
rect 13780 14560 13786 14572
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 14642 14600 14648 14612
rect 14603 14572 14648 14600
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 15105 14603 15163 14609
rect 15105 14569 15117 14603
rect 15151 14600 15163 14603
rect 15654 14600 15660 14612
rect 15151 14572 15660 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 18782 14600 18788 14612
rect 18743 14572 18788 14600
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 19889 14603 19947 14609
rect 19889 14569 19901 14603
rect 19935 14600 19947 14603
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 19935 14572 20453 14600
rect 19935 14569 19947 14572
rect 19889 14563 19947 14569
rect 20441 14569 20453 14572
rect 20487 14600 20499 14603
rect 20530 14600 20536 14612
rect 20487 14572 20536 14600
rect 20487 14569 20499 14572
rect 20441 14563 20499 14569
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 21910 14600 21916 14612
rect 21871 14572 21916 14600
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 10873 14535 10931 14541
rect 10873 14532 10885 14535
rect 10836 14504 10885 14532
rect 10836 14492 10842 14504
rect 10873 14501 10885 14504
rect 10919 14501 10931 14535
rect 10873 14495 10931 14501
rect 11609 14535 11667 14541
rect 11609 14501 11621 14535
rect 11655 14501 11667 14535
rect 15746 14532 15752 14544
rect 15707 14504 15752 14532
rect 11609 14495 11667 14501
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 18874 14492 18880 14544
rect 18932 14532 18938 14544
rect 19290 14535 19348 14541
rect 19290 14532 19302 14535
rect 18932 14504 19302 14532
rect 18932 14492 18938 14504
rect 19290 14501 19302 14504
rect 19336 14532 19348 14535
rect 20254 14532 20260 14544
rect 19336 14504 20260 14532
rect 19336 14501 19348 14504
rect 19290 14495 19348 14501
rect 20254 14492 20260 14504
rect 20312 14492 20318 14544
rect 21082 14532 21088 14544
rect 21043 14504 21088 14532
rect 21082 14492 21088 14504
rect 21140 14492 21146 14544
rect 22649 14535 22707 14541
rect 22649 14501 22661 14535
rect 22695 14532 22707 14535
rect 23014 14532 23020 14544
rect 22695 14504 23020 14532
rect 22695 14501 22707 14504
rect 22649 14495 22707 14501
rect 23014 14492 23020 14504
rect 23072 14492 23078 14544
rect 2409 14467 2467 14473
rect 2409 14433 2421 14467
rect 2455 14464 2467 14467
rect 2685 14467 2743 14473
rect 2455 14436 2630 14464
rect 2455 14433 2467 14436
rect 2409 14427 2467 14433
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 2498 14328 2504 14340
rect 2459 14300 2504 14328
rect 2498 14288 2504 14300
rect 2556 14288 2562 14340
rect 2602 14260 2630 14436
rect 2685 14433 2697 14467
rect 2731 14433 2743 14467
rect 2685 14427 2743 14433
rect 3694 14424 3700 14476
rect 3752 14464 3758 14476
rect 3789 14467 3847 14473
rect 3789 14464 3801 14467
rect 3752 14436 3801 14464
rect 3752 14424 3758 14436
rect 3789 14433 3801 14436
rect 3835 14433 3847 14467
rect 3789 14427 3847 14433
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4430 14464 4436 14476
rect 4111 14436 4436 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4430 14424 4436 14436
rect 4488 14464 4494 14476
rect 5350 14464 5356 14476
rect 4488 14436 5356 14464
rect 4488 14424 4494 14436
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 5534 14424 5540 14476
rect 5592 14424 5598 14476
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 5902 14464 5908 14476
rect 5675 14436 5908 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 6984 14467 7042 14473
rect 6984 14433 6996 14467
rect 7030 14464 7042 14467
rect 7190 14464 7196 14476
rect 7030 14436 7196 14464
rect 7030 14433 7042 14436
rect 6984 14427 7042 14433
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 7742 14424 7748 14476
rect 7800 14464 7806 14476
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 7800 14436 8033 14464
rect 7800 14424 7806 14436
rect 8021 14433 8033 14436
rect 8067 14433 8079 14467
rect 8478 14464 8484 14476
rect 8439 14436 8484 14464
rect 8021 14427 8079 14433
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 8846 14424 8852 14476
rect 8904 14464 8910 14476
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 8904 14436 11253 14464
rect 8904 14424 8910 14436
rect 11241 14433 11253 14436
rect 11287 14433 11299 14467
rect 17402 14464 17408 14476
rect 17363 14436 17408 14464
rect 11241 14427 11299 14433
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 17586 14424 17592 14476
rect 17644 14464 17650 14476
rect 17865 14467 17923 14473
rect 17865 14464 17877 14467
rect 17644 14436 17877 14464
rect 17644 14424 17650 14436
rect 17865 14433 17877 14436
rect 17911 14464 17923 14467
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 17911 14436 18429 14464
rect 17911 14433 17923 14436
rect 17865 14427 17923 14433
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 18506 14424 18512 14476
rect 18564 14464 18570 14476
rect 18969 14467 19027 14473
rect 18969 14464 18981 14467
rect 18564 14436 18981 14464
rect 18564 14424 18570 14436
rect 18969 14433 18981 14436
rect 19015 14464 19027 14467
rect 19886 14464 19892 14476
rect 19015 14436 19892 14464
rect 19015 14433 19027 14436
rect 18969 14427 19027 14433
rect 19886 14424 19892 14436
rect 19944 14424 19950 14476
rect 3145 14399 3203 14405
rect 3145 14365 3157 14399
rect 3191 14396 3203 14399
rect 3970 14396 3976 14408
rect 3191 14368 3976 14396
rect 3191 14365 3203 14368
rect 3145 14359 3203 14365
rect 3970 14356 3976 14368
rect 4028 14396 4034 14408
rect 5994 14396 6000 14408
rect 4028 14368 6000 14396
rect 4028 14356 4034 14368
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14396 6147 14399
rect 7834 14396 7840 14408
rect 6135 14368 7840 14396
rect 6135 14365 6147 14368
rect 6089 14359 6147 14365
rect 7834 14356 7840 14368
rect 7892 14356 7898 14408
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 9490 14396 9496 14408
rect 8803 14368 9496 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 9490 14356 9496 14368
rect 9548 14396 9554 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 9548 14368 9689 14396
rect 9548 14356 9554 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 11517 14399 11575 14405
rect 11517 14396 11529 14399
rect 11204 14368 11529 14396
rect 11204 14356 11210 14368
rect 11517 14365 11529 14368
rect 11563 14365 11575 14399
rect 11974 14396 11980 14408
rect 11935 14368 11980 14396
rect 11517 14359 11575 14365
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14396 12587 14399
rect 13170 14396 13176 14408
rect 12575 14368 13176 14396
rect 12575 14365 12587 14368
rect 12529 14359 12587 14365
rect 13170 14356 13176 14368
rect 13228 14396 13234 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13228 14368 13277 14396
rect 13228 14356 13234 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 15654 14396 15660 14408
rect 15615 14368 15660 14396
rect 13265 14359 13323 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14396 16359 14399
rect 16482 14396 16488 14408
rect 16347 14368 16488 14396
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14396 18199 14399
rect 20438 14396 20444 14408
rect 18187 14368 20444 14396
rect 18187 14365 18199 14368
rect 18141 14359 18199 14365
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 20990 14396 20996 14408
rect 20951 14368 20996 14396
rect 20990 14356 20996 14368
rect 21048 14356 21054 14408
rect 21266 14396 21272 14408
rect 21227 14368 21272 14396
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 22557 14399 22615 14405
rect 22557 14396 22569 14399
rect 22152 14368 22569 14396
rect 22152 14356 22158 14368
rect 22557 14365 22569 14368
rect 22603 14365 22615 14399
rect 22830 14396 22836 14408
rect 22791 14368 22836 14396
rect 22557 14359 22615 14365
rect 22830 14356 22836 14368
rect 22888 14356 22894 14408
rect 3510 14328 3516 14340
rect 3471 14300 3516 14328
rect 3510 14288 3516 14300
rect 3568 14288 3574 14340
rect 5442 14288 5448 14340
rect 5500 14328 5506 14340
rect 6457 14331 6515 14337
rect 6457 14328 6469 14331
rect 5500 14300 6469 14328
rect 5500 14288 5506 14300
rect 6457 14297 6469 14300
rect 6503 14328 6515 14331
rect 6546 14328 6552 14340
rect 6503 14300 6552 14328
rect 6503 14297 6515 14300
rect 6457 14291 6515 14297
rect 6546 14288 6552 14300
rect 6604 14288 6610 14340
rect 20162 14288 20168 14340
rect 20220 14328 20226 14340
rect 21008 14328 21036 14356
rect 20220 14300 21036 14328
rect 20220 14288 20226 14300
rect 3602 14260 3608 14272
rect 2602 14232 3608 14260
rect 3602 14220 3608 14232
rect 3660 14260 3666 14272
rect 4065 14263 4123 14269
rect 4065 14260 4077 14263
rect 3660 14232 4077 14260
rect 3660 14220 3666 14232
rect 4065 14229 4077 14232
rect 4111 14229 4123 14263
rect 4246 14260 4252 14272
rect 4207 14232 4252 14260
rect 4065 14223 4123 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 4893 14263 4951 14269
rect 4893 14229 4905 14263
rect 4939 14260 4951 14263
rect 5350 14260 5356 14272
rect 4939 14232 5356 14260
rect 4939 14229 4951 14232
rect 4893 14223 4951 14229
rect 5350 14220 5356 14232
rect 5408 14260 5414 14272
rect 7006 14260 7012 14272
rect 5408 14232 7012 14260
rect 5408 14220 5414 14232
rect 7006 14220 7012 14232
rect 7064 14260 7070 14272
rect 7377 14263 7435 14269
rect 7377 14260 7389 14263
rect 7064 14232 7389 14260
rect 7064 14220 7070 14232
rect 7377 14229 7389 14232
rect 7423 14229 7435 14263
rect 9030 14260 9036 14272
rect 8991 14232 9036 14260
rect 7377 14223 7435 14229
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 14185 14263 14243 14269
rect 14185 14229 14197 14263
rect 14231 14260 14243 14263
rect 14366 14260 14372 14272
rect 14231 14232 14372 14260
rect 14231 14229 14243 14232
rect 14185 14223 14243 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 16298 14220 16304 14272
rect 16356 14260 16362 14272
rect 16577 14263 16635 14269
rect 16577 14260 16589 14263
rect 16356 14232 16589 14260
rect 16356 14220 16362 14232
rect 16577 14229 16589 14232
rect 16623 14229 16635 14263
rect 16577 14223 16635 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 8021 14059 8079 14065
rect 8021 14056 8033 14059
rect 7800 14028 8033 14056
rect 7800 14016 7806 14028
rect 8021 14025 8033 14028
rect 8067 14025 8079 14059
rect 9582 14056 9588 14068
rect 9543 14028 9588 14056
rect 8021 14019 8079 14025
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 11422 14056 11428 14068
rect 11383 14028 11428 14056
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 12342 14056 12348 14068
rect 12299 14028 12348 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12526 14056 12532 14068
rect 12487 14028 12532 14056
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 13354 14016 13360 14068
rect 13412 14016 13418 14068
rect 13630 14016 13636 14068
rect 13688 14056 13694 14068
rect 13725 14059 13783 14065
rect 13725 14056 13737 14059
rect 13688 14028 13737 14056
rect 13688 14016 13694 14028
rect 13725 14025 13737 14028
rect 13771 14025 13783 14059
rect 13725 14019 13783 14025
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 14424 14028 14473 14056
rect 14424 14016 14430 14028
rect 14461 14025 14473 14028
rect 14507 14056 14519 14059
rect 15746 14056 15752 14068
rect 14507 14028 15752 14056
rect 14507 14025 14519 14028
rect 14461 14019 14519 14025
rect 15746 14016 15752 14028
rect 15804 14056 15810 14068
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15804 14028 15945 14056
rect 15804 14016 15810 14028
rect 15933 14025 15945 14028
rect 15979 14025 15991 14059
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 15933 14019 15991 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 17586 14016 17592 14068
rect 17644 14056 17650 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17644 14028 17785 14056
rect 17644 14016 17650 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 19613 14059 19671 14065
rect 19613 14025 19625 14059
rect 19659 14056 19671 14059
rect 21082 14056 21088 14068
rect 19659 14028 21088 14056
rect 19659 14025 19671 14028
rect 19613 14019 19671 14025
rect 21082 14016 21088 14028
rect 21140 14056 21146 14068
rect 21637 14059 21695 14065
rect 21637 14056 21649 14059
rect 21140 14028 21649 14056
rect 21140 14016 21146 14028
rect 21637 14025 21649 14028
rect 21683 14025 21695 14059
rect 22738 14056 22744 14068
rect 22699 14028 22744 14056
rect 21637 14019 21695 14025
rect 22738 14016 22744 14028
rect 22796 14016 22802 14068
rect 23014 14056 23020 14068
rect 22975 14028 23020 14056
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 2133 13991 2191 13997
rect 2133 13957 2145 13991
rect 2179 13988 2191 13991
rect 3510 13988 3516 14000
rect 2179 13960 3516 13988
rect 2179 13957 2191 13960
rect 2133 13951 2191 13957
rect 3510 13948 3516 13960
rect 3568 13948 3574 14000
rect 5166 13988 5172 14000
rect 4172 13960 5172 13988
rect 2866 13880 2872 13932
rect 2924 13920 2930 13932
rect 3786 13920 3792 13932
rect 2924 13892 3792 13920
rect 2924 13880 2930 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1670 13852 1676 13864
rect 1443 13824 1676 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 3160 13861 3188 13892
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13821 3203 13855
rect 3145 13815 3203 13821
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13821 3663 13855
rect 3605 13815 3663 13821
rect 1486 13744 1492 13796
rect 1544 13784 1550 13796
rect 2409 13787 2467 13793
rect 2409 13784 2421 13787
rect 1544 13756 2421 13784
rect 1544 13744 1550 13756
rect 2409 13753 2421 13756
rect 2455 13784 2467 13787
rect 2498 13784 2504 13796
rect 2455 13756 2504 13784
rect 2455 13753 2467 13756
rect 2409 13747 2467 13753
rect 2498 13744 2504 13756
rect 2556 13784 2562 13796
rect 2556 13756 3188 13784
rect 2556 13744 2562 13756
rect 1118 13676 1124 13728
rect 1176 13716 1182 13728
rect 1581 13719 1639 13725
rect 1581 13716 1593 13719
rect 1176 13688 1593 13716
rect 1176 13676 1182 13688
rect 1581 13685 1593 13688
rect 1627 13685 1639 13719
rect 2958 13716 2964 13728
rect 2919 13688 2964 13716
rect 1581 13679 1639 13685
rect 2958 13676 2964 13688
rect 3016 13676 3022 13728
rect 3160 13716 3188 13756
rect 3510 13744 3516 13796
rect 3568 13784 3574 13796
rect 3620 13784 3648 13815
rect 3694 13812 3700 13864
rect 3752 13852 3758 13864
rect 3752 13824 3797 13852
rect 3752 13812 3758 13824
rect 4172 13784 4200 13960
rect 5166 13948 5172 13960
rect 5224 13988 5230 14000
rect 5261 13991 5319 13997
rect 5261 13988 5273 13991
rect 5224 13960 5273 13988
rect 5224 13948 5230 13960
rect 5261 13957 5273 13960
rect 5307 13957 5319 13991
rect 10778 13988 10784 14000
rect 5261 13951 5319 13957
rect 10244 13960 10784 13988
rect 4982 13880 4988 13932
rect 5040 13920 5046 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5040 13892 5641 13920
rect 5040 13880 5046 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13920 7159 13923
rect 7466 13920 7472 13932
rect 7147 13892 7472 13920
rect 7147 13889 7159 13892
rect 7101 13883 7159 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13920 7803 13923
rect 8478 13920 8484 13932
rect 7791 13892 8484 13920
rect 7791 13889 7803 13892
rect 7745 13883 7803 13889
rect 8478 13880 8484 13892
rect 8536 13880 8542 13932
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13920 8723 13923
rect 9030 13920 9036 13932
rect 8711 13892 9036 13920
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 5169 13855 5227 13861
rect 4295 13824 4476 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 4448 13796 4476 13824
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5350 13852 5356 13864
rect 5215 13824 5356 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13852 5503 13855
rect 5534 13852 5540 13864
rect 5491 13824 5540 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 7006 13852 7012 13864
rect 6967 13824 7012 13852
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7282 13852 7288 13864
rect 7243 13824 7288 13852
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 3568 13756 4200 13784
rect 3568 13744 3574 13756
rect 4430 13744 4436 13796
rect 4488 13784 4494 13796
rect 4617 13787 4675 13793
rect 4617 13784 4629 13787
rect 4488 13756 4629 13784
rect 4488 13744 4494 13756
rect 4617 13753 4629 13756
rect 4663 13753 4675 13787
rect 4617 13747 4675 13753
rect 8294 13744 8300 13796
rect 8352 13784 8358 13796
rect 8573 13787 8631 13793
rect 8573 13784 8585 13787
rect 8352 13756 8585 13784
rect 8352 13744 8358 13756
rect 8573 13753 8585 13756
rect 8619 13784 8631 13787
rect 9027 13787 9085 13793
rect 9027 13784 9039 13787
rect 8619 13756 9039 13784
rect 8619 13753 8631 13756
rect 8573 13747 8631 13753
rect 9027 13753 9039 13756
rect 9073 13784 9085 13787
rect 10244 13784 10272 13960
rect 10778 13948 10784 13960
rect 10836 13948 10842 14000
rect 12544 13988 12572 14016
rect 13372 13988 13400 14016
rect 14001 13991 14059 13997
rect 14001 13988 14013 13991
rect 12544 13960 14013 13988
rect 14001 13957 14013 13960
rect 14047 13957 14059 13991
rect 14001 13951 14059 13957
rect 15657 13991 15715 13997
rect 15657 13957 15669 13991
rect 15703 13988 15715 13991
rect 15838 13988 15844 14000
rect 15703 13960 15844 13988
rect 15703 13957 15715 13960
rect 15657 13951 15715 13957
rect 15838 13948 15844 13960
rect 15896 13948 15902 14000
rect 19886 13988 19892 14000
rect 19847 13960 19892 13988
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 20254 13988 20260 14000
rect 20215 13960 20260 13988
rect 20254 13948 20260 13960
rect 20312 13948 20318 14000
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13920 10379 13923
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 10367 13892 10517 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 10505 13889 10517 13892
rect 10551 13920 10563 13923
rect 10686 13920 10692 13932
rect 10551 13892 10692 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 11146 13920 11152 13932
rect 11107 13892 11152 13920
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 13357 13923 13415 13929
rect 12584 13892 12940 13920
rect 12584 13880 12590 13892
rect 12912 13861 12940 13892
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 14734 13920 14740 13932
rect 13403 13892 14740 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 16206 13920 16212 13932
rect 15335 13892 16212 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 15856 13864 15884 13892
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 16482 13920 16488 13932
rect 16443 13892 16488 13920
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 18693 13923 18751 13929
rect 18693 13889 18705 13923
rect 18739 13920 18751 13923
rect 18782 13920 18788 13932
rect 18739 13892 18788 13920
rect 18739 13889 18751 13892
rect 18693 13883 18751 13889
rect 18782 13880 18788 13892
rect 18840 13880 18846 13932
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13821 12771 13855
rect 12713 13815 12771 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 10597 13787 10655 13793
rect 10597 13784 10609 13787
rect 9073 13756 9996 13784
rect 10244 13756 10609 13784
rect 9073 13753 9085 13756
rect 9027 13747 9085 13753
rect 9968 13728 9996 13756
rect 10597 13753 10609 13756
rect 10643 13753 10655 13787
rect 10597 13747 10655 13753
rect 4985 13719 5043 13725
rect 4985 13716 4997 13719
rect 3160 13688 4997 13716
rect 4985 13685 4997 13688
rect 5031 13716 5043 13719
rect 5442 13716 5448 13728
rect 5031 13688 5448 13716
rect 5031 13685 5043 13688
rect 4985 13679 5043 13685
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 6181 13719 6239 13725
rect 6181 13716 6193 13719
rect 6052 13688 6193 13716
rect 6052 13676 6058 13688
rect 6181 13685 6193 13688
rect 6227 13685 6239 13719
rect 6181 13679 6239 13685
rect 6641 13719 6699 13725
rect 6641 13685 6653 13719
rect 6687 13716 6699 13719
rect 7190 13716 7196 13728
rect 6687 13688 7196 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 9950 13716 9956 13728
rect 9911 13688 9956 13716
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 11885 13719 11943 13725
rect 11885 13685 11897 13719
rect 11931 13716 11943 13719
rect 12618 13716 12624 13728
rect 11931 13688 12624 13716
rect 11931 13685 11943 13688
rect 11885 13679 11943 13685
rect 12618 13676 12624 13688
rect 12676 13716 12682 13728
rect 12728 13716 12756 13815
rect 15838 13812 15844 13864
rect 15896 13812 15902 13864
rect 14642 13784 14648 13796
rect 14603 13756 14648 13784
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 14737 13787 14795 13793
rect 14737 13753 14749 13787
rect 14783 13753 14795 13787
rect 16206 13784 16212 13796
rect 16167 13756 16212 13784
rect 14737 13747 14795 13753
rect 12676 13688 12756 13716
rect 12676 13676 12682 13688
rect 14366 13676 14372 13728
rect 14424 13716 14430 13728
rect 14752 13716 14780 13747
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 16301 13787 16359 13793
rect 16301 13753 16313 13787
rect 16347 13784 16359 13787
rect 16390 13784 16396 13796
rect 16347 13756 16396 13784
rect 16347 13753 16359 13756
rect 16301 13747 16359 13753
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 19014 13787 19072 13793
rect 19014 13753 19026 13787
rect 19060 13753 19072 13787
rect 19014 13747 19072 13753
rect 14424 13688 14780 13716
rect 14424 13676 14430 13688
rect 18414 13676 18420 13728
rect 18472 13716 18478 13728
rect 18509 13719 18567 13725
rect 18509 13716 18521 13719
rect 18472 13688 18521 13716
rect 18472 13676 18478 13688
rect 18509 13685 18521 13688
rect 18555 13716 18567 13719
rect 18874 13716 18880 13728
rect 18555 13688 18880 13716
rect 18555 13685 18567 13688
rect 18509 13679 18567 13685
rect 18874 13676 18880 13688
rect 18932 13716 18938 13728
rect 19029 13716 19057 13747
rect 18932 13688 19057 13716
rect 20272 13716 20300 13948
rect 20438 13920 20444 13932
rect 20399 13892 20444 13920
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 22256 13855 22314 13861
rect 22256 13821 22268 13855
rect 22302 13852 22314 13855
rect 22738 13852 22744 13864
rect 22302 13824 22744 13852
rect 22302 13821 22314 13824
rect 22256 13815 22314 13821
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 23382 13812 23388 13864
rect 23440 13852 23446 13864
rect 23712 13855 23770 13861
rect 23712 13852 23724 13855
rect 23440 13824 23724 13852
rect 23440 13812 23446 13824
rect 23712 13821 23724 13824
rect 23758 13852 23770 13855
rect 24121 13855 24179 13861
rect 24121 13852 24133 13855
rect 23758 13824 24133 13852
rect 23758 13821 23770 13824
rect 23712 13815 23770 13821
rect 24121 13821 24133 13824
rect 24167 13821 24179 13855
rect 24121 13815 24179 13821
rect 20530 13744 20536 13796
rect 20588 13784 20594 13796
rect 23799 13787 23857 13793
rect 23799 13784 23811 13787
rect 20588 13756 23811 13784
rect 20588 13744 20594 13756
rect 23799 13753 23811 13756
rect 23845 13753 23857 13787
rect 23799 13747 23857 13753
rect 20809 13719 20867 13725
rect 20809 13716 20821 13719
rect 20272 13688 20821 13716
rect 18932 13676 18938 13688
rect 20809 13685 20821 13688
rect 20855 13685 20867 13719
rect 21358 13716 21364 13728
rect 21319 13688 21364 13716
rect 20809 13679 20867 13685
rect 21358 13676 21364 13688
rect 21416 13676 21422 13728
rect 22094 13716 22100 13728
rect 22055 13688 22100 13716
rect 22094 13676 22100 13688
rect 22152 13676 22158 13728
rect 22186 13676 22192 13728
rect 22244 13716 22250 13728
rect 22327 13719 22385 13725
rect 22327 13716 22339 13719
rect 22244 13688 22339 13716
rect 22244 13676 22250 13688
rect 22327 13685 22339 13688
rect 22373 13685 22385 13719
rect 22327 13679 22385 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1670 13512 1676 13524
rect 1583 13484 1676 13512
rect 1670 13472 1676 13484
rect 1728 13512 1734 13524
rect 9490 13512 9496 13524
rect 1728 13484 9352 13512
rect 9451 13484 9496 13512
rect 1728 13472 1734 13484
rect 2587 13447 2645 13453
rect 2587 13413 2599 13447
rect 2633 13444 2645 13447
rect 2774 13444 2780 13456
rect 2633 13416 2780 13444
rect 2633 13413 2645 13416
rect 2587 13407 2645 13413
rect 2774 13404 2780 13416
rect 2832 13404 2838 13456
rect 4246 13444 4252 13456
rect 3160 13416 4252 13444
rect 2682 13336 2688 13388
rect 2740 13376 2746 13388
rect 3160 13385 3188 13416
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 5442 13404 5448 13456
rect 5500 13444 5506 13456
rect 9324 13444 9352 13484
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 13170 13512 13176 13524
rect 10612 13484 13032 13512
rect 13131 13484 13176 13512
rect 10612 13444 10640 13484
rect 5500 13416 5764 13444
rect 9324 13416 10640 13444
rect 10689 13447 10747 13453
rect 5500 13404 5506 13416
rect 5736 13385 5764 13416
rect 10689 13413 10701 13447
rect 10735 13444 10747 13447
rect 11701 13447 11759 13453
rect 11701 13444 11713 13447
rect 10735 13416 11713 13444
rect 10735 13413 10747 13416
rect 10689 13407 10747 13413
rect 11701 13413 11713 13416
rect 11747 13444 11759 13447
rect 11790 13444 11796 13456
rect 11747 13416 11796 13444
rect 11747 13413 11759 13416
rect 11701 13407 11759 13413
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 12618 13404 12624 13456
rect 12676 13444 12682 13456
rect 12805 13447 12863 13453
rect 12805 13444 12817 13447
rect 12676 13416 12817 13444
rect 12676 13404 12682 13416
rect 12805 13413 12817 13416
rect 12851 13413 12863 13447
rect 13004 13444 13032 13484
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 15105 13515 15163 13521
rect 15105 13481 15117 13515
rect 15151 13512 15163 13515
rect 15562 13512 15568 13524
rect 15151 13484 15568 13512
rect 15151 13481 15163 13484
rect 15105 13475 15163 13481
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 16022 13512 16028 13524
rect 15672 13484 16028 13512
rect 13446 13444 13452 13456
rect 13004 13416 13452 13444
rect 12805 13407 12863 13413
rect 13446 13404 13452 13416
rect 13504 13404 13510 13456
rect 15672 13453 15700 13484
rect 16022 13472 16028 13484
rect 16080 13512 16086 13524
rect 16390 13512 16396 13524
rect 16080 13484 16396 13512
rect 16080 13472 16086 13484
rect 16390 13472 16396 13484
rect 16448 13512 16454 13524
rect 16485 13515 16543 13521
rect 16485 13512 16497 13515
rect 16448 13484 16497 13512
rect 16448 13472 16454 13484
rect 16485 13481 16497 13484
rect 16531 13481 16543 13515
rect 16485 13475 16543 13481
rect 18414 13472 18420 13524
rect 18472 13512 18478 13524
rect 18509 13515 18567 13521
rect 18509 13512 18521 13515
rect 18472 13484 18521 13512
rect 18472 13472 18478 13484
rect 18509 13481 18521 13484
rect 18555 13512 18567 13515
rect 19337 13515 19395 13521
rect 19337 13512 19349 13515
rect 18555 13484 19349 13512
rect 18555 13481 18567 13484
rect 18509 13475 18567 13481
rect 19337 13481 19349 13484
rect 19383 13481 19395 13515
rect 20162 13512 20168 13524
rect 20123 13484 20168 13512
rect 19337 13475 19395 13481
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 20438 13512 20444 13524
rect 20399 13484 20444 13512
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 22094 13472 22100 13524
rect 22152 13512 22158 13524
rect 24167 13515 24225 13521
rect 24167 13512 24179 13515
rect 22152 13484 24179 13512
rect 22152 13472 22158 13484
rect 24167 13481 24179 13484
rect 24213 13481 24225 13515
rect 24167 13475 24225 13481
rect 15657 13447 15715 13453
rect 15657 13413 15669 13447
rect 15703 13413 15715 13447
rect 15657 13407 15715 13413
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 19797 13447 19855 13453
rect 19797 13444 19809 13447
rect 19484 13416 19809 13444
rect 19484 13404 19490 13416
rect 19797 13413 19809 13416
rect 19843 13444 19855 13447
rect 20530 13444 20536 13456
rect 19843 13416 20536 13444
rect 19843 13413 19855 13416
rect 19797 13407 19855 13413
rect 20530 13404 20536 13416
rect 20588 13404 20594 13456
rect 20714 13404 20720 13456
rect 20772 13444 20778 13456
rect 21085 13447 21143 13453
rect 21085 13444 21097 13447
rect 20772 13416 21097 13444
rect 20772 13404 20778 13416
rect 21085 13413 21097 13416
rect 21131 13444 21143 13447
rect 21358 13444 21364 13456
rect 21131 13416 21364 13444
rect 21131 13413 21143 13416
rect 21085 13407 21143 13413
rect 21358 13404 21364 13416
rect 21416 13404 21422 13456
rect 22646 13444 22652 13456
rect 22607 13416 22652 13444
rect 22646 13404 22652 13416
rect 22704 13404 22710 13456
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 2740 13348 3157 13376
rect 2740 13336 2746 13348
rect 3145 13345 3157 13348
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 5629 13379 5687 13385
rect 5629 13345 5641 13379
rect 5675 13345 5687 13379
rect 5629 13339 5687 13345
rect 5721 13379 5779 13385
rect 5721 13345 5733 13379
rect 5767 13345 5779 13379
rect 5721 13339 5779 13345
rect 5905 13379 5963 13385
rect 5905 13345 5917 13379
rect 5951 13376 5963 13379
rect 5994 13376 6000 13388
rect 5951 13348 6000 13376
rect 5951 13345 5963 13348
rect 5905 13339 5963 13345
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13308 2283 13311
rect 3510 13308 3516 13320
rect 2271 13280 3516 13308
rect 2271 13277 2283 13280
rect 2225 13271 2283 13277
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 4212 13280 4257 13308
rect 4212 13268 4218 13280
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 4433 13311 4491 13317
rect 4433 13308 4445 13311
rect 4396 13280 4445 13308
rect 4396 13268 4402 13280
rect 4433 13277 4445 13280
rect 4479 13277 4491 13311
rect 5644 13308 5672 13339
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 7834 13376 7840 13388
rect 7795 13348 7840 13376
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13376 8355 13379
rect 8478 13376 8484 13388
rect 8343 13348 8484 13376
rect 8343 13345 8355 13348
rect 8297 13339 8355 13345
rect 8478 13336 8484 13348
rect 8536 13376 8542 13388
rect 8849 13379 8907 13385
rect 8849 13376 8861 13379
rect 8536 13348 8861 13376
rect 8536 13336 8542 13348
rect 8849 13345 8861 13348
rect 8895 13345 8907 13379
rect 10134 13376 10140 13388
rect 10095 13348 10140 13376
rect 8849 13339 8907 13345
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 13262 13376 13268 13388
rect 13223 13348 13268 13376
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13630 13376 13636 13388
rect 13543 13348 13636 13376
rect 13630 13336 13636 13348
rect 13688 13376 13694 13388
rect 14001 13379 14059 13385
rect 14001 13376 14013 13379
rect 13688 13348 14013 13376
rect 13688 13336 13694 13348
rect 14001 13345 14013 13348
rect 14047 13345 14059 13379
rect 15378 13376 15384 13388
rect 14001 13339 14059 13345
rect 15028 13348 15384 13376
rect 6086 13308 6092 13320
rect 5644 13280 6092 13308
rect 4433 13271 4491 13277
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 6328 13280 6377 13308
rect 6328 13268 6334 13280
rect 6365 13277 6377 13280
rect 6411 13308 6423 13311
rect 7374 13308 7380 13320
rect 6411 13280 7380 13308
rect 6411 13277 6423 13280
rect 6365 13271 6423 13277
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 8386 13308 8392 13320
rect 8347 13280 8392 13308
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 11882 13308 11888 13320
rect 11843 13280 11888 13308
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 13280 13308 13308 13336
rect 14366 13308 14372 13320
rect 13280 13280 14372 13308
rect 14366 13268 14372 13280
rect 14424 13308 14430 13320
rect 15028 13308 15056 13348
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 17034 13376 17040 13388
rect 16995 13348 17040 13376
rect 17034 13336 17040 13348
rect 17092 13336 17098 13388
rect 24096 13379 24154 13385
rect 24096 13345 24108 13379
rect 24142 13376 24154 13379
rect 24210 13376 24216 13388
rect 24142 13348 24216 13376
rect 24142 13345 24154 13348
rect 24096 13339 24154 13345
rect 24210 13336 24216 13348
rect 24268 13336 24274 13388
rect 15562 13308 15568 13320
rect 14424 13280 15056 13308
rect 15523 13280 15568 13308
rect 14424 13268 14430 13280
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 15838 13308 15844 13320
rect 15799 13280 15844 13308
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 17862 13268 17868 13320
rect 17920 13308 17926 13320
rect 18141 13311 18199 13317
rect 18141 13308 18153 13311
rect 17920 13280 18153 13308
rect 17920 13268 17926 13280
rect 18141 13277 18153 13280
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13308 21051 13311
rect 21450 13308 21456 13320
rect 21039 13280 21456 13308
rect 21039 13277 21051 13280
rect 20993 13271 21051 13277
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 22554 13308 22560 13320
rect 22515 13280 22560 13308
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 22830 13308 22836 13320
rect 22791 13280 22836 13308
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 7009 13243 7067 13249
rect 7009 13240 7021 13243
rect 4126 13212 7021 13240
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 3326 13172 3332 13184
rect 2179 13144 3332 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 3326 13132 3332 13144
rect 3384 13172 3390 13184
rect 3421 13175 3479 13181
rect 3421 13172 3433 13175
rect 3384 13144 3433 13172
rect 3384 13132 3390 13144
rect 3421 13141 3433 13144
rect 3467 13141 3479 13175
rect 3421 13135 3479 13141
rect 3786 13132 3792 13184
rect 3844 13172 3850 13184
rect 3881 13175 3939 13181
rect 3881 13172 3893 13175
rect 3844 13144 3893 13172
rect 3844 13132 3850 13144
rect 3881 13141 3893 13144
rect 3927 13172 3939 13175
rect 3970 13172 3976 13184
rect 3927 13144 3976 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 3970 13132 3976 13144
rect 4028 13172 4034 13184
rect 4126 13172 4154 13212
rect 7009 13209 7021 13212
rect 7055 13240 7067 13243
rect 7282 13240 7288 13252
rect 7055 13212 7288 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 11900 13240 11928 13268
rect 14458 13240 14464 13252
rect 11900 13212 14464 13240
rect 14458 13200 14464 13212
rect 14516 13200 14522 13252
rect 14642 13240 14648 13252
rect 14555 13212 14648 13240
rect 14642 13200 14648 13212
rect 14700 13240 14706 13252
rect 17175 13243 17233 13249
rect 17175 13240 17187 13243
rect 14700 13212 17187 13240
rect 14700 13200 14706 13212
rect 17175 13209 17187 13212
rect 17221 13209 17233 13243
rect 17175 13203 17233 13209
rect 21266 13200 21272 13252
rect 21324 13240 21330 13252
rect 21545 13243 21603 13249
rect 21545 13240 21557 13243
rect 21324 13212 21557 13240
rect 21324 13200 21330 13212
rect 21545 13209 21557 13212
rect 21591 13240 21603 13243
rect 23934 13240 23940 13252
rect 21591 13212 23940 13240
rect 21591 13209 21603 13212
rect 21545 13203 21603 13209
rect 23934 13200 23940 13212
rect 23992 13200 23998 13252
rect 5166 13172 5172 13184
rect 4028 13144 4154 13172
rect 5127 13144 5172 13172
rect 4028 13132 4034 13144
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 6730 13172 6736 13184
rect 6691 13144 6736 13172
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 7098 13132 7104 13184
rect 7156 13172 7162 13184
rect 7377 13175 7435 13181
rect 7377 13172 7389 13175
rect 7156 13144 7389 13172
rect 7156 13132 7162 13144
rect 7377 13141 7389 13144
rect 7423 13172 7435 13175
rect 7466 13172 7472 13184
rect 7423 13144 7472 13172
rect 7423 13141 7435 13144
rect 7377 13135 7435 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 10870 13132 10876 13184
rect 10928 13172 10934 13184
rect 10965 13175 11023 13181
rect 10965 13172 10977 13175
rect 10928 13144 10977 13172
rect 10928 13132 10934 13144
rect 10965 13141 10977 13144
rect 11011 13141 11023 13175
rect 10965 13135 11023 13141
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 11333 13175 11391 13181
rect 11333 13172 11345 13175
rect 11296 13144 11345 13172
rect 11296 13132 11302 13144
rect 11333 13141 11345 13144
rect 11379 13141 11391 13175
rect 12618 13172 12624 13184
rect 12579 13144 12624 13172
rect 11333 13135 11391 13141
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 12805 13175 12863 13181
rect 12805 13141 12817 13175
rect 12851 13172 12863 13175
rect 12989 13175 13047 13181
rect 12989 13172 13001 13175
rect 12851 13144 13001 13172
rect 12851 13141 12863 13144
rect 12805 13135 12863 13141
rect 12989 13141 13001 13144
rect 13035 13172 13047 13175
rect 13170 13172 13176 13184
rect 13035 13144 13176 13172
rect 13035 13141 13047 13144
rect 12989 13135 13047 13141
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 14001 13175 14059 13181
rect 14001 13141 14013 13175
rect 14047 13172 14059 13175
rect 14185 13175 14243 13181
rect 14185 13172 14197 13175
rect 14047 13144 14197 13172
rect 14047 13141 14059 13144
rect 14001 13135 14059 13141
rect 14185 13141 14197 13144
rect 14231 13172 14243 13175
rect 17494 13172 17500 13184
rect 14231 13144 17500 13172
rect 14231 13141 14243 13144
rect 14185 13135 14243 13141
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 19058 13172 19064 13184
rect 19019 13144 19064 13172
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 3145 12971 3203 12977
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 3234 12968 3240 12980
rect 3191 12940 3240 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 5442 12968 5448 12980
rect 5403 12940 5448 12968
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 7834 12968 7840 12980
rect 7795 12940 7840 12968
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 14366 12968 14372 12980
rect 14327 12940 14372 12968
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 16666 12977 16672 12980
rect 16623 12971 16672 12977
rect 16623 12968 16635 12971
rect 15620 12940 16635 12968
rect 15620 12928 15626 12940
rect 16623 12937 16635 12940
rect 16669 12937 16672 12971
rect 16623 12931 16672 12937
rect 16666 12928 16672 12931
rect 16724 12928 16730 12980
rect 20714 12968 20720 12980
rect 20675 12940 20720 12968
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 21085 12971 21143 12977
rect 21085 12937 21097 12971
rect 21131 12968 21143 12971
rect 21358 12968 21364 12980
rect 21131 12940 21364 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 21358 12928 21364 12940
rect 21416 12968 21422 12980
rect 22557 12971 22615 12977
rect 22557 12968 22569 12971
rect 21416 12940 22569 12968
rect 21416 12928 21422 12940
rect 22557 12937 22569 12940
rect 22603 12968 22615 12971
rect 22646 12968 22652 12980
rect 22603 12940 22652 12968
rect 22603 12937 22615 12940
rect 22557 12931 22615 12937
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 24121 12971 24179 12977
rect 24121 12937 24133 12971
rect 24167 12968 24179 12971
rect 24210 12968 24216 12980
rect 24167 12940 24216 12968
rect 24167 12937 24179 12940
rect 24121 12931 24179 12937
rect 24210 12928 24216 12940
rect 24268 12928 24274 12980
rect 24765 12971 24823 12977
rect 24765 12937 24777 12971
rect 24811 12968 24823 12971
rect 24946 12968 24952 12980
rect 24811 12940 24952 12968
rect 24811 12937 24823 12940
rect 24765 12931 24823 12937
rect 24946 12928 24952 12940
rect 25004 12928 25010 12980
rect 2774 12900 2780 12912
rect 2687 12872 2780 12900
rect 2774 12860 2780 12872
rect 2832 12900 2838 12912
rect 5534 12900 5540 12912
rect 2832 12872 5540 12900
rect 2832 12860 2838 12872
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 6822 12860 6828 12912
rect 6880 12900 6886 12912
rect 6880 12872 7236 12900
rect 6880 12860 6886 12872
rect 1394 12792 1400 12844
rect 1452 12832 1458 12844
rect 1765 12835 1823 12841
rect 1765 12832 1777 12835
rect 1452 12804 1777 12832
rect 1452 12792 1458 12804
rect 1765 12801 1777 12804
rect 1811 12801 1823 12835
rect 2406 12832 2412 12844
rect 2367 12804 2412 12832
rect 1765 12795 1823 12801
rect 2406 12792 2412 12804
rect 2464 12832 2470 12844
rect 4338 12832 4344 12844
rect 2464 12804 4344 12832
rect 2464 12792 2470 12804
rect 4338 12792 4344 12804
rect 4396 12792 4402 12844
rect 5767 12835 5825 12841
rect 5767 12801 5779 12835
rect 5813 12832 5825 12835
rect 6730 12832 6736 12844
rect 5813 12804 6736 12832
rect 5813 12801 5825 12804
rect 5767 12795 5825 12801
rect 6730 12792 6736 12804
rect 6788 12832 6794 12844
rect 7208 12841 7236 12872
rect 7374 12860 7380 12912
rect 7432 12900 7438 12912
rect 8297 12903 8355 12909
rect 8297 12900 8309 12903
rect 7432 12872 8309 12900
rect 7432 12860 7438 12872
rect 8297 12869 8309 12872
rect 8343 12900 8355 12903
rect 13630 12900 13636 12912
rect 8343 12872 13636 12900
rect 8343 12869 8355 12872
rect 8297 12863 8355 12869
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 6788 12804 6929 12832
rect 6788 12792 6794 12804
rect 6917 12801 6929 12804
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 3234 12764 3240 12776
rect 3195 12736 3240 12764
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3694 12764 3700 12776
rect 3655 12736 3700 12764
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 4246 12764 4252 12776
rect 4207 12736 4252 12764
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 4430 12764 4436 12776
rect 4391 12736 4436 12764
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12764 5227 12767
rect 5680 12767 5738 12773
rect 5680 12764 5692 12767
rect 5215 12736 5692 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 5680 12733 5692 12736
rect 5726 12764 5738 12767
rect 6178 12764 6184 12776
rect 5726 12736 6184 12764
rect 5726 12733 5738 12736
rect 5680 12727 5738 12733
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 8404 12773 8432 12872
rect 13630 12860 13636 12872
rect 13688 12860 13694 12912
rect 16022 12900 16028 12912
rect 13786 12872 15792 12900
rect 15983 12872 16028 12900
rect 9030 12832 9036 12844
rect 8991 12804 9036 12832
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 11882 12832 11888 12844
rect 11563 12804 11888 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 13786 12832 13814 12872
rect 12032 12804 13814 12832
rect 12032 12792 12038 12804
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 15289 12835 15347 12841
rect 15289 12832 15301 12835
rect 14884 12804 15301 12832
rect 14884 12792 14890 12804
rect 15289 12801 15301 12804
rect 15335 12832 15347 12835
rect 15654 12832 15660 12844
rect 15335 12804 15660 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 8389 12767 8447 12773
rect 8389 12733 8401 12767
rect 8435 12733 8447 12767
rect 8389 12727 8447 12733
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 8849 12767 8907 12773
rect 8849 12764 8861 12767
rect 8536 12736 8861 12764
rect 8536 12724 8542 12736
rect 8849 12733 8861 12736
rect 8895 12733 8907 12767
rect 8849 12727 8907 12733
rect 12529 12767 12587 12773
rect 12529 12733 12541 12767
rect 12575 12733 12587 12767
rect 13170 12764 13176 12776
rect 13131 12736 13176 12764
rect 12529 12727 12587 12733
rect 1854 12656 1860 12708
rect 1912 12696 1918 12708
rect 1912 12668 1957 12696
rect 1912 12656 1918 12668
rect 4706 12656 4712 12708
rect 4764 12696 4770 12708
rect 5994 12696 6000 12708
rect 4764 12668 6000 12696
rect 4764 12656 4770 12668
rect 5994 12656 6000 12668
rect 6052 12696 6058 12708
rect 6457 12699 6515 12705
rect 6457 12696 6469 12699
rect 6052 12668 6469 12696
rect 6052 12656 6058 12668
rect 6457 12665 6469 12668
rect 6503 12665 6515 12699
rect 7006 12696 7012 12708
rect 6967 12668 7012 12696
rect 6457 12659 6515 12665
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 10870 12696 10876 12708
rect 10831 12668 10876 12696
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 10965 12699 11023 12705
rect 10965 12665 10977 12699
rect 11011 12696 11023 12699
rect 11146 12696 11152 12708
rect 11011 12668 11152 12696
rect 11011 12665 11023 12668
rect 10965 12659 11023 12665
rect 3510 12628 3516 12640
rect 3471 12600 3516 12628
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 6086 12628 6092 12640
rect 6047 12600 6092 12628
rect 6086 12588 6092 12600
rect 6144 12588 6150 12640
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10134 12628 10140 12640
rect 10091 12600 10140 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10134 12588 10140 12600
rect 10192 12628 10198 12640
rect 10689 12631 10747 12637
rect 10689 12628 10701 12631
rect 10192 12600 10701 12628
rect 10192 12588 10198 12600
rect 10689 12597 10701 12600
rect 10735 12628 10747 12631
rect 10980 12628 11008 12659
rect 11146 12656 11152 12668
rect 11204 12656 11210 12708
rect 10735 12600 11008 12628
rect 10735 12597 10747 12600
rect 10689 12591 10747 12597
rect 11882 12588 11888 12640
rect 11940 12628 11946 12640
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 11940 12600 12173 12628
rect 11940 12588 11946 12600
rect 12161 12597 12173 12600
rect 12207 12628 12219 12631
rect 12544 12628 12572 12727
rect 13170 12724 13176 12736
rect 13228 12724 13234 12776
rect 13354 12764 13360 12776
rect 13315 12736 13360 12764
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 13725 12767 13783 12773
rect 13725 12733 13737 12767
rect 13771 12764 13783 12767
rect 14090 12764 14096 12776
rect 13771 12736 14096 12764
rect 13771 12733 13783 12736
rect 13725 12727 13783 12733
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 13740 12696 13768 12727
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 15764 12764 15792 12872
rect 16022 12860 16028 12872
rect 16080 12860 16086 12912
rect 17402 12860 17408 12912
rect 17460 12900 17466 12912
rect 18417 12903 18475 12909
rect 18417 12900 18429 12903
rect 17460 12872 18429 12900
rect 17460 12860 17466 12872
rect 18417 12869 18429 12872
rect 18463 12869 18475 12903
rect 18417 12863 18475 12869
rect 18506 12860 18512 12912
rect 18564 12900 18570 12912
rect 23382 12900 23388 12912
rect 18564 12872 23388 12900
rect 18564 12860 18570 12872
rect 23382 12860 23388 12872
rect 23440 12860 23446 12912
rect 19426 12832 19432 12844
rect 19387 12804 19432 12832
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12832 20131 12835
rect 20162 12832 20168 12844
rect 20119 12804 20168 12832
rect 20119 12801 20131 12804
rect 20073 12795 20131 12801
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 16393 12767 16451 12773
rect 16393 12764 16405 12767
rect 15764 12736 16405 12764
rect 16393 12733 16405 12736
rect 16439 12764 16451 12767
rect 16482 12764 16488 12776
rect 16540 12773 16546 12776
rect 16540 12767 16578 12773
rect 16439 12736 16488 12764
rect 16439 12733 16451 12736
rect 16393 12727 16451 12733
rect 16482 12724 16488 12736
rect 16566 12733 16578 12767
rect 18230 12764 18236 12776
rect 18191 12736 18236 12764
rect 16540 12727 16578 12733
rect 16540 12724 16546 12727
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12764 24639 12767
rect 25130 12764 25136 12776
rect 24627 12736 25136 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 25130 12724 25136 12736
rect 25188 12724 25194 12776
rect 13998 12696 14004 12708
rect 12676 12668 13768 12696
rect 13959 12668 14004 12696
rect 12676 12656 12682 12668
rect 13998 12656 14004 12668
rect 14056 12656 14062 12708
rect 15010 12696 15016 12708
rect 14971 12668 15016 12696
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 15105 12699 15163 12705
rect 15105 12665 15117 12699
rect 15151 12665 15163 12699
rect 15105 12659 15163 12665
rect 13078 12628 13084 12640
rect 12207 12600 13084 12628
rect 12207 12597 12219 12600
rect 12161 12591 12219 12597
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 14642 12588 14648 12640
rect 14700 12628 14706 12640
rect 14737 12631 14795 12637
rect 14737 12628 14749 12631
rect 14700 12600 14749 12628
rect 14700 12588 14706 12600
rect 14737 12597 14749 12600
rect 14783 12628 14795 12631
rect 15120 12628 15148 12659
rect 17310 12656 17316 12708
rect 17368 12696 17374 12708
rect 17770 12696 17776 12708
rect 17368 12668 17776 12696
rect 17368 12656 17374 12668
rect 17770 12656 17776 12668
rect 17828 12656 17834 12708
rect 19521 12699 19579 12705
rect 19521 12665 19533 12699
rect 19567 12665 19579 12699
rect 21266 12696 21272 12708
rect 21227 12668 21272 12696
rect 19521 12659 19579 12665
rect 14783 12600 15148 12628
rect 14783 12597 14795 12600
rect 14737 12591 14795 12597
rect 15930 12588 15936 12640
rect 15988 12628 15994 12640
rect 17034 12628 17040 12640
rect 15988 12600 17040 12628
rect 15988 12588 15994 12600
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 17862 12628 17868 12640
rect 17823 12600 17868 12628
rect 17862 12588 17868 12600
rect 17920 12588 17926 12640
rect 18414 12588 18420 12640
rect 18472 12628 18478 12640
rect 18785 12631 18843 12637
rect 18785 12628 18797 12631
rect 18472 12600 18797 12628
rect 18472 12588 18478 12600
rect 18785 12597 18797 12600
rect 18831 12597 18843 12631
rect 18785 12591 18843 12597
rect 19058 12588 19064 12640
rect 19116 12628 19122 12640
rect 19245 12631 19303 12637
rect 19245 12628 19257 12631
rect 19116 12600 19257 12628
rect 19116 12588 19122 12600
rect 19245 12597 19257 12600
rect 19291 12628 19303 12631
rect 19536 12628 19564 12659
rect 21266 12656 21272 12668
rect 21324 12656 21330 12708
rect 21358 12656 21364 12708
rect 21416 12696 21422 12708
rect 21416 12668 21461 12696
rect 21416 12656 21422 12668
rect 21542 12656 21548 12708
rect 21600 12696 21606 12708
rect 21910 12696 21916 12708
rect 21600 12668 21916 12696
rect 21600 12656 21606 12668
rect 21910 12656 21916 12668
rect 21968 12656 21974 12708
rect 22002 12656 22008 12708
rect 22060 12696 22066 12708
rect 23198 12696 23204 12708
rect 22060 12668 23204 12696
rect 22060 12656 22066 12668
rect 23198 12656 23204 12668
rect 23256 12696 23262 12708
rect 24210 12696 24216 12708
rect 23256 12668 24216 12696
rect 23256 12656 23262 12668
rect 24210 12656 24216 12668
rect 24268 12656 24274 12708
rect 21376 12628 21404 12656
rect 22830 12628 22836 12640
rect 19291 12600 21404 12628
rect 22791 12600 22836 12628
rect 19291 12597 19303 12600
rect 19245 12591 19303 12597
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 24026 12588 24032 12640
rect 24084 12628 24090 12640
rect 24670 12628 24676 12640
rect 24084 12600 24676 12628
rect 24084 12588 24090 12600
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 3326 12424 3332 12436
rect 3287 12396 3332 12424
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 3694 12424 3700 12436
rect 3655 12396 3700 12424
rect 3694 12384 3700 12396
rect 3752 12424 3758 12436
rect 4338 12424 4344 12436
rect 3752 12396 4344 12424
rect 3752 12384 3758 12396
rect 4338 12384 4344 12396
rect 4396 12424 4402 12436
rect 4798 12424 4804 12436
rect 4396 12396 4804 12424
rect 4396 12384 4402 12396
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 4982 12424 4988 12436
rect 4943 12396 4988 12424
rect 4982 12384 4988 12396
rect 5040 12384 5046 12436
rect 6917 12427 6975 12433
rect 6917 12393 6929 12427
rect 6963 12424 6975 12427
rect 7006 12424 7012 12436
rect 6963 12396 7012 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 8113 12427 8171 12433
rect 8113 12393 8125 12427
rect 8159 12424 8171 12427
rect 8478 12424 8484 12436
rect 8159 12396 8484 12424
rect 8159 12393 8171 12396
rect 8113 12387 8171 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8711 12427 8769 12433
rect 8711 12393 8723 12427
rect 8757 12424 8769 12427
rect 8846 12424 8852 12436
rect 8757 12396 8852 12424
rect 8757 12393 8769 12396
rect 8711 12387 8769 12393
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 11146 12424 11152 12436
rect 11107 12396 11152 12424
rect 11146 12384 11152 12396
rect 11204 12384 11210 12436
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 12897 12427 12955 12433
rect 12897 12424 12909 12427
rect 12676 12396 12909 12424
rect 12676 12384 12682 12396
rect 12897 12393 12909 12396
rect 12943 12393 12955 12427
rect 12897 12387 12955 12393
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 15010 12424 15016 12436
rect 13872 12396 13917 12424
rect 14971 12396 15016 12424
rect 13872 12384 13878 12396
rect 15010 12384 15016 12396
rect 15068 12424 15074 12436
rect 15286 12424 15292 12436
rect 15068 12396 15292 12424
rect 15068 12384 15074 12396
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 16666 12424 16672 12436
rect 16627 12396 16672 12424
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 17862 12384 17868 12436
rect 17920 12424 17926 12436
rect 18785 12427 18843 12433
rect 18785 12424 18797 12427
rect 17920 12396 18797 12424
rect 17920 12384 17926 12396
rect 18785 12393 18797 12396
rect 18831 12393 18843 12427
rect 18785 12387 18843 12393
rect 21821 12427 21879 12433
rect 21821 12393 21833 12427
rect 21867 12424 21879 12427
rect 21910 12424 21916 12436
rect 21867 12396 21916 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 22051 12427 22109 12433
rect 22051 12393 22063 12427
rect 22097 12424 22109 12427
rect 22554 12424 22560 12436
rect 22097 12396 22560 12424
rect 22097 12393 22109 12396
rect 22051 12387 22109 12393
rect 22554 12384 22560 12396
rect 22612 12424 22618 12436
rect 22830 12424 22836 12436
rect 22612 12396 22836 12424
rect 22612 12384 22618 12396
rect 22830 12384 22836 12396
rect 22888 12384 22894 12436
rect 25130 12424 25136 12436
rect 25091 12396 25136 12424
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 4154 12316 4160 12368
rect 4212 12356 4218 12368
rect 6457 12359 6515 12365
rect 6457 12356 6469 12359
rect 4212 12328 6469 12356
rect 4212 12316 4218 12328
rect 6457 12325 6469 12328
rect 6503 12356 6515 12359
rect 6822 12356 6828 12368
rect 6503 12328 6828 12356
rect 6503 12325 6515 12328
rect 6457 12319 6515 12325
rect 6822 12316 6828 12328
rect 6880 12316 6886 12368
rect 7190 12356 7196 12368
rect 7151 12328 7196 12356
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 9950 12316 9956 12368
rect 10008 12356 10014 12368
rect 10591 12359 10649 12365
rect 10591 12356 10603 12359
rect 10008 12328 10603 12356
rect 10008 12316 10014 12328
rect 10591 12325 10603 12328
rect 10637 12356 10649 12359
rect 11054 12356 11060 12368
rect 10637 12328 11060 12356
rect 10637 12325 10649 12328
rect 10591 12319 10649 12325
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 12158 12356 12164 12368
rect 12071 12328 12164 12356
rect 12158 12316 12164 12328
rect 12216 12356 12222 12368
rect 13354 12356 13360 12368
rect 12216 12328 13360 12356
rect 12216 12316 12222 12328
rect 13354 12316 13360 12328
rect 13412 12316 13418 12368
rect 15470 12356 15476 12368
rect 14384 12328 15476 12356
rect 14384 12300 14412 12328
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 17310 12356 17316 12368
rect 17271 12328 17316 12356
rect 17310 12316 17316 12328
rect 17368 12316 17374 12368
rect 17494 12316 17500 12368
rect 17552 12356 17558 12368
rect 17552 12328 17908 12356
rect 17552 12316 17558 12328
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12288 1823 12291
rect 1854 12288 1860 12300
rect 1811 12260 1860 12288
rect 1811 12257 1823 12260
rect 1765 12251 1823 12257
rect 1854 12248 1860 12260
rect 1912 12288 1918 12300
rect 2041 12291 2099 12297
rect 2041 12288 2053 12291
rect 1912 12260 2053 12288
rect 1912 12248 1918 12260
rect 2041 12257 2053 12260
rect 2087 12257 2099 12291
rect 2682 12288 2688 12300
rect 2643 12260 2688 12288
rect 2041 12251 2099 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 3234 12248 3240 12300
rect 3292 12288 3298 12300
rect 4614 12288 4620 12300
rect 3292 12260 4620 12288
rect 3292 12248 3298 12260
rect 4614 12248 4620 12260
rect 4672 12288 4678 12300
rect 4709 12291 4767 12297
rect 4709 12288 4721 12291
rect 4672 12260 4721 12288
rect 4672 12248 4678 12260
rect 4709 12257 4721 12260
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 5169 12291 5227 12297
rect 5169 12288 5181 12291
rect 4856 12260 5181 12288
rect 4856 12248 4862 12260
rect 5169 12257 5181 12260
rect 5215 12257 5227 12291
rect 5442 12288 5448 12300
rect 5169 12251 5227 12257
rect 5276 12260 5448 12288
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4304 12192 4537 12220
rect 4304 12180 4310 12192
rect 4525 12189 4537 12192
rect 4571 12220 4583 12223
rect 5276 12220 5304 12260
rect 5442 12248 5448 12260
rect 5500 12288 5506 12300
rect 5537 12291 5595 12297
rect 5537 12288 5549 12291
rect 5500 12260 5549 12288
rect 5500 12248 5506 12260
rect 5537 12257 5549 12260
rect 5583 12257 5595 12291
rect 5537 12251 5595 12257
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12288 5963 12291
rect 6086 12288 6092 12300
rect 5951 12260 6092 12288
rect 5951 12257 5963 12260
rect 5905 12251 5963 12257
rect 4571 12192 5304 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 5350 12180 5356 12232
rect 5408 12220 5414 12232
rect 5920 12220 5948 12251
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 8110 12248 8116 12300
rect 8168 12288 8174 12300
rect 8608 12291 8666 12297
rect 8608 12288 8620 12291
rect 8168 12260 8620 12288
rect 8168 12248 8174 12260
rect 8608 12257 8620 12260
rect 8654 12257 8666 12291
rect 12250 12288 12256 12300
rect 12211 12260 12256 12288
rect 8608 12251 8666 12257
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 14366 12288 14372 12300
rect 14279 12260 14372 12288
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 17880 12288 17908 12328
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 18325 12359 18383 12365
rect 18325 12356 18337 12359
rect 18288 12328 18337 12356
rect 18288 12316 18294 12328
rect 18325 12325 18337 12328
rect 18371 12356 18383 12359
rect 24075 12359 24133 12365
rect 24075 12356 24087 12359
rect 18371 12328 24087 12356
rect 18371 12325 18383 12328
rect 18325 12319 18383 12325
rect 24075 12325 24087 12328
rect 24121 12325 24133 12359
rect 24075 12319 24133 12325
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 17880 12260 18981 12288
rect 18969 12257 18981 12260
rect 19015 12288 19027 12291
rect 19058 12288 19064 12300
rect 19015 12260 19064 12288
rect 19015 12257 19027 12260
rect 18969 12251 19027 12257
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 19242 12288 19248 12300
rect 19203 12260 19248 12288
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 21980 12291 22038 12297
rect 21980 12257 21992 12291
rect 22026 12288 22038 12291
rect 22278 12288 22284 12300
rect 22026 12260 22284 12288
rect 22026 12257 22038 12260
rect 21980 12251 22038 12257
rect 22278 12248 22284 12260
rect 22336 12248 22342 12300
rect 22925 12291 22983 12297
rect 22925 12257 22937 12291
rect 22971 12288 22983 12291
rect 23014 12288 23020 12300
rect 22971 12260 23020 12288
rect 22971 12257 22983 12260
rect 22925 12251 22983 12257
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 23934 12288 23940 12300
rect 23895 12260 23940 12288
rect 23934 12248 23940 12260
rect 23992 12248 23998 12300
rect 25016 12291 25074 12297
rect 25016 12257 25028 12291
rect 25062 12288 25074 12291
rect 25498 12288 25504 12300
rect 25062 12260 25504 12288
rect 25062 12257 25074 12260
rect 25016 12251 25074 12257
rect 25498 12248 25504 12260
rect 25556 12248 25562 12300
rect 5408 12192 5948 12220
rect 7101 12223 7159 12229
rect 5408 12180 5414 12192
rect 7101 12189 7113 12223
rect 7147 12220 7159 12223
rect 7834 12220 7840 12232
rect 7147 12192 7840 12220
rect 7147 12189 7159 12192
rect 7101 12183 7159 12189
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12220 10287 12223
rect 10962 12220 10968 12232
rect 10275 12192 10968 12220
rect 10275 12189 10287 12192
rect 10229 12183 10287 12189
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 13998 12220 14004 12232
rect 13495 12192 14004 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 15378 12220 15384 12232
rect 14516 12192 15384 12220
rect 14516 12180 14522 12192
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 15654 12220 15660 12232
rect 15615 12192 15660 12220
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 16942 12180 16948 12232
rect 17000 12220 17006 12232
rect 17221 12223 17279 12229
rect 17221 12220 17233 12223
rect 17000 12192 17233 12220
rect 17000 12180 17006 12192
rect 17221 12189 17233 12192
rect 17267 12189 17279 12223
rect 17221 12183 17279 12189
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12220 17923 12223
rect 18782 12220 18788 12232
rect 17911 12192 18788 12220
rect 17911 12189 17923 12192
rect 17865 12183 17923 12189
rect 18782 12180 18788 12192
rect 18840 12180 18846 12232
rect 20898 12220 20904 12232
rect 20859 12192 20904 12220
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 106 12112 112 12164
rect 164 12152 170 12164
rect 4062 12152 4068 12164
rect 164 12124 4068 12152
rect 164 12112 170 12124
rect 4062 12112 4068 12124
rect 4120 12112 4126 12164
rect 6822 12112 6828 12164
rect 6880 12152 6886 12164
rect 7653 12155 7711 12161
rect 7653 12152 7665 12155
rect 6880 12124 7665 12152
rect 6880 12112 6886 12124
rect 7653 12121 7665 12124
rect 7699 12121 7711 12155
rect 7653 12115 7711 12121
rect 9214 12112 9220 12164
rect 9272 12152 9278 12164
rect 11517 12155 11575 12161
rect 11517 12152 11529 12155
rect 9272 12124 11529 12152
rect 9272 12112 9278 12124
rect 11517 12121 11529 12124
rect 11563 12152 11575 12155
rect 11606 12152 11612 12164
rect 11563 12124 11612 12152
rect 11563 12121 11575 12124
rect 11517 12115 11575 12121
rect 11606 12112 11612 12124
rect 11664 12112 11670 12164
rect 12437 12155 12495 12161
rect 12437 12121 12449 12155
rect 12483 12152 12495 12155
rect 18598 12152 18604 12164
rect 12483 12124 18604 12152
rect 12483 12121 12495 12124
rect 12437 12115 12495 12121
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 21266 12112 21272 12164
rect 21324 12152 21330 12164
rect 21453 12155 21511 12161
rect 21453 12152 21465 12155
rect 21324 12124 21465 12152
rect 21324 12112 21330 12124
rect 21453 12121 21465 12124
rect 21499 12152 21511 12155
rect 23063 12155 23121 12161
rect 23063 12152 23075 12155
rect 21499 12124 23075 12152
rect 21499 12121 21511 12124
rect 21453 12115 21511 12121
rect 23063 12121 23075 12124
rect 23109 12121 23121 12155
rect 23063 12115 23121 12121
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 3786 12084 3792 12096
rect 3384 12056 3792 12084
rect 3384 12044 3390 12056
rect 3786 12044 3792 12056
rect 3844 12084 3850 12096
rect 4430 12084 4436 12096
rect 3844 12056 4436 12084
rect 3844 12044 3850 12056
rect 4430 12044 4436 12056
rect 4488 12044 4494 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 9953 12087 10011 12093
rect 9953 12084 9965 12087
rect 7156 12056 9965 12084
rect 7156 12044 7162 12056
rect 9953 12053 9965 12056
rect 9999 12084 10011 12087
rect 10226 12084 10232 12096
rect 9999 12056 10232 12084
rect 9999 12053 10011 12056
rect 9953 12047 10011 12053
rect 10226 12044 10232 12056
rect 10284 12084 10290 12096
rect 13170 12084 13176 12096
rect 10284 12056 13176 12084
rect 10284 12044 10290 12056
rect 13170 12044 13176 12056
rect 13228 12084 13234 12096
rect 13357 12087 13415 12093
rect 13357 12084 13369 12087
rect 13228 12056 13369 12084
rect 13228 12044 13234 12056
rect 13357 12053 13369 12056
rect 13403 12084 13415 12087
rect 13538 12084 13544 12096
rect 13403 12056 13544 12084
rect 13403 12053 13415 12056
rect 13357 12047 13415 12053
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 13722 12044 13728 12096
rect 13780 12084 13786 12096
rect 14366 12084 14372 12096
rect 13780 12056 14372 12084
rect 13780 12044 13786 12056
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 16390 12084 16396 12096
rect 16351 12056 16396 12084
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 19797 12087 19855 12093
rect 19797 12053 19809 12087
rect 19843 12084 19855 12087
rect 20346 12084 20352 12096
rect 19843 12056 20352 12084
rect 19843 12053 19855 12056
rect 19797 12047 19855 12053
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1302 11840 1308 11892
rect 1360 11880 1366 11892
rect 1854 11880 1860 11892
rect 1360 11852 1860 11880
rect 1360 11840 1366 11852
rect 1854 11840 1860 11852
rect 1912 11880 1918 11892
rect 2133 11883 2191 11889
rect 2133 11880 2145 11883
rect 1912 11852 2145 11880
rect 1912 11840 1918 11852
rect 2133 11849 2145 11852
rect 2179 11880 2191 11883
rect 2590 11880 2596 11892
rect 2179 11852 2596 11880
rect 2179 11849 2191 11852
rect 2133 11843 2191 11849
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 4062 11880 4068 11892
rect 4023 11852 4068 11880
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 6181 11883 6239 11889
rect 6181 11880 6193 11883
rect 4856 11852 6193 11880
rect 4856 11840 4862 11852
rect 6181 11849 6193 11852
rect 6227 11880 6239 11883
rect 7098 11880 7104 11892
rect 6227 11852 7104 11880
rect 6227 11849 6239 11852
rect 6181 11843 6239 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11880 8171 11883
rect 8941 11883 8999 11889
rect 8941 11880 8953 11883
rect 8159 11852 8953 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 8941 11849 8953 11852
rect 8987 11880 8999 11883
rect 9490 11880 9496 11892
rect 8987 11852 9496 11880
rect 8987 11849 8999 11852
rect 8941 11843 8999 11849
rect 9490 11840 9496 11852
rect 9548 11880 9554 11892
rect 11882 11880 11888 11892
rect 9548 11852 11888 11880
rect 9548 11840 9554 11852
rect 11882 11840 11888 11852
rect 11940 11880 11946 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 11940 11852 12725 11880
rect 11940 11840 11946 11852
rect 12713 11849 12725 11852
rect 12759 11880 12771 11883
rect 12759 11852 12940 11880
rect 12759 11849 12771 11852
rect 12713 11843 12771 11849
rect 3142 11772 3148 11824
rect 3200 11812 3206 11824
rect 3789 11815 3847 11821
rect 3789 11812 3801 11815
rect 3200 11784 3801 11812
rect 3200 11772 3206 11784
rect 3789 11781 3801 11784
rect 3835 11812 3847 11815
rect 4246 11812 4252 11824
rect 3835 11784 4252 11812
rect 3835 11781 3847 11784
rect 3789 11775 3847 11781
rect 4246 11772 4252 11784
rect 4304 11772 4310 11824
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 6420 11784 12173 11812
rect 6420 11772 6426 11784
rect 12161 11781 12173 11784
rect 12207 11812 12219 11815
rect 12250 11812 12256 11824
rect 12207 11784 12256 11812
rect 12207 11781 12219 11784
rect 12161 11775 12219 11781
rect 12250 11772 12256 11784
rect 12308 11772 12314 11824
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 2409 11747 2467 11753
rect 2409 11744 2421 11747
rect 1903 11716 2421 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 2409 11713 2421 11716
rect 2455 11744 2467 11747
rect 2498 11744 2504 11756
rect 2455 11716 2504 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 4982 11744 4988 11756
rect 4943 11716 4988 11744
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6687 11716 6837 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 6825 11713 6837 11716
rect 6871 11744 6883 11747
rect 7190 11744 7196 11756
rect 6871 11716 7196 11744
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 7190 11704 7196 11716
rect 7248 11704 7254 11756
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 8527 11747 8585 11753
rect 8527 11744 8539 11747
rect 7892 11716 8539 11744
rect 7892 11704 7898 11716
rect 8527 11713 8539 11716
rect 8573 11713 8585 11747
rect 8527 11707 8585 11713
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 11333 11747 11391 11753
rect 11333 11744 11345 11747
rect 8904 11716 11345 11744
rect 8904 11704 8910 11716
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11645 2375 11679
rect 2590 11676 2596 11688
rect 2551 11648 2596 11676
rect 2317 11639 2375 11645
rect 2332 11608 2360 11639
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 3878 11676 3884 11688
rect 3839 11648 3884 11676
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 5905 11679 5963 11685
rect 4126 11648 5856 11676
rect 2406 11608 2412 11620
rect 2332 11580 2412 11608
rect 2406 11568 2412 11580
rect 2464 11568 2470 11620
rect 3053 11611 3111 11617
rect 3053 11577 3065 11611
rect 3099 11608 3111 11611
rect 4126 11608 4154 11648
rect 3099 11580 4154 11608
rect 5347 11611 5405 11617
rect 3099 11577 3111 11580
rect 3053 11571 3111 11577
rect 5347 11577 5359 11611
rect 5393 11608 5405 11611
rect 5534 11608 5540 11620
rect 5393 11580 5540 11608
rect 5393 11577 5405 11580
rect 5347 11571 5405 11577
rect 5534 11568 5540 11580
rect 5592 11568 5598 11620
rect 5828 11608 5856 11648
rect 5905 11645 5917 11679
rect 5951 11676 5963 11679
rect 7006 11676 7012 11688
rect 5951 11648 7012 11676
rect 5951 11645 5963 11648
rect 5905 11639 5963 11645
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11676 7987 11679
rect 8110 11676 8116 11688
rect 7975 11648 8116 11676
rect 7975 11645 7987 11648
rect 7929 11639 7987 11645
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 8424 11679 8482 11685
rect 8424 11645 8436 11679
rect 8470 11645 8482 11679
rect 9490 11676 9496 11688
rect 9451 11648 9496 11676
rect 8424 11639 8482 11645
rect 8297 11611 8355 11617
rect 5828 11580 8248 11608
rect 3418 11540 3424 11552
rect 3379 11512 3424 11540
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 4801 11543 4859 11549
rect 4801 11509 4813 11543
rect 4847 11540 4859 11543
rect 5258 11540 5264 11552
rect 4847 11512 5264 11540
rect 4847 11509 4859 11512
rect 4801 11503 4859 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 8113 11543 8171 11549
rect 8113 11540 8125 11543
rect 6696 11512 8125 11540
rect 6696 11500 6702 11512
rect 8113 11509 8125 11512
rect 8159 11509 8171 11543
rect 8220 11540 8248 11580
rect 8297 11577 8309 11611
rect 8343 11608 8355 11611
rect 8439 11608 8467 11639
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 10226 11676 10232 11688
rect 10187 11648 10232 11676
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 10520 11685 10548 11716
rect 11333 11713 11345 11716
rect 11379 11744 11391 11747
rect 12066 11744 12072 11756
rect 11379 11716 12072 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 10505 11679 10563 11685
rect 10505 11645 10517 11679
rect 10551 11645 10563 11679
rect 10686 11676 10692 11688
rect 10647 11648 10692 11676
rect 10505 11639 10563 11645
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 11974 11676 11980 11688
rect 10796 11648 11980 11676
rect 9674 11608 9680 11620
rect 8343 11580 9680 11608
rect 8343 11577 8355 11580
rect 8297 11571 8355 11577
rect 9674 11568 9680 11580
rect 9732 11608 9738 11620
rect 10796 11608 10824 11648
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 12802 11636 12808 11688
rect 12860 11676 12866 11688
rect 12912 11685 12940 11852
rect 13998 11840 14004 11892
rect 14056 11880 14062 11892
rect 15013 11883 15071 11889
rect 15013 11880 15025 11883
rect 14056 11852 15025 11880
rect 14056 11840 14062 11852
rect 15013 11849 15025 11852
rect 15059 11849 15071 11883
rect 15013 11843 15071 11849
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15657 11883 15715 11889
rect 15657 11880 15669 11883
rect 15528 11852 15669 11880
rect 15528 11840 15534 11852
rect 15657 11849 15669 11852
rect 15703 11849 15715 11883
rect 19058 11880 19064 11892
rect 19019 11852 19064 11880
rect 15657 11843 15715 11849
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 19242 11840 19248 11892
rect 19300 11880 19306 11892
rect 19429 11883 19487 11889
rect 19429 11880 19441 11883
rect 19300 11852 19441 11880
rect 19300 11840 19306 11852
rect 19429 11849 19441 11852
rect 19475 11849 19487 11883
rect 23934 11880 23940 11892
rect 23895 11852 23940 11880
rect 19429 11843 19487 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 14645 11815 14703 11821
rect 14645 11812 14657 11815
rect 13872 11784 14657 11812
rect 13872 11772 13878 11784
rect 14645 11781 14657 11784
rect 14691 11812 14703 11815
rect 14826 11812 14832 11824
rect 14691 11784 14832 11812
rect 14691 11781 14703 11784
rect 14645 11775 14703 11781
rect 14826 11772 14832 11784
rect 14884 11772 14890 11824
rect 16942 11812 16948 11824
rect 16903 11784 16948 11812
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 17310 11772 17316 11824
rect 17368 11812 17374 11824
rect 17405 11815 17463 11821
rect 17405 11812 17417 11815
rect 17368 11784 17417 11812
rect 17368 11772 17374 11784
rect 17405 11781 17417 11784
rect 17451 11812 17463 11815
rect 24762 11812 24768 11824
rect 17451 11784 21220 11812
rect 24723 11784 24768 11812
rect 17451 11781 17463 11784
rect 17405 11775 17463 11781
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11744 15255 11747
rect 15286 11744 15292 11756
rect 15243 11716 15292 11744
rect 15243 11713 15255 11716
rect 15197 11707 15255 11713
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 18782 11744 18788 11756
rect 18743 11716 18788 11744
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12860 11648 12909 11676
rect 12860 11636 12866 11648
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 13538 11676 13544 11688
rect 13499 11648 13544 11676
rect 12897 11639 12955 11645
rect 13538 11636 13544 11648
rect 13596 11636 13602 11688
rect 13814 11676 13820 11688
rect 13786 11636 13820 11676
rect 13872 11676 13878 11688
rect 14090 11676 14096 11688
rect 13872 11648 13917 11676
rect 14051 11648 14096 11676
rect 13872 11636 13878 11648
rect 14090 11636 14096 11648
rect 14148 11636 14154 11688
rect 20346 11676 20352 11688
rect 20307 11648 20352 11676
rect 20346 11636 20352 11648
rect 20404 11636 20410 11688
rect 21192 11685 21220 11784
rect 24762 11772 24768 11784
rect 24820 11772 24826 11824
rect 25498 11744 25504 11756
rect 25459 11716 25504 11744
rect 25498 11704 25504 11716
rect 25556 11704 25562 11756
rect 21177 11679 21235 11685
rect 21177 11645 21189 11679
rect 21223 11676 21235 11679
rect 21361 11679 21419 11685
rect 21361 11676 21373 11679
rect 21223 11648 21373 11676
rect 21223 11645 21235 11648
rect 21177 11639 21235 11645
rect 21361 11645 21373 11648
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 24118 11636 24124 11688
rect 24176 11676 24182 11688
rect 24581 11679 24639 11685
rect 24581 11676 24593 11679
rect 24176 11648 24593 11676
rect 24176 11636 24182 11648
rect 24581 11645 24593 11648
rect 24627 11676 24639 11679
rect 25133 11679 25191 11685
rect 25133 11676 25145 11679
rect 24627 11648 25145 11676
rect 24627 11645 24639 11648
rect 24581 11639 24639 11645
rect 25133 11645 25145 11648
rect 25179 11645 25191 11679
rect 25133 11639 25191 11645
rect 10962 11608 10968 11620
rect 9732 11580 10824 11608
rect 10923 11580 10968 11608
rect 9732 11568 9738 11580
rect 10962 11568 10968 11580
rect 11020 11568 11026 11620
rect 13786 11608 13814 11636
rect 14366 11608 14372 11620
rect 11808 11580 13814 11608
rect 14327 11580 14372 11608
rect 8846 11540 8852 11552
rect 8220 11512 8852 11540
rect 8113 11503 8171 11509
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 9401 11543 9459 11549
rect 9401 11509 9413 11543
rect 9447 11540 9459 11543
rect 9490 11540 9496 11552
rect 9447 11512 9496 11540
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 9490 11500 9496 11512
rect 9548 11540 9554 11552
rect 10686 11540 10692 11552
rect 9548 11512 10692 11540
rect 9548 11500 9554 11512
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 11808 11549 11836 11580
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 16390 11608 16396 11620
rect 16351 11580 16396 11608
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 16485 11611 16543 11617
rect 16485 11577 16497 11611
rect 16531 11608 16543 11611
rect 17770 11608 17776 11620
rect 16531 11580 17776 11608
rect 16531 11577 16543 11580
rect 16485 11571 16543 11577
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11756 11512 11805 11540
rect 11756 11500 11762 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 16209 11543 16267 11549
rect 16209 11509 16221 11543
rect 16255 11540 16267 11543
rect 16500 11540 16528 11571
rect 17770 11568 17776 11580
rect 17828 11568 17834 11620
rect 18138 11608 18144 11620
rect 18099 11580 18144 11608
rect 18138 11568 18144 11580
rect 18196 11568 18202 11620
rect 18233 11611 18291 11617
rect 18233 11577 18245 11611
rect 18279 11577 18291 11611
rect 21269 11611 21327 11617
rect 21269 11608 21281 11611
rect 18233 11571 18291 11577
rect 18937 11580 21281 11608
rect 16255 11512 16528 11540
rect 17865 11543 17923 11549
rect 16255 11509 16267 11512
rect 16209 11503 16267 11509
rect 17865 11509 17877 11543
rect 17911 11540 17923 11543
rect 18248 11540 18276 11571
rect 18937 11540 18965 11580
rect 21269 11577 21281 11580
rect 21315 11577 21327 11611
rect 21269 11571 21327 11577
rect 20162 11540 20168 11552
rect 17911 11512 18965 11540
rect 20123 11512 20168 11540
rect 17911 11509 17923 11512
rect 17865 11503 17923 11509
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 22278 11540 22284 11552
rect 22239 11512 22284 11540
rect 22278 11500 22284 11512
rect 22336 11500 22342 11552
rect 23014 11540 23020 11552
rect 22927 11512 23020 11540
rect 23014 11500 23020 11512
rect 23072 11540 23078 11552
rect 23566 11540 23572 11552
rect 23072 11512 23572 11540
rect 23072 11500 23078 11512
rect 23566 11500 23572 11512
rect 23624 11500 23630 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 1673 11339 1731 11345
rect 1673 11336 1685 11339
rect 1452 11308 1685 11336
rect 1452 11296 1458 11308
rect 1673 11305 1685 11308
rect 1719 11305 1731 11339
rect 1673 11299 1731 11305
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 2682 11336 2688 11348
rect 2179 11308 2688 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 3510 11336 3516 11348
rect 3471 11308 3516 11336
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 3878 11336 3884 11348
rect 3839 11308 3884 11336
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 4890 11336 4896 11348
rect 4672 11308 4896 11336
rect 4672 11296 4678 11308
rect 4890 11296 4896 11308
rect 4948 11336 4954 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 4948 11308 5181 11336
rect 4948 11296 4954 11308
rect 5169 11305 5181 11308
rect 5215 11336 5227 11339
rect 6638 11336 6644 11348
rect 5215 11308 6644 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 6733 11339 6791 11345
rect 6733 11305 6745 11339
rect 6779 11336 6791 11339
rect 7006 11336 7012 11348
rect 6779 11308 7012 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7834 11336 7840 11348
rect 7795 11308 7840 11336
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11379 11339 11437 11345
rect 11379 11336 11391 11339
rect 10928 11308 11391 11336
rect 10928 11296 10934 11308
rect 11379 11305 11391 11308
rect 11425 11305 11437 11339
rect 12158 11336 12164 11348
rect 12119 11308 12164 11336
rect 11379 11299 11437 11305
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 12526 11336 12532 11348
rect 12487 11308 12532 11336
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 15378 11296 15384 11348
rect 15436 11336 15442 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 15436 11308 15485 11336
rect 15436 11296 15442 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 16206 11296 16212 11348
rect 16264 11336 16270 11348
rect 17543 11339 17601 11345
rect 17543 11336 17555 11339
rect 16264 11308 17555 11336
rect 16264 11296 16270 11308
rect 17543 11305 17555 11308
rect 17589 11305 17601 11339
rect 17543 11299 17601 11305
rect 19613 11339 19671 11345
rect 19613 11305 19625 11339
rect 19659 11305 19671 11339
rect 19613 11299 19671 11305
rect 4065 11271 4123 11277
rect 4065 11268 4077 11271
rect 2516 11240 4077 11268
rect 2516 11212 2544 11240
rect 4065 11237 4077 11240
rect 4111 11237 4123 11271
rect 4065 11231 4123 11237
rect 5951 11271 6009 11277
rect 5951 11237 5963 11271
rect 5997 11268 6009 11271
rect 9214 11268 9220 11280
rect 5997 11240 9220 11268
rect 5997 11237 6009 11240
rect 5951 11231 6009 11237
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 9306 11228 9312 11280
rect 9364 11268 9370 11280
rect 9861 11271 9919 11277
rect 9861 11268 9873 11271
rect 9364 11240 9873 11268
rect 9364 11228 9370 11240
rect 9861 11237 9873 11240
rect 9907 11268 9919 11271
rect 10226 11268 10232 11280
rect 9907 11240 10232 11268
rect 9907 11237 9919 11240
rect 9861 11231 9919 11237
rect 10226 11228 10232 11240
rect 10284 11228 10290 11280
rect 10962 11228 10968 11280
rect 11020 11268 11026 11280
rect 11057 11271 11115 11277
rect 11057 11268 11069 11271
rect 11020 11240 11069 11268
rect 11020 11228 11026 11240
rect 11057 11237 11069 11240
rect 11103 11237 11115 11271
rect 11057 11231 11115 11237
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 2682 11200 2688 11212
rect 2556 11172 2601 11200
rect 2643 11172 2688 11200
rect 2556 11160 2562 11172
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 4246 11200 4252 11212
rect 4207 11172 4252 11200
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 5864 11203 5922 11209
rect 5864 11169 5876 11203
rect 5910 11200 5922 11203
rect 6362 11200 6368 11212
rect 5910 11172 6368 11200
rect 5910 11169 5922 11172
rect 5864 11163 5922 11169
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 7469 11203 7527 11209
rect 7469 11169 7481 11203
rect 7515 11200 7527 11203
rect 8018 11200 8024 11212
rect 7515 11172 8024 11200
rect 7515 11169 7527 11172
rect 7469 11163 7527 11169
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 8570 11200 8576 11212
rect 8531 11172 8576 11200
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 10410 11160 10416 11212
rect 10468 11200 10474 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 10468 11172 11253 11200
rect 10468 11160 10474 11172
rect 11241 11169 11253 11172
rect 11287 11200 11299 11203
rect 11330 11200 11336 11212
rect 11287 11172 11336 11200
rect 11287 11169 11299 11172
rect 11241 11163 11299 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 12544 11200 12572 11296
rect 14826 11228 14832 11280
rect 14884 11268 14890 11280
rect 15978 11271 16036 11277
rect 15978 11268 15990 11271
rect 14884 11240 15990 11268
rect 14884 11228 14890 11240
rect 15978 11237 15990 11240
rect 16024 11237 16036 11271
rect 15978 11231 16036 11237
rect 18414 11228 18420 11280
rect 18472 11268 18478 11280
rect 19014 11271 19072 11277
rect 19014 11268 19026 11271
rect 18472 11240 19026 11268
rect 18472 11228 18478 11240
rect 19014 11237 19026 11240
rect 19060 11237 19072 11271
rect 19628 11268 19656 11299
rect 20346 11268 20352 11280
rect 19628 11240 20352 11268
rect 19014 11231 19072 11237
rect 20346 11228 20352 11240
rect 20404 11268 20410 11280
rect 21085 11271 21143 11277
rect 21085 11268 21097 11271
rect 20404 11240 21097 11268
rect 20404 11228 20410 11240
rect 21085 11237 21097 11240
rect 21131 11268 21143 11271
rect 21450 11268 21456 11280
rect 21131 11240 21456 11268
rect 21131 11237 21143 11240
rect 21085 11231 21143 11237
rect 21450 11228 21456 11240
rect 21508 11228 21514 11280
rect 12713 11203 12771 11209
rect 12713 11200 12725 11203
rect 12544 11172 12725 11200
rect 12713 11169 12725 11172
rect 12759 11169 12771 11203
rect 12713 11163 12771 11169
rect 12986 11160 12992 11212
rect 13044 11200 13050 11212
rect 13173 11203 13231 11209
rect 13173 11200 13185 11203
rect 13044 11172 13185 11200
rect 13044 11160 13050 11172
rect 13173 11169 13185 11172
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 13354 11160 13360 11212
rect 13412 11200 13418 11212
rect 13541 11203 13599 11209
rect 13541 11200 13553 11203
rect 13412 11172 13553 11200
rect 13412 11160 13418 11172
rect 13541 11169 13553 11172
rect 13587 11200 13599 11203
rect 13630 11200 13636 11212
rect 13587 11172 13636 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 14090 11200 14096 11212
rect 14051 11172 14096 11200
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 14366 11160 14372 11212
rect 14424 11200 14430 11212
rect 15654 11200 15660 11212
rect 14424 11172 15660 11200
rect 14424 11160 14430 11172
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 16577 11203 16635 11209
rect 16577 11169 16589 11203
rect 16623 11200 16635 11203
rect 17310 11200 17316 11212
rect 16623 11172 17316 11200
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 17494 11209 17500 11212
rect 17472 11203 17500 11209
rect 17472 11200 17484 11203
rect 17407 11172 17484 11200
rect 17472 11169 17484 11172
rect 17552 11200 17558 11212
rect 18506 11200 18512 11212
rect 17552 11172 18512 11200
rect 17472 11163 17500 11169
rect 17494 11160 17500 11163
rect 17552 11160 17558 11172
rect 18506 11160 18512 11172
rect 18564 11160 18570 11212
rect 22532 11203 22590 11209
rect 22532 11169 22544 11203
rect 22578 11200 22590 11203
rect 22830 11200 22836 11212
rect 22578 11172 22836 11200
rect 22578 11169 22590 11172
rect 22532 11163 22590 11169
rect 22830 11160 22836 11172
rect 22888 11160 22894 11212
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 8711 11135 8769 11141
rect 3191 11104 3924 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3896 11064 3924 11104
rect 8711 11101 8723 11135
rect 8757 11132 8769 11135
rect 9122 11132 9128 11144
rect 8757 11104 9128 11132
rect 8757 11101 8769 11104
rect 8711 11095 8769 11101
rect 9122 11092 9128 11104
rect 9180 11132 9186 11144
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9180 11104 9781 11132
rect 9180 11092 9186 11104
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 10042 11132 10048 11144
rect 10003 11104 10048 11132
rect 9769 11095 9827 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 14185 11135 14243 11141
rect 14185 11101 14197 11135
rect 14231 11132 14243 11135
rect 18693 11135 18751 11141
rect 18693 11132 18705 11135
rect 14231 11104 18705 11132
rect 14231 11101 14243 11104
rect 14185 11095 14243 11101
rect 18693 11101 18705 11104
rect 18739 11132 18751 11135
rect 19150 11132 19156 11144
rect 18739 11104 19156 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11132 21051 11135
rect 21266 11132 21272 11144
rect 21039 11104 21272 11132
rect 21039 11101 21051 11104
rect 20993 11095 21051 11101
rect 21266 11092 21272 11104
rect 21324 11092 21330 11144
rect 10870 11064 10876 11076
rect 3896 11036 10876 11064
rect 10870 11024 10876 11036
rect 10928 11064 10934 11076
rect 11698 11064 11704 11076
rect 10928 11036 11704 11064
rect 10928 11024 10934 11036
rect 11698 11024 11704 11036
rect 11756 11024 11762 11076
rect 20438 11024 20444 11076
rect 20496 11064 20502 11076
rect 21082 11064 21088 11076
rect 20496 11036 21088 11064
rect 20496 11024 20502 11036
rect 21082 11024 21088 11036
rect 21140 11064 21146 11076
rect 21545 11067 21603 11073
rect 21545 11064 21557 11067
rect 21140 11036 21557 11064
rect 21140 11024 21146 11036
rect 21545 11033 21557 11036
rect 21591 11033 21603 11067
rect 21545 11027 21603 11033
rect 5534 10996 5540 11008
rect 5447 10968 5540 10996
rect 5534 10956 5540 10968
rect 5592 10996 5598 11008
rect 6638 10996 6644 11008
rect 5592 10968 6644 10996
rect 5592 10956 5598 10968
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 7098 10996 7104 11008
rect 7059 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 9306 10996 9312 11008
rect 9267 10968 9312 10996
rect 9306 10956 9312 10968
rect 9364 10956 9370 11008
rect 10781 10999 10839 11005
rect 10781 10965 10793 10999
rect 10827 10996 10839 10999
rect 11054 10996 11060 11008
rect 10827 10968 11060 10996
rect 10827 10965 10839 10968
rect 10781 10959 10839 10965
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 11790 10996 11796 11008
rect 11751 10968 11796 10996
rect 11790 10956 11796 10968
rect 11848 10956 11854 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 17129 10999 17187 11005
rect 17129 10996 17141 10999
rect 17000 10968 17141 10996
rect 17000 10956 17006 10968
rect 17129 10965 17141 10968
rect 17175 10965 17187 10999
rect 18046 10996 18052 11008
rect 18007 10968 18052 10996
rect 17129 10959 17187 10965
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 18138 10956 18144 11008
rect 18196 10996 18202 11008
rect 22603 10999 22661 11005
rect 22603 10996 22615 10999
rect 18196 10968 22615 10996
rect 18196 10956 18202 10968
rect 22603 10965 22615 10968
rect 22649 10965 22661 10999
rect 22603 10959 22661 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2222 10792 2228 10804
rect 2183 10764 2228 10792
rect 2222 10752 2228 10764
rect 2280 10792 2286 10804
rect 2590 10792 2596 10804
rect 2280 10764 2596 10792
rect 2280 10752 2286 10764
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 3418 10792 3424 10804
rect 3379 10764 3424 10792
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 5040 10764 5457 10792
rect 5040 10752 5046 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6362 10792 6368 10804
rect 5951 10764 6368 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9582 10792 9588 10804
rect 9171 10764 9588 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 10226 10792 10232 10804
rect 10187 10764 10232 10792
rect 10226 10752 10232 10764
rect 10284 10792 10290 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 10284 10764 10609 10792
rect 10284 10752 10290 10764
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 10597 10755 10655 10761
rect 2406 10724 2412 10736
rect 2319 10696 2412 10724
rect 2406 10684 2412 10696
rect 2464 10724 2470 10736
rect 3436 10724 3464 10752
rect 2464 10696 3464 10724
rect 2464 10684 2470 10696
rect 8570 10684 8576 10736
rect 8628 10724 8634 10736
rect 8665 10727 8723 10733
rect 8665 10724 8677 10727
rect 8628 10696 8677 10724
rect 8628 10684 8634 10696
rect 8665 10693 8677 10696
rect 8711 10724 8723 10727
rect 10410 10724 10416 10736
rect 8711 10696 10416 10724
rect 8711 10693 8723 10696
rect 8665 10687 8723 10693
rect 10410 10684 10416 10696
rect 10468 10684 10474 10736
rect 2424 10597 2452 10684
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10656 2559 10659
rect 2590 10656 2596 10668
rect 2547 10628 2596 10656
rect 2547 10625 2559 10628
rect 2501 10619 2559 10625
rect 2590 10616 2596 10628
rect 2648 10656 2654 10668
rect 3142 10656 3148 10668
rect 2648 10628 2912 10656
rect 3103 10628 3148 10656
rect 2648 10616 2654 10628
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10557 2467 10591
rect 2409 10551 2467 10557
rect 2682 10548 2688 10600
rect 2740 10588 2746 10600
rect 2884 10588 2912 10628
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 5166 10656 5172 10668
rect 5079 10628 5172 10656
rect 4065 10591 4123 10597
rect 4065 10588 4077 10591
rect 2740 10560 2833 10588
rect 2884 10560 4077 10588
rect 2740 10548 2746 10560
rect 4065 10557 4077 10560
rect 4111 10588 4123 10591
rect 4246 10588 4252 10600
rect 4111 10560 4252 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 4522 10548 4528 10600
rect 4580 10588 4586 10600
rect 5092 10597 5120 10628
rect 5166 10616 5172 10628
rect 5224 10656 5230 10668
rect 6270 10656 6276 10668
rect 5224 10628 6276 10656
rect 5224 10616 5230 10628
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 6638 10656 6644 10668
rect 6551 10628 6644 10656
rect 6638 10616 6644 10628
rect 6696 10656 6702 10668
rect 7466 10656 7472 10668
rect 6696 10628 7472 10656
rect 6696 10616 6702 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10656 10011 10659
rect 10042 10656 10048 10668
rect 9999 10628 10048 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 4580 10560 5089 10588
rect 4580 10548 4586 10560
rect 5077 10557 5089 10560
rect 5123 10557 5135 10591
rect 6822 10588 6828 10600
rect 6783 10560 6828 10588
rect 5077 10551 5135 10557
rect 6822 10548 6828 10560
rect 6880 10588 6886 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 6880 10560 8033 10588
rect 6880 10548 6886 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 1949 10523 2007 10529
rect 1949 10489 1961 10523
rect 1995 10520 2007 10523
rect 2314 10520 2320 10532
rect 1995 10492 2320 10520
rect 1995 10489 2007 10492
rect 1949 10483 2007 10489
rect 2314 10480 2320 10492
rect 2372 10520 2378 10532
rect 2700 10520 2728 10548
rect 4430 10520 4436 10532
rect 2372 10492 2728 10520
rect 4391 10492 4436 10520
rect 2372 10480 2378 10492
rect 4430 10480 4436 10492
rect 4488 10480 4494 10532
rect 6273 10523 6331 10529
rect 6273 10489 6285 10523
rect 6319 10520 6331 10523
rect 7187 10523 7245 10529
rect 6319 10492 7052 10520
rect 6319 10489 6331 10492
rect 6273 10483 6331 10489
rect 7024 10452 7052 10492
rect 7187 10489 7199 10523
rect 7233 10520 7245 10523
rect 7466 10520 7472 10532
rect 7233 10492 7472 10520
rect 7233 10489 7245 10492
rect 7187 10483 7245 10489
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 9306 10520 9312 10532
rect 9267 10492 9312 10520
rect 9306 10480 9312 10492
rect 9364 10480 9370 10532
rect 9410 10523 9468 10529
rect 9410 10489 9422 10523
rect 9456 10520 9468 10523
rect 9582 10520 9588 10532
rect 9456 10492 9588 10520
rect 9456 10489 9468 10492
rect 9410 10483 9468 10489
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 10612 10520 10640 10755
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 14461 10795 14519 10801
rect 14461 10792 14473 10795
rect 14240 10764 14473 10792
rect 14240 10752 14246 10764
rect 14461 10761 14473 10764
rect 14507 10761 14519 10795
rect 14826 10792 14832 10804
rect 14787 10764 14832 10792
rect 14461 10755 14519 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 16390 10752 16396 10804
rect 16448 10792 16454 10804
rect 16448 10764 18736 10792
rect 16448 10752 16454 10764
rect 11790 10724 11796 10736
rect 10888 10696 11796 10724
rect 10888 10665 10916 10696
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 14093 10727 14151 10733
rect 14093 10693 14105 10727
rect 14139 10724 14151 10727
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 14139 10696 17785 10724
rect 14139 10693 14151 10696
rect 14093 10687 14151 10693
rect 17773 10693 17785 10696
rect 17819 10724 17831 10727
rect 18708 10724 18736 10764
rect 20162 10752 20168 10804
rect 20220 10792 20226 10804
rect 20257 10795 20315 10801
rect 20257 10792 20269 10795
rect 20220 10764 20269 10792
rect 20220 10752 20226 10764
rect 20257 10761 20269 10764
rect 20303 10761 20315 10795
rect 21450 10792 21456 10804
rect 20257 10755 20315 10761
rect 20364 10764 21312 10792
rect 21411 10764 21456 10792
rect 20364 10724 20392 10764
rect 21082 10724 21088 10736
rect 17819 10696 18644 10724
rect 18708 10696 20392 10724
rect 21043 10696 21088 10724
rect 17819 10693 17831 10696
rect 17773 10687 17831 10693
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 11146 10656 11152 10668
rect 11107 10628 11152 10656
rect 10873 10619 10931 10625
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10656 17003 10659
rect 18046 10656 18052 10668
rect 16991 10628 18052 10656
rect 16991 10625 17003 10628
rect 16945 10619 17003 10625
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18616 10665 18644 10696
rect 21082 10684 21088 10696
rect 21140 10684 21146 10736
rect 21284 10724 21312 10764
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 22830 10792 22836 10804
rect 22791 10764 22836 10792
rect 22830 10752 22836 10764
rect 22888 10752 22894 10804
rect 22143 10727 22201 10733
rect 22143 10724 22155 10727
rect 21284 10696 22155 10724
rect 22143 10693 22155 10696
rect 22189 10693 22201 10727
rect 22143 10687 22201 10693
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 20530 10656 20536 10668
rect 20443 10628 20536 10656
rect 18601 10619 18659 10625
rect 20530 10616 20536 10628
rect 20588 10656 20594 10668
rect 20898 10656 20904 10668
rect 20588 10628 20904 10656
rect 20588 10616 20594 10628
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 12713 10591 12771 10597
rect 12713 10588 12725 10591
rect 12584 10560 12725 10588
rect 12584 10548 12590 10560
rect 12713 10557 12725 10560
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 12986 10548 12992 10600
rect 13044 10588 13050 10600
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 13044 10560 13185 10588
rect 13044 10548 13050 10560
rect 13173 10557 13185 10560
rect 13219 10557 13231 10591
rect 13630 10588 13636 10600
rect 13591 10560 13636 10588
rect 13173 10551 13231 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10557 13967 10591
rect 15010 10588 15016 10600
rect 14971 10560 15016 10588
rect 13909 10551 13967 10557
rect 10965 10523 11023 10529
rect 10965 10520 10977 10523
rect 10612 10492 10977 10520
rect 10965 10489 10977 10492
rect 11011 10489 11023 10523
rect 10965 10483 11023 10489
rect 11885 10523 11943 10529
rect 11885 10489 11897 10523
rect 11931 10520 11943 10523
rect 12253 10523 12311 10529
rect 12253 10520 12265 10523
rect 11931 10492 12265 10520
rect 11931 10489 11943 10492
rect 11885 10483 11943 10489
rect 12253 10489 12265 10492
rect 12299 10520 12311 10523
rect 13004 10520 13032 10548
rect 12299 10492 13032 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 7024 10424 7757 10452
rect 7745 10421 7757 10424
rect 7791 10452 7803 10455
rect 8018 10452 8024 10464
rect 7791 10424 8024 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 11900 10452 11928 10483
rect 10744 10424 11928 10452
rect 13924 10452 13952 10551
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 15933 10591 15991 10597
rect 15933 10557 15945 10591
rect 15979 10588 15991 10591
rect 16390 10588 16396 10600
rect 15979 10560 16396 10588
rect 15979 10557 15991 10560
rect 15933 10551 15991 10557
rect 16390 10548 16396 10560
rect 16448 10548 16454 10600
rect 17494 10588 17500 10600
rect 17455 10560 17500 10588
rect 17494 10548 17500 10560
rect 17552 10588 17558 10600
rect 17954 10588 17960 10600
rect 17552 10560 17960 10588
rect 17552 10548 17558 10560
rect 17954 10548 17960 10560
rect 18012 10548 18018 10600
rect 22072 10591 22130 10597
rect 22072 10557 22084 10591
rect 22118 10588 22130 10591
rect 22462 10588 22468 10600
rect 22118 10560 22468 10588
rect 22118 10557 22130 10560
rect 22072 10551 22130 10557
rect 22462 10548 22468 10560
rect 22520 10548 22526 10600
rect 14826 10480 14832 10532
rect 14884 10520 14890 10532
rect 15334 10523 15392 10529
rect 15334 10520 15346 10523
rect 14884 10492 15346 10520
rect 14884 10480 14890 10492
rect 15334 10489 15346 10492
rect 15380 10520 15392 10523
rect 15562 10520 15568 10532
rect 15380 10492 15568 10520
rect 15380 10489 15392 10492
rect 15334 10483 15392 10489
rect 15562 10480 15568 10492
rect 15620 10520 15626 10532
rect 16209 10523 16267 10529
rect 16209 10520 16221 10523
rect 15620 10492 16221 10520
rect 15620 10480 15626 10492
rect 16209 10489 16221 10492
rect 16255 10520 16267 10523
rect 18414 10520 18420 10532
rect 16255 10492 18420 10520
rect 16255 10489 16267 10492
rect 16209 10483 16267 10489
rect 18414 10480 18420 10492
rect 18472 10520 18478 10532
rect 18922 10523 18980 10529
rect 18922 10520 18934 10523
rect 18472 10492 18934 10520
rect 18472 10480 18478 10492
rect 18922 10489 18934 10492
rect 18968 10489 18980 10523
rect 18922 10483 18980 10489
rect 20625 10523 20683 10529
rect 20625 10489 20637 10523
rect 20671 10489 20683 10523
rect 20625 10483 20683 10489
rect 14090 10452 14096 10464
rect 13924 10424 14096 10452
rect 10744 10412 10750 10424
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 19518 10452 19524 10464
rect 19479 10424 19524 10452
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 20162 10412 20168 10464
rect 20220 10452 20226 10464
rect 20640 10452 20668 10483
rect 21266 10480 21272 10532
rect 21324 10520 21330 10532
rect 21821 10523 21879 10529
rect 21821 10520 21833 10523
rect 21324 10492 21833 10520
rect 21324 10480 21330 10492
rect 21821 10489 21833 10492
rect 21867 10489 21879 10523
rect 21821 10483 21879 10489
rect 20220 10424 20668 10452
rect 20220 10412 20226 10424
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2556 10220 2789 10248
rect 2556 10208 2562 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 3418 10248 3424 10260
rect 3283 10220 3424 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 2133 10183 2191 10189
rect 2133 10149 2145 10183
rect 2179 10180 2191 10183
rect 2314 10180 2320 10192
rect 2179 10152 2320 10180
rect 2179 10149 2191 10152
rect 2133 10143 2191 10149
rect 2314 10140 2320 10152
rect 2372 10180 2378 10192
rect 3252 10180 3280 10211
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 3602 10208 3608 10260
rect 3660 10248 3666 10260
rect 4522 10248 4528 10260
rect 3660 10220 4528 10248
rect 3660 10208 3666 10220
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 6880 10220 6929 10248
rect 6880 10208 6886 10220
rect 6917 10217 6929 10220
rect 6963 10217 6975 10251
rect 9122 10248 9128 10260
rect 9083 10220 9128 10248
rect 6917 10211 6975 10217
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 11563 10251 11621 10257
rect 11563 10248 11575 10251
rect 9364 10220 11575 10248
rect 9364 10208 9370 10220
rect 11563 10217 11575 10220
rect 11609 10217 11621 10251
rect 11563 10211 11621 10217
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 12158 10248 12164 10260
rect 12115 10220 12164 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 12526 10248 12532 10260
rect 12483 10220 12532 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 2372 10152 3280 10180
rect 3789 10183 3847 10189
rect 2372 10140 2378 10152
rect 3789 10149 3801 10183
rect 3835 10180 3847 10183
rect 4062 10180 4068 10192
rect 3835 10152 4068 10180
rect 3835 10149 3847 10152
rect 3789 10143 3847 10149
rect 4062 10140 4068 10152
rect 4120 10180 4126 10192
rect 4430 10180 4436 10192
rect 4120 10152 4436 10180
rect 4120 10140 4126 10152
rect 4430 10140 4436 10152
rect 4488 10140 4494 10192
rect 5442 10140 5448 10192
rect 5500 10180 5506 10192
rect 6638 10180 6644 10192
rect 5500 10152 6644 10180
rect 5500 10140 5506 10152
rect 1302 10072 1308 10124
rect 1360 10112 1366 10124
rect 1489 10115 1547 10121
rect 1489 10112 1501 10115
rect 1360 10084 1501 10112
rect 1360 10072 1366 10084
rect 1489 10081 1501 10084
rect 1535 10081 1547 10115
rect 1489 10075 1547 10081
rect 5813 10115 5871 10121
rect 5813 10081 5825 10115
rect 5859 10081 5871 10115
rect 6270 10112 6276 10124
rect 6231 10084 6276 10112
rect 5813 10075 5871 10081
rect 5828 9976 5856 10075
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6380 10121 6408 10152
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 8018 10180 8024 10192
rect 7979 10152 8024 10180
rect 8018 10140 8024 10152
rect 8076 10140 8082 10192
rect 9493 10183 9551 10189
rect 9493 10149 9505 10183
rect 9539 10180 9551 10183
rect 9582 10180 9588 10192
rect 9539 10152 9588 10180
rect 9539 10149 9551 10152
rect 9493 10143 9551 10149
rect 9582 10140 9588 10152
rect 9640 10180 9646 10192
rect 10045 10183 10103 10189
rect 10045 10180 10057 10183
rect 9640 10152 10057 10180
rect 9640 10140 9646 10152
rect 10045 10149 10057 10152
rect 10091 10149 10103 10183
rect 10045 10143 10103 10149
rect 10597 10183 10655 10189
rect 10597 10149 10609 10183
rect 10643 10180 10655 10183
rect 11146 10180 11152 10192
rect 10643 10152 11152 10180
rect 10643 10149 10655 10152
rect 10597 10143 10655 10149
rect 11146 10140 11152 10152
rect 11204 10140 11210 10192
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10081 6423 10115
rect 6365 10075 6423 10081
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 6512 10084 6929 10112
rect 6512 10072 6518 10084
rect 6917 10081 6929 10084
rect 6963 10112 6975 10115
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 6963 10084 7481 10112
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 7469 10081 7481 10084
rect 7515 10081 7527 10115
rect 10870 10112 10876 10124
rect 10831 10084 10876 10112
rect 7469 10075 7527 10081
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 11492 10115 11550 10121
rect 11492 10081 11504 10115
rect 11538 10112 11550 10115
rect 11882 10112 11888 10124
rect 11538 10084 11888 10112
rect 11538 10081 11550 10084
rect 11492 10075 11550 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 7926 10044 7932 10056
rect 7887 10016 7932 10044
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 8202 10044 8208 10056
rect 8163 10016 8208 10044
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 7190 9976 7196 9988
rect 5828 9948 7196 9976
rect 7190 9936 7196 9948
rect 7248 9976 7254 9988
rect 7653 9979 7711 9985
rect 7653 9976 7665 9979
rect 7248 9948 7665 9976
rect 7248 9936 7254 9948
rect 7653 9945 7665 9948
rect 7699 9976 7711 9979
rect 9214 9976 9220 9988
rect 7699 9948 9220 9976
rect 7699 9945 7711 9948
rect 7653 9939 7711 9945
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 9968 9976 9996 10007
rect 10318 10004 10324 10056
rect 10376 10044 10382 10056
rect 12452 10044 12480 10211
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 15654 10248 15660 10260
rect 15615 10220 15660 10248
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 16022 10248 16028 10260
rect 15983 10220 16028 10248
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 18414 10208 18420 10260
rect 18472 10248 18478 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 18472 10220 18797 10248
rect 18472 10208 18478 10220
rect 18785 10217 18797 10220
rect 18831 10217 18843 10251
rect 19150 10248 19156 10260
rect 19111 10220 19156 10248
rect 18785 10211 18843 10217
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 20530 10248 20536 10260
rect 20491 10220 20536 10248
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 23707 10251 23765 10257
rect 20916 10220 23474 10248
rect 14369 10183 14427 10189
rect 14369 10149 14381 10183
rect 14415 10180 14427 10183
rect 15010 10180 15016 10192
rect 14415 10152 15016 10180
rect 14415 10149 14427 10152
rect 14369 10143 14427 10149
rect 15010 10140 15016 10152
rect 15068 10140 15074 10192
rect 16390 10180 16396 10192
rect 16351 10152 16396 10180
rect 16390 10140 16396 10152
rect 16448 10140 16454 10192
rect 16942 10180 16948 10192
rect 16903 10152 16948 10180
rect 16942 10140 16948 10152
rect 17000 10140 17006 10192
rect 17770 10180 17776 10192
rect 17731 10152 17776 10180
rect 17770 10140 17776 10152
rect 17828 10140 17834 10192
rect 20916 10180 20944 10220
rect 21082 10180 21088 10192
rect 19996 10152 20944 10180
rect 21043 10152 21088 10180
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 12860 10084 12909 10112
rect 12860 10072 12866 10084
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 13630 10112 13636 10124
rect 13591 10084 13636 10112
rect 12897 10075 12955 10081
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14090 10112 14096 10124
rect 13872 10084 13917 10112
rect 14051 10084 14096 10112
rect 13872 10072 13878 10084
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 17494 10072 17500 10124
rect 17552 10112 17558 10124
rect 17865 10115 17923 10121
rect 17865 10112 17877 10115
rect 17552 10084 17877 10112
rect 17552 10072 17558 10084
rect 17865 10081 17877 10084
rect 17911 10081 17923 10115
rect 17865 10075 17923 10081
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19648 10115 19706 10121
rect 19648 10112 19660 10115
rect 19484 10084 19660 10112
rect 19484 10072 19490 10084
rect 19648 10081 19660 10084
rect 19694 10112 19706 10115
rect 19996 10112 20024 10152
rect 21082 10140 21088 10152
rect 21140 10140 21146 10192
rect 23446 10180 23474 10220
rect 23707 10217 23719 10251
rect 23753 10248 23765 10251
rect 24026 10248 24032 10260
rect 23753 10220 24032 10248
rect 23753 10217 23765 10220
rect 23707 10211 23765 10217
rect 24026 10208 24032 10220
rect 24084 10208 24090 10260
rect 24762 10248 24768 10260
rect 24723 10220 24768 10248
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 25222 10180 25228 10192
rect 23446 10152 25228 10180
rect 25222 10140 25228 10152
rect 25280 10140 25286 10192
rect 19694 10084 20024 10112
rect 19694 10081 19706 10084
rect 19648 10075 19706 10081
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 23604 10115 23662 10121
rect 23604 10112 23616 10115
rect 23440 10084 23616 10112
rect 23440 10072 23446 10084
rect 23604 10081 23616 10084
rect 23650 10081 23662 10115
rect 23604 10075 23662 10081
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10112 24639 10115
rect 25130 10112 25136 10124
rect 24627 10084 25136 10112
rect 24627 10081 24639 10084
rect 24581 10075 24639 10081
rect 16298 10044 16304 10056
rect 10376 10016 12480 10044
rect 16259 10016 16304 10044
rect 10376 10004 10382 10016
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 20990 10044 20996 10056
rect 20951 10016 20996 10044
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 21266 10044 21272 10056
rect 21227 10016 21272 10044
rect 21266 10004 21272 10016
rect 21324 10004 21330 10056
rect 23290 10004 23296 10056
rect 23348 10044 23354 10056
rect 24596 10044 24624 10075
rect 25130 10072 25136 10084
rect 25188 10072 25194 10124
rect 23348 10016 24624 10044
rect 23348 10004 23354 10016
rect 11422 9976 11428 9988
rect 9968 9948 11428 9976
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 2406 9908 2412 9920
rect 2367 9880 2412 9908
rect 2406 9868 2412 9880
rect 2464 9868 2470 9920
rect 7374 9908 7380 9920
rect 7335 9880 7380 9908
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 9490 9908 9496 9920
rect 7515 9880 9496 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 11330 9908 11336 9920
rect 11291 9880 11336 9908
rect 11330 9868 11336 9880
rect 11388 9868 11394 9920
rect 12710 9908 12716 9920
rect 12671 9880 12716 9908
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 19751 9911 19809 9917
rect 19751 9877 19763 9911
rect 19797 9908 19809 9911
rect 19978 9908 19984 9920
rect 19797 9880 19984 9908
rect 19797 9877 19809 9880
rect 19751 9871 19809 9877
rect 19978 9868 19984 9880
rect 20036 9868 20042 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1854 9704 1860 9716
rect 1815 9676 1860 9704
rect 1854 9664 1860 9676
rect 1912 9664 1918 9716
rect 2406 9704 2412 9716
rect 2367 9676 2412 9704
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 3237 9707 3295 9713
rect 3237 9673 3249 9707
rect 3283 9704 3295 9707
rect 3510 9704 3516 9716
rect 3283 9676 3516 9704
rect 3283 9673 3295 9676
rect 3237 9667 3295 9673
rect 1854 9460 1860 9512
rect 1912 9500 1918 9512
rect 2041 9503 2099 9509
rect 2041 9500 2053 9503
rect 1912 9472 2053 9500
rect 1912 9460 1918 9472
rect 2041 9469 2053 9472
rect 2087 9469 2099 9503
rect 2041 9463 2099 9469
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 3436 9432 3464 9676
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 5350 9664 5356 9716
rect 5408 9704 5414 9716
rect 5629 9707 5687 9713
rect 5629 9704 5641 9707
rect 5408 9676 5641 9704
rect 5408 9664 5414 9676
rect 5629 9673 5641 9676
rect 5675 9704 5687 9707
rect 6454 9704 6460 9716
rect 5675 9676 6460 9704
rect 5675 9673 5687 9676
rect 5629 9667 5687 9673
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 12802 9664 12808 9716
rect 12860 9704 12866 9716
rect 13265 9707 13323 9713
rect 13265 9704 13277 9707
rect 12860 9676 13277 9704
rect 12860 9664 12866 9676
rect 13265 9673 13277 9676
rect 13311 9673 13323 9707
rect 13630 9704 13636 9716
rect 13591 9676 13636 9704
rect 13265 9667 13323 9673
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 16390 9664 16396 9716
rect 16448 9704 16454 9716
rect 16577 9707 16635 9713
rect 16577 9704 16589 9707
rect 16448 9676 16589 9704
rect 16448 9664 16454 9676
rect 16577 9673 16589 9676
rect 16623 9704 16635 9707
rect 17494 9704 17500 9716
rect 16623 9676 17500 9704
rect 16623 9673 16635 9676
rect 16577 9667 16635 9673
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 18966 9664 18972 9716
rect 19024 9704 19030 9716
rect 23382 9704 23388 9716
rect 19024 9676 23388 9704
rect 19024 9664 19030 9676
rect 23382 9664 23388 9676
rect 23440 9704 23446 9716
rect 23845 9707 23903 9713
rect 23845 9704 23857 9707
rect 23440 9676 23857 9704
rect 23440 9664 23446 9676
rect 23845 9673 23857 9676
rect 23891 9673 23903 9707
rect 23845 9667 23903 9673
rect 24670 9664 24676 9716
rect 24728 9704 24734 9716
rect 24765 9707 24823 9713
rect 24765 9704 24777 9707
rect 24728 9676 24777 9704
rect 24728 9664 24734 9676
rect 24765 9673 24777 9676
rect 24811 9673 24823 9707
rect 25130 9704 25136 9716
rect 25091 9676 25136 9704
rect 24765 9667 24823 9673
rect 25130 9664 25136 9676
rect 25188 9664 25194 9716
rect 3786 9596 3792 9648
rect 3844 9636 3850 9648
rect 5997 9639 6055 9645
rect 3844 9608 5120 9636
rect 3844 9596 3850 9608
rect 4246 9568 4252 9580
rect 3988 9540 4252 9568
rect 3988 9509 4016 9540
rect 4246 9528 4252 9540
rect 4304 9568 4310 9580
rect 4890 9568 4896 9580
rect 4304 9540 4896 9568
rect 4304 9528 4310 9540
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 5092 9568 5120 9608
rect 5997 9605 6009 9639
rect 6043 9636 6055 9639
rect 6270 9636 6276 9648
rect 6043 9608 6276 9636
rect 6043 9605 6055 9608
rect 5997 9599 6055 9605
rect 6270 9596 6276 9608
rect 6328 9636 6334 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 6328 9608 6653 9636
rect 6328 9596 6334 9608
rect 6641 9605 6653 9608
rect 6687 9636 6699 9639
rect 7558 9636 7564 9648
rect 6687 9608 7564 9636
rect 6687 9605 6699 9608
rect 6641 9599 6699 9605
rect 7558 9596 7564 9608
rect 7616 9596 7622 9648
rect 14182 9636 14188 9648
rect 11532 9608 14188 9636
rect 7374 9568 7380 9580
rect 5092 9540 7380 9568
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3651 9472 3985 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4120 9472 4445 9500
rect 4120 9460 4126 9472
rect 4433 9469 4445 9472
rect 4479 9500 4491 9503
rect 4522 9500 4528 9512
rect 4479 9472 4528 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4522 9460 4528 9472
rect 4580 9460 4586 9512
rect 4706 9500 4712 9512
rect 4667 9472 4712 9500
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 5092 9509 5120 9540
rect 7374 9528 7380 9540
rect 7432 9568 7438 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 7432 9540 9597 9568
rect 7432 9528 7438 9540
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 7101 9503 7159 9509
rect 7101 9469 7113 9503
rect 7147 9500 7159 9503
rect 7190 9500 7196 9512
rect 7147 9472 7196 9500
rect 7147 9469 7159 9472
rect 7101 9463 7159 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7558 9500 7564 9512
rect 7519 9472 7564 9500
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 8220 9509 8248 9540
rect 9585 9537 9597 9540
rect 9631 9568 9643 9571
rect 11532 9568 11560 9608
rect 14182 9596 14188 9608
rect 14240 9596 14246 9648
rect 16298 9596 16304 9648
rect 16356 9636 16362 9648
rect 16945 9639 17003 9645
rect 16945 9636 16957 9639
rect 16356 9608 16957 9636
rect 16356 9596 16362 9608
rect 16945 9605 16957 9608
rect 16991 9636 17003 9639
rect 18138 9636 18144 9648
rect 16991 9608 18144 9636
rect 16991 9605 17003 9608
rect 16945 9599 17003 9605
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 20533 9639 20591 9645
rect 20533 9605 20545 9639
rect 20579 9636 20591 9639
rect 21266 9636 21272 9648
rect 20579 9608 21272 9636
rect 20579 9605 20591 9608
rect 20533 9599 20591 9605
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 9631 9540 11560 9568
rect 9631 9537 9643 9540
rect 9585 9531 9643 9537
rect 11532 9512 11560 9540
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12768 9540 12909 9568
rect 12768 9528 12774 9540
rect 12897 9537 12909 9540
rect 12943 9568 12955 9571
rect 14090 9568 14096 9580
rect 12943 9540 14096 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 14642 9568 14648 9580
rect 14603 9540 14648 9568
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9568 15623 9571
rect 16022 9568 16028 9580
rect 15611 9540 16028 9568
rect 15611 9537 15623 9540
rect 15565 9531 15623 9537
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 19337 9571 19395 9577
rect 19337 9537 19349 9571
rect 19383 9568 19395 9571
rect 19978 9568 19984 9580
rect 19383 9540 19984 9568
rect 19383 9537 19395 9540
rect 19337 9531 19395 9537
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 20993 9571 21051 9577
rect 20993 9537 21005 9571
rect 21039 9568 21051 9571
rect 21082 9568 21088 9580
rect 21039 9540 21088 9568
rect 21039 9537 21051 9540
rect 20993 9531 21051 9537
rect 21082 9528 21088 9540
rect 21140 9568 21146 9580
rect 21453 9571 21511 9577
rect 21453 9568 21465 9571
rect 21140 9540 21465 9568
rect 21140 9528 21146 9540
rect 21453 9537 21465 9540
rect 21499 9537 21511 9571
rect 21453 9531 21511 9537
rect 21818 9528 21824 9580
rect 21876 9568 21882 9580
rect 23290 9568 23296 9580
rect 21876 9540 23296 9568
rect 21876 9528 21882 9540
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9469 8263 9503
rect 9214 9500 9220 9512
rect 9127 9472 9220 9500
rect 8205 9463 8263 9469
rect 4724 9432 4752 9460
rect 2924 9404 4752 9432
rect 2924 9392 2930 9404
rect 6638 9392 6644 9444
rect 6696 9432 6702 9444
rect 7852 9432 7880 9463
rect 9214 9460 9220 9472
rect 9272 9500 9278 9512
rect 9950 9500 9956 9512
rect 9272 9472 9956 9500
rect 9272 9460 9278 9472
rect 9950 9460 9956 9472
rect 10008 9500 10014 9512
rect 10318 9500 10324 9512
rect 10008 9472 10324 9500
rect 10008 9460 10014 9472
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 10594 9500 10600 9512
rect 10555 9472 10600 9500
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10870 9500 10876 9512
rect 10831 9472 10876 9500
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 11425 9503 11483 9509
rect 11425 9469 11437 9503
rect 11471 9500 11483 9503
rect 11514 9500 11520 9512
rect 11471 9472 11520 9500
rect 11471 9469 11483 9472
rect 11425 9463 11483 9469
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 11882 9500 11888 9512
rect 11843 9472 11888 9500
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 13780 9472 14565 9500
rect 13780 9460 13786 9472
rect 14553 9469 14565 9472
rect 14599 9500 14611 9503
rect 14921 9503 14979 9509
rect 14921 9500 14933 9503
rect 14599 9472 14933 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 14921 9469 14933 9472
rect 14967 9469 14979 9503
rect 21545 9503 21603 9509
rect 21545 9500 21557 9503
rect 14921 9463 14979 9469
rect 21284 9472 21557 9500
rect 8573 9435 8631 9441
rect 8573 9432 8585 9435
rect 6696 9404 8585 9432
rect 6696 9392 6702 9404
rect 8573 9401 8585 9404
rect 8619 9401 8631 9435
rect 8573 9395 8631 9401
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3568 9336 3801 9364
rect 3568 9324 3574 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 6914 9364 6920 9376
rect 6875 9336 6920 9364
rect 3789 9327 3847 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 7616 9336 9965 9364
rect 7616 9324 7622 9336
rect 9953 9333 9965 9336
rect 9999 9364 10011 9367
rect 10134 9364 10140 9376
rect 9999 9336 10140 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10134 9324 10140 9336
rect 10192 9364 10198 9376
rect 10612 9364 10640 9460
rect 10888 9432 10916 9460
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 10888 9404 12173 9432
rect 12161 9401 12173 9404
rect 12207 9432 12219 9435
rect 12342 9432 12348 9444
rect 12207 9404 12348 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 12342 9392 12348 9404
rect 12400 9392 12406 9444
rect 15657 9435 15715 9441
rect 15657 9401 15669 9435
rect 15703 9401 15715 9435
rect 15657 9395 15715 9401
rect 16209 9435 16267 9441
rect 16209 9401 16221 9435
rect 16255 9432 16267 9435
rect 17310 9432 17316 9444
rect 16255 9404 17316 9432
rect 16255 9401 16267 9404
rect 16209 9395 16267 9401
rect 10192 9336 10640 9364
rect 10192 9324 10198 9336
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 10836 9336 11253 9364
rect 10836 9324 10842 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 12434 9364 12440 9376
rect 12395 9336 12440 9364
rect 11241 9327 11299 9333
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 15381 9367 15439 9373
rect 15381 9333 15393 9367
rect 15427 9364 15439 9367
rect 15672 9364 15700 9395
rect 17310 9392 17316 9404
rect 17368 9432 17374 9444
rect 18141 9435 18199 9441
rect 18141 9432 18153 9435
rect 17368 9404 18153 9432
rect 17368 9392 17374 9404
rect 18141 9401 18153 9404
rect 18187 9401 18199 9435
rect 18141 9395 18199 9401
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 18233 9395 18291 9401
rect 18785 9435 18843 9441
rect 18785 9401 18797 9435
rect 18831 9432 18843 9435
rect 18966 9432 18972 9444
rect 18831 9404 18972 9432
rect 18831 9401 18843 9404
rect 18785 9395 18843 9401
rect 16114 9364 16120 9376
rect 15427 9336 16120 9364
rect 15427 9333 15439 9336
rect 15381 9327 15439 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 17770 9324 17776 9336
rect 17828 9364 17834 9376
rect 18248 9364 18276 9395
rect 18966 9392 18972 9404
rect 19024 9392 19030 9444
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 19978 9432 19984 9444
rect 19576 9404 19984 9432
rect 19576 9392 19582 9404
rect 19978 9392 19984 9404
rect 20036 9432 20042 9444
rect 21284 9441 21312 9472
rect 21545 9469 21557 9472
rect 21591 9469 21603 9503
rect 24581 9503 24639 9509
rect 24581 9500 24593 9503
rect 21545 9463 21603 9469
rect 24412 9472 24593 9500
rect 20073 9435 20131 9441
rect 20073 9432 20085 9435
rect 20036 9404 20085 9432
rect 20036 9392 20042 9404
rect 20073 9401 20085 9404
rect 20119 9432 20131 9435
rect 21269 9435 21327 9441
rect 21269 9432 21281 9435
rect 20119 9404 21281 9432
rect 20119 9401 20131 9404
rect 20073 9395 20131 9401
rect 21269 9401 21281 9404
rect 21315 9401 21327 9435
rect 21269 9395 21327 9401
rect 24412 9376 24440 9472
rect 24581 9469 24593 9472
rect 24627 9469 24639 9503
rect 24581 9463 24639 9469
rect 17828 9336 18276 9364
rect 17828 9324 17834 9336
rect 19426 9324 19432 9376
rect 19484 9364 19490 9376
rect 19613 9367 19671 9373
rect 19613 9364 19625 9367
rect 19484 9336 19625 9364
rect 19484 9324 19490 9336
rect 19613 9333 19625 9336
rect 19659 9333 19671 9367
rect 24394 9364 24400 9376
rect 24355 9336 24400 9364
rect 19613 9327 19671 9333
rect 24394 9324 24400 9336
rect 24452 9324 24458 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 3786 9160 3792 9172
rect 3747 9132 3792 9160
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 6273 9163 6331 9169
rect 4212 9132 4257 9160
rect 4212 9120 4218 9132
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 6638 9160 6644 9172
rect 6319 9132 6644 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7926 9120 7932 9172
rect 7984 9160 7990 9172
rect 8389 9163 8447 9169
rect 8389 9160 8401 9163
rect 7984 9132 8401 9160
rect 7984 9120 7990 9132
rect 8389 9129 8401 9132
rect 8435 9160 8447 9163
rect 8711 9163 8769 9169
rect 8711 9160 8723 9163
rect 8435 9132 8723 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 8711 9129 8723 9132
rect 8757 9129 8769 9163
rect 8711 9123 8769 9129
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 9364 9132 9413 9160
rect 9364 9120 9370 9132
rect 9401 9129 9413 9132
rect 9447 9160 9459 9163
rect 9769 9163 9827 9169
rect 9769 9160 9781 9163
rect 9447 9132 9781 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 9769 9129 9781 9132
rect 9815 9129 9827 9163
rect 12342 9160 12348 9172
rect 12303 9132 12348 9160
rect 9769 9123 9827 9129
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 12802 9160 12808 9172
rect 12763 9132 12808 9160
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 15562 9120 15568 9172
rect 15620 9160 15626 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 15620 9132 15669 9160
rect 15620 9120 15626 9132
rect 15657 9129 15669 9132
rect 15703 9129 15715 9163
rect 15657 9123 15715 9129
rect 16209 9163 16267 9169
rect 16209 9129 16221 9163
rect 16255 9160 16267 9163
rect 17770 9160 17776 9172
rect 16255 9132 17776 9160
rect 16255 9129 16267 9132
rect 16209 9123 16267 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 19978 9160 19984 9172
rect 19939 9132 19984 9160
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 23707 9163 23765 9169
rect 23707 9129 23719 9163
rect 23753 9160 23765 9163
rect 24394 9160 24400 9172
rect 23753 9132 24400 9160
rect 23753 9129 23765 9132
rect 23707 9123 23765 9129
rect 24394 9120 24400 9132
rect 24452 9120 24458 9172
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3970 9092 3976 9104
rect 3191 9064 3976 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3970 9052 3976 9064
rect 4028 9092 4034 9104
rect 4028 9064 5948 9092
rect 4028 9052 4034 9064
rect 1464 9027 1522 9033
rect 1464 8993 1476 9027
rect 1510 9024 1522 9027
rect 1578 9024 1584 9036
rect 1510 8996 1584 9024
rect 1510 8993 1522 8996
rect 1464 8987 1522 8993
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 9024 3111 9027
rect 4246 9024 4252 9036
rect 3099 8996 4252 9024
rect 3099 8993 3111 8996
rect 3053 8987 3111 8993
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 4614 9024 4620 9036
rect 4575 8996 4620 9024
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 4893 9027 4951 9033
rect 4893 9024 4905 9027
rect 4764 8996 4905 9024
rect 4764 8984 4770 8996
rect 4893 8993 4905 8996
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 5261 9027 5319 9033
rect 5261 8993 5273 9027
rect 5307 9024 5319 9027
rect 5350 9024 5356 9036
rect 5307 8996 5356 9024
rect 5307 8993 5319 8996
rect 5261 8987 5319 8993
rect 3786 8916 3792 8968
rect 3844 8956 3850 8968
rect 5276 8956 5304 8987
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 5920 8965 5948 9064
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 7146 9095 7204 9101
rect 7146 9092 7158 9095
rect 6788 9064 7158 9092
rect 6788 9052 6794 9064
rect 7146 9061 7158 9064
rect 7192 9092 7204 9095
rect 7466 9092 7472 9104
rect 7192 9064 7472 9092
rect 7192 9061 7204 9064
rect 7146 9055 7204 9061
rect 7466 9052 7472 9064
rect 7524 9052 7530 9104
rect 8018 9092 8024 9104
rect 7979 9064 8024 9092
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 11882 9092 11888 9104
rect 8655 9064 11888 9092
rect 8655 9036 8683 9064
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 9024 6883 9027
rect 6914 9024 6920 9036
rect 6871 8996 6920 9024
rect 6871 8993 6883 8996
rect 6825 8987 6883 8993
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 8655 9033 8668 9036
rect 8640 9027 8668 9033
rect 8640 9024 8652 9027
rect 8575 8996 8652 9024
rect 8640 8993 8652 8996
rect 8640 8987 8668 8993
rect 8662 8984 8668 8987
rect 8720 8984 8726 9036
rect 9950 9024 9956 9036
rect 9911 8996 9956 9024
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 10134 9024 10140 9036
rect 10095 8996 10140 9024
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10686 9024 10692 9036
rect 10647 8996 10692 9024
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 10962 9024 10968 9036
rect 10923 8996 10968 9024
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 12820 9024 12848 9120
rect 17218 9092 17224 9104
rect 17179 9064 17224 9092
rect 17218 9052 17224 9064
rect 17276 9052 17282 9104
rect 18414 9052 18420 9104
rect 18472 9092 18478 9104
rect 18693 9095 18751 9101
rect 18693 9092 18705 9095
rect 18472 9064 18705 9092
rect 18472 9052 18478 9064
rect 18693 9061 18705 9064
rect 18739 9061 18751 9095
rect 18693 9055 18751 9061
rect 18785 9095 18843 9101
rect 18785 9061 18797 9095
rect 18831 9092 18843 9095
rect 19058 9092 19064 9104
rect 18831 9064 19064 9092
rect 18831 9061 18843 9064
rect 18785 9055 18843 9061
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 12897 9027 12955 9033
rect 12897 9024 12909 9027
rect 12820 8996 12909 9024
rect 12897 8993 12909 8996
rect 12943 8993 12955 9027
rect 12897 8987 12955 8993
rect 12986 8984 12992 9036
rect 13044 9024 13050 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 13044 8996 13369 9024
rect 13044 8984 13050 8996
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13722 9024 13728 9036
rect 13683 8996 13728 9024
rect 13357 8987 13415 8993
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 14182 9024 14188 9036
rect 14143 8996 14188 9024
rect 14182 8984 14188 8996
rect 14240 8984 14246 9036
rect 23636 9027 23694 9033
rect 23636 8993 23648 9027
rect 23682 9024 23694 9027
rect 23750 9024 23756 9036
rect 23682 8996 23756 9024
rect 23682 8993 23694 8996
rect 23636 8987 23694 8993
rect 23750 8984 23756 8996
rect 23808 8984 23814 9036
rect 24581 9027 24639 9033
rect 24581 8993 24593 9027
rect 24627 9024 24639 9027
rect 24670 9024 24676 9036
rect 24627 8996 24676 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 24670 8984 24676 8996
rect 24728 8984 24734 9036
rect 3844 8928 5304 8956
rect 5905 8959 5963 8965
rect 3844 8916 3850 8928
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 7190 8956 7196 8968
rect 5951 8928 7196 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 14369 8959 14427 8965
rect 14369 8925 14381 8959
rect 14415 8956 14427 8959
rect 14826 8956 14832 8968
rect 14415 8928 14832 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 14826 8916 14832 8928
rect 14884 8956 14890 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14884 8928 15301 8956
rect 14884 8916 14890 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 17126 8956 17132 8968
rect 17087 8928 17132 8956
rect 15289 8919 15347 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 17368 8928 17417 8956
rect 17368 8916 17374 8928
rect 17405 8925 17417 8928
rect 17451 8956 17463 8959
rect 18417 8959 18475 8965
rect 18417 8956 18429 8959
rect 17451 8928 18429 8956
rect 17451 8925 17463 8928
rect 17405 8919 17463 8925
rect 18417 8925 18429 8928
rect 18463 8925 18475 8959
rect 18966 8956 18972 8968
rect 18927 8928 18972 8956
rect 18417 8919 18475 8925
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 1302 8848 1308 8900
rect 1360 8888 1366 8900
rect 1857 8891 1915 8897
rect 1857 8888 1869 8891
rect 1360 8860 1869 8888
rect 1360 8848 1366 8860
rect 1857 8857 1869 8860
rect 1903 8857 1915 8891
rect 1857 8851 1915 8857
rect 20990 8848 20996 8900
rect 21048 8888 21054 8900
rect 21177 8891 21235 8897
rect 21177 8888 21189 8891
rect 21048 8860 21189 8888
rect 21048 8848 21054 8860
rect 21177 8857 21189 8860
rect 21223 8888 21235 8891
rect 24719 8891 24777 8897
rect 24719 8888 24731 8891
rect 21223 8860 24731 8888
rect 21223 8857 21235 8860
rect 21177 8851 21235 8857
rect 24719 8857 24731 8860
rect 24765 8857 24777 8891
rect 24719 8851 24777 8857
rect 1535 8823 1593 8829
rect 1535 8789 1547 8823
rect 1581 8820 1593 8823
rect 1762 8820 1768 8832
rect 1581 8792 1768 8820
rect 1581 8789 1593 8792
rect 1535 8783 1593 8789
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 7742 8820 7748 8832
rect 7703 8792 7748 8820
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 11422 8820 11428 8832
rect 11383 8792 11428 8820
rect 11422 8780 11428 8792
rect 11480 8780 11486 8832
rect 18046 8820 18052 8832
rect 18007 8792 18052 8820
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 22278 8820 22284 8832
rect 18932 8792 22284 8820
rect 18932 8780 18938 8792
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 1854 8576 1860 8628
rect 1912 8616 1918 8628
rect 1949 8619 2007 8625
rect 1949 8616 1961 8619
rect 1912 8588 1961 8616
rect 1912 8576 1918 8588
rect 1949 8585 1961 8588
rect 1995 8585 2007 8619
rect 1949 8579 2007 8585
rect 3237 8619 3295 8625
rect 3237 8585 3249 8619
rect 3283 8616 3295 8619
rect 3789 8619 3847 8625
rect 3789 8616 3801 8619
rect 3283 8588 3801 8616
rect 3283 8585 3295 8588
rect 3237 8579 3295 8585
rect 3789 8585 3801 8588
rect 3835 8616 3847 8619
rect 4246 8616 4252 8628
rect 3835 8588 4252 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 4614 8576 4620 8628
rect 4672 8616 4678 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 4672 8588 5825 8616
rect 4672 8576 4678 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 8662 8616 8668 8628
rect 8623 8588 8668 8616
rect 5813 8579 5871 8585
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 9217 8619 9275 8625
rect 9217 8585 9229 8619
rect 9263 8616 9275 8619
rect 10134 8616 10140 8628
rect 9263 8588 10140 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10744 8588 10885 8616
rect 10744 8576 10750 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12986 8616 12992 8628
rect 12299 8588 12992 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13078 8576 13084 8628
rect 13136 8616 13142 8628
rect 15105 8619 15163 8625
rect 15105 8616 15117 8619
rect 13136 8588 15117 8616
rect 13136 8576 13142 8588
rect 15105 8585 15117 8588
rect 15151 8616 15163 8619
rect 15562 8616 15568 8628
rect 15151 8588 15568 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 16114 8616 16120 8628
rect 16075 8588 16120 8616
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 24670 8616 24676 8628
rect 24631 8588 24676 8616
rect 24670 8576 24676 8588
rect 24728 8576 24734 8628
rect 1762 8508 1768 8560
rect 1820 8548 1826 8560
rect 7469 8551 7527 8557
rect 1820 8520 6960 8548
rect 1820 8508 1826 8520
rect 2314 8480 2320 8492
rect 2148 8452 2320 8480
rect 2148 8421 2176 8452
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 2866 8480 2872 8492
rect 2827 8452 2872 8480
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 6932 8489 6960 8520
rect 7469 8517 7481 8551
rect 7515 8548 7527 8551
rect 8202 8548 8208 8560
rect 7515 8520 8208 8548
rect 7515 8517 7527 8520
rect 7469 8511 7527 8517
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 10505 8551 10563 8557
rect 10505 8548 10517 8551
rect 9548 8520 10517 8548
rect 9548 8508 9554 8520
rect 10505 8517 10517 8520
rect 10551 8548 10563 8551
rect 10962 8548 10968 8560
rect 10551 8520 10968 8548
rect 10551 8517 10563 8520
rect 10505 8511 10563 8517
rect 10962 8508 10968 8520
rect 11020 8548 11026 8560
rect 12710 8548 12716 8560
rect 11020 8520 12716 8548
rect 11020 8508 11026 8520
rect 12710 8508 12716 8520
rect 12768 8508 12774 8560
rect 12802 8508 12808 8560
rect 12860 8548 12866 8560
rect 14645 8551 14703 8557
rect 14645 8548 14657 8551
rect 12860 8520 14657 8548
rect 12860 8508 12866 8520
rect 14645 8517 14657 8520
rect 14691 8517 14703 8551
rect 15580 8548 15608 8576
rect 16393 8551 16451 8557
rect 16393 8548 16405 8551
rect 15580 8520 16405 8548
rect 14645 8511 14703 8517
rect 16393 8517 16405 8520
rect 16439 8517 16451 8551
rect 18046 8548 18052 8560
rect 16393 8511 16451 8517
rect 17011 8520 18052 8548
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 3568 8452 4261 8480
rect 3568 8440 3574 8452
rect 4249 8449 4261 8452
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8480 6975 8483
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 6963 8452 7849 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 9306 8480 9312 8492
rect 9267 8452 9312 8480
rect 7837 8443 7895 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 12342 8440 12348 8492
rect 12400 8480 12406 8492
rect 12400 8452 13768 8480
rect 12400 8440 12406 8452
rect 13740 8424 13768 8452
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 17011 8480 17039 8520
rect 18046 8508 18052 8520
rect 18104 8548 18110 8560
rect 18877 8551 18935 8557
rect 18104 8520 18184 8548
rect 18104 8508 18110 8520
rect 18156 8489 18184 8520
rect 18877 8517 18889 8551
rect 18923 8548 18935 8551
rect 21818 8548 21824 8560
rect 18923 8520 21824 8548
rect 18923 8517 18935 8520
rect 18877 8511 18935 8517
rect 21818 8508 21824 8520
rect 21876 8508 21882 8560
rect 15528 8452 17039 8480
rect 18141 8483 18199 8489
rect 15528 8440 15534 8452
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18414 8480 18420 8492
rect 18375 8452 18420 8480
rect 18141 8443 18199 8449
rect 18414 8440 18420 8452
rect 18472 8480 18478 8492
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 18472 8452 19441 8480
rect 18472 8440 18478 8452
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8381 2191 8415
rect 2133 8375 2191 8381
rect 2222 8372 2228 8424
rect 2280 8412 2286 8424
rect 2409 8415 2467 8421
rect 2280 8384 2325 8412
rect 2280 8372 2286 8384
rect 2409 8381 2421 8415
rect 2455 8381 2467 8415
rect 2409 8375 2467 8381
rect 11124 8415 11182 8421
rect 11124 8381 11136 8415
rect 11170 8412 11182 8415
rect 11170 8384 11652 8412
rect 11170 8381 11182 8384
rect 11124 8375 11182 8381
rect 1854 8304 1860 8356
rect 1912 8344 1918 8356
rect 2424 8344 2452 8375
rect 5445 8347 5503 8353
rect 5445 8344 5457 8347
rect 1912 8316 2452 8344
rect 4632 8316 5457 8344
rect 1912 8304 1918 8316
rect 4632 8288 4660 8316
rect 5445 8313 5457 8316
rect 5491 8313 5503 8347
rect 5445 8307 5503 8313
rect 6273 8347 6331 8353
rect 6273 8313 6285 8347
rect 6319 8344 6331 8347
rect 7009 8347 7067 8353
rect 7009 8344 7021 8347
rect 6319 8316 7021 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 7009 8313 7021 8316
rect 7055 8344 7067 8347
rect 7098 8344 7104 8356
rect 7055 8316 7104 8344
rect 7055 8313 7067 8316
rect 7009 8307 7067 8313
rect 3786 8236 3792 8288
rect 3844 8276 3850 8288
rect 4065 8279 4123 8285
rect 4065 8276 4077 8279
rect 3844 8248 4077 8276
rect 3844 8236 3850 8248
rect 4065 8245 4077 8248
rect 4111 8245 4123 8279
rect 4614 8276 4620 8288
rect 4575 8248 4620 8276
rect 4065 8239 4123 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 5166 8276 5172 8288
rect 5127 8248 5172 8276
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 5460 8276 5488 8307
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 9582 8344 9588 8356
rect 9543 8316 9588 8344
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 11624 8344 11652 8384
rect 12802 8372 12808 8424
rect 12860 8412 12866 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12860 8384 12909 8412
rect 12860 8372 12866 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 12986 8372 12992 8424
rect 13044 8412 13050 8424
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 13044 8384 13369 8412
rect 13044 8372 13050 8384
rect 13357 8381 13369 8384
rect 13403 8412 13415 8415
rect 13538 8412 13544 8424
rect 13403 8384 13544 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 13722 8412 13728 8424
rect 13635 8384 13728 8412
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 14090 8412 14096 8424
rect 14051 8384 14096 8412
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14369 8415 14427 8421
rect 14369 8381 14381 8415
rect 14415 8412 14427 8415
rect 15194 8412 15200 8424
rect 14415 8384 15200 8412
rect 14415 8381 14427 8384
rect 14369 8375 14427 8381
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 15930 8412 15936 8424
rect 15396 8384 15936 8412
rect 15396 8344 15424 8384
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 16942 8412 16948 8424
rect 16903 8384 16948 8412
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 17218 8372 17224 8424
rect 17276 8412 17282 8424
rect 17313 8415 17371 8421
rect 17313 8412 17325 8415
rect 17276 8384 17325 8412
rect 17276 8372 17282 8384
rect 17313 8381 17325 8384
rect 17359 8412 17371 8415
rect 17773 8415 17831 8421
rect 17773 8412 17785 8415
rect 17359 8384 17785 8412
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 17773 8381 17785 8384
rect 17819 8381 17831 8415
rect 17773 8375 17831 8381
rect 17126 8353 17132 8356
rect 17083 8347 17132 8353
rect 17083 8344 17095 8347
rect 11624 8316 15424 8344
rect 17039 8316 17095 8344
rect 11624 8288 11652 8316
rect 17083 8313 17095 8316
rect 17129 8313 17132 8347
rect 17083 8307 17132 8313
rect 17126 8304 17132 8307
rect 17184 8344 17190 8356
rect 17494 8344 17500 8356
rect 17184 8316 17500 8344
rect 17184 8304 17190 8316
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 17788 8344 17816 8375
rect 18233 8347 18291 8353
rect 18233 8344 18245 8347
rect 17788 8316 18245 8344
rect 18233 8313 18245 8316
rect 18279 8313 18291 8347
rect 18233 8307 18291 8313
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 5460 8248 6561 8276
rect 6549 8245 6561 8248
rect 6595 8276 6607 8279
rect 6730 8276 6736 8288
rect 6595 8248 6736 8276
rect 6595 8245 6607 8248
rect 6549 8239 6607 8245
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 10229 8279 10287 8285
rect 10229 8276 10241 8279
rect 10100 8248 10241 8276
rect 10100 8236 10106 8248
rect 10229 8245 10241 8248
rect 10275 8245 10287 8279
rect 10229 8239 10287 8245
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 11195 8279 11253 8285
rect 11195 8276 11207 8279
rect 11020 8248 11207 8276
rect 11020 8236 11026 8248
rect 11195 8245 11207 8248
rect 11241 8245 11253 8279
rect 11606 8276 11612 8288
rect 11567 8248 11612 8276
rect 11195 8239 11253 8245
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 15562 8276 15568 8288
rect 15523 8248 15568 8276
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 16574 8236 16580 8288
rect 16632 8276 16638 8288
rect 16761 8279 16819 8285
rect 16761 8276 16773 8279
rect 16632 8248 16773 8276
rect 16632 8236 16638 8248
rect 16761 8245 16773 8248
rect 16807 8276 16819 8279
rect 17313 8279 17371 8285
rect 17313 8276 17325 8279
rect 16807 8248 17325 8276
rect 16807 8245 16819 8248
rect 16761 8239 16819 8245
rect 17313 8245 17325 8248
rect 17359 8245 17371 8279
rect 17313 8239 17371 8245
rect 17405 8279 17463 8285
rect 17405 8245 17417 8279
rect 17451 8276 17463 8279
rect 17586 8276 17592 8288
rect 17451 8248 17592 8276
rect 17451 8245 17463 8248
rect 17405 8239 17463 8245
rect 17586 8236 17592 8248
rect 17644 8276 17650 8288
rect 18877 8279 18935 8285
rect 18877 8276 18889 8279
rect 17644 8248 18889 8276
rect 17644 8236 17650 8248
rect 18877 8245 18889 8248
rect 18923 8245 18935 8279
rect 19058 8276 19064 8288
rect 19019 8248 19064 8276
rect 18877 8239 18935 8245
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 23750 8236 23756 8288
rect 23808 8276 23814 8288
rect 23845 8279 23903 8285
rect 23845 8276 23857 8279
rect 23808 8248 23857 8276
rect 23808 8236 23814 8248
rect 23845 8245 23857 8248
rect 23891 8245 23903 8279
rect 23845 8239 23903 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 1670 8072 1676 8084
rect 1627 8044 1676 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 2222 8072 2228 8084
rect 2183 8044 2228 8072
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 3510 8072 3516 8084
rect 3471 8044 3516 8072
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 4614 8072 4620 8084
rect 4575 8044 4620 8072
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 6972 8044 7297 8072
rect 6972 8032 6978 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 7524 8044 9321 8072
rect 7524 8032 7530 8044
rect 9309 8041 9321 8044
rect 9355 8072 9367 8075
rect 9582 8072 9588 8084
rect 9355 8044 9588 8072
rect 9355 8041 9367 8044
rect 9309 8035 9367 8041
rect 9582 8032 9588 8044
rect 9640 8072 9646 8084
rect 9640 8032 9674 8072
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 10008 8044 10149 8072
rect 10008 8032 10014 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8072 10655 8075
rect 10962 8072 10968 8084
rect 10643 8044 10968 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11146 8072 11152 8084
rect 11107 8044 11152 8072
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 11572 8044 12357 8072
rect 11572 8032 11578 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 13538 8072 13544 8084
rect 13499 8044 13544 8072
rect 12345 8035 12403 8041
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 15933 8075 15991 8081
rect 15933 8072 15945 8075
rect 15252 8044 15945 8072
rect 15252 8032 15258 8044
rect 15933 8041 15945 8044
rect 15979 8041 15991 8075
rect 17494 8072 17500 8084
rect 17455 8044 17500 8072
rect 15933 8035 15991 8041
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 2866 7964 2872 8016
rect 2924 8004 2930 8016
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 2924 7976 3801 8004
rect 2924 7964 2930 7976
rect 3789 7973 3801 7976
rect 3835 7973 3847 8007
rect 7742 8004 7748 8016
rect 3789 7967 3847 7973
rect 6932 7976 7748 8004
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 2222 7936 2228 7948
rect 1443 7908 2228 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 2406 7936 2412 7948
rect 2367 7908 2412 7936
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 6932 7945 6960 7976
rect 7742 7964 7748 7976
rect 7800 8004 7806 8016
rect 8021 8007 8079 8013
rect 8021 8004 8033 8007
rect 7800 7976 8033 8004
rect 7800 7964 7806 7976
rect 8021 7973 8033 7976
rect 8067 7973 8079 8007
rect 9646 8004 9674 8032
rect 11164 8004 11192 8032
rect 9646 7976 11192 8004
rect 8021 7967 8079 7973
rect 12434 7964 12440 8016
rect 12492 8004 12498 8016
rect 12621 8007 12679 8013
rect 12621 8004 12633 8007
rect 12492 7976 12633 8004
rect 12492 7964 12498 7976
rect 12621 7973 12633 7976
rect 12667 7973 12679 8007
rect 12621 7967 12679 7973
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 15470 8004 15476 8016
rect 12768 7976 12813 8004
rect 15431 7976 15476 8004
rect 12768 7964 12774 7976
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 16114 7964 16120 8016
rect 16172 8004 16178 8016
rect 16669 8007 16727 8013
rect 16669 8004 16681 8007
rect 16172 7976 16681 8004
rect 16172 7964 16178 7976
rect 16669 7973 16681 7976
rect 16715 7973 16727 8007
rect 16669 7967 16727 7973
rect 17221 8007 17279 8013
rect 17221 7973 17233 8007
rect 17267 8004 17279 8007
rect 18414 8004 18420 8016
rect 17267 7976 18420 8004
rect 17267 7973 17279 7976
rect 17221 7967 17279 7973
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 18785 8007 18843 8013
rect 18785 7973 18797 8007
rect 18831 8004 18843 8007
rect 19058 8004 19064 8016
rect 18831 7976 19064 8004
rect 18831 7973 18843 7976
rect 18785 7967 18843 7973
rect 19058 7964 19064 7976
rect 19116 7964 19122 8016
rect 4249 7939 4307 7945
rect 4249 7936 4261 7939
rect 4212 7908 4261 7936
rect 4212 7896 4218 7908
rect 4249 7905 4261 7908
rect 4295 7905 4307 7939
rect 4249 7899 4307 7905
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 9712 7939 9770 7945
rect 9712 7936 9724 7939
rect 9640 7908 9724 7936
rect 9640 7896 9646 7908
rect 9712 7905 9724 7908
rect 9758 7905 9770 7939
rect 9712 7899 9770 7905
rect 9815 7939 9873 7945
rect 9815 7905 9827 7939
rect 9861 7936 9873 7939
rect 12069 7939 12127 7945
rect 9861 7908 11145 7936
rect 9861 7905 9873 7908
rect 9815 7899 9873 7905
rect 7006 7868 7012 7880
rect 6967 7840 7012 7868
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8202 7868 8208 7880
rect 7975 7840 8208 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 10778 7868 10784 7880
rect 10739 7840 10784 7868
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 11117 7868 11145 7908
rect 12069 7905 12081 7939
rect 12115 7936 12127 7939
rect 12342 7936 12348 7948
rect 12115 7908 12348 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 17770 7896 17776 7948
rect 17828 7936 17834 7948
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 17828 7908 18153 7936
rect 17828 7896 17834 7908
rect 18141 7905 18153 7908
rect 18187 7936 18199 7939
rect 18230 7936 18236 7948
rect 18187 7908 18236 7936
rect 18187 7905 18199 7908
rect 18141 7899 18199 7905
rect 18230 7896 18236 7908
rect 18288 7896 18294 7948
rect 23198 7896 23204 7948
rect 23256 7936 23262 7948
rect 24581 7939 24639 7945
rect 24581 7936 24593 7939
rect 23256 7908 24593 7936
rect 23256 7896 23262 7908
rect 24581 7905 24593 7908
rect 24627 7936 24639 7939
rect 24670 7936 24676 7948
rect 24627 7908 24676 7936
rect 24627 7905 24639 7908
rect 24581 7899 24639 7905
rect 24670 7896 24676 7908
rect 24728 7896 24734 7948
rect 16390 7868 16396 7880
rect 11117 7840 16396 7868
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 17310 7868 17316 7880
rect 16623 7840 17316 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 17310 7828 17316 7840
rect 17368 7828 17374 7880
rect 8478 7800 8484 7812
rect 8439 7772 8484 7800
rect 8478 7760 8484 7772
rect 8536 7760 8542 7812
rect 12158 7760 12164 7812
rect 12216 7800 12222 7812
rect 13173 7803 13231 7809
rect 13173 7800 13185 7803
rect 12216 7772 13185 7800
rect 12216 7760 12222 7772
rect 13173 7769 13185 7772
rect 13219 7800 13231 7803
rect 13446 7800 13452 7812
rect 13219 7772 13452 7800
rect 13219 7769 13231 7772
rect 13173 7763 13231 7769
rect 13446 7760 13452 7772
rect 13504 7760 13510 7812
rect 2222 7692 2228 7744
rect 2280 7732 2286 7744
rect 2639 7735 2697 7741
rect 2639 7732 2651 7735
rect 2280 7704 2651 7732
rect 2280 7692 2286 7704
rect 2639 7701 2651 7704
rect 2685 7701 2697 7735
rect 2639 7695 2697 7701
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 5169 7735 5227 7741
rect 5169 7732 5181 7735
rect 4856 7704 5181 7732
rect 4856 7692 4862 7704
rect 5169 7701 5181 7704
rect 5215 7701 5227 7735
rect 5169 7695 5227 7701
rect 5258 7692 5264 7744
rect 5316 7732 5322 7744
rect 5445 7735 5503 7741
rect 5445 7732 5457 7735
rect 5316 7704 5457 7732
rect 5316 7692 5322 7704
rect 5445 7701 5457 7704
rect 5491 7701 5503 7735
rect 11698 7732 11704 7744
rect 11659 7704 11704 7732
rect 5445 7695 5503 7701
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 24765 7735 24823 7741
rect 24765 7701 24777 7735
rect 24811 7732 24823 7735
rect 27614 7732 27620 7744
rect 24811 7704 27620 7732
rect 24811 7701 24823 7704
rect 24765 7695 24823 7701
rect 27614 7692 27620 7704
rect 27672 7692 27678 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1673 7531 1731 7537
rect 1673 7497 1685 7531
rect 1719 7528 1731 7531
rect 2222 7528 2228 7540
rect 1719 7500 2228 7528
rect 1719 7497 1731 7500
rect 1673 7491 1731 7497
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7064 7500 7849 7528
rect 7064 7488 7070 7500
rect 7837 7497 7849 7500
rect 7883 7528 7895 7531
rect 8202 7528 8208 7540
rect 7883 7500 8208 7528
rect 7883 7497 7895 7500
rect 7837 7491 7895 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 10042 7528 10048 7540
rect 10003 7500 10048 7528
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 11146 7528 11152 7540
rect 11059 7500 11152 7528
rect 11146 7488 11152 7500
rect 11204 7528 11210 7540
rect 13078 7528 13084 7540
rect 11204 7500 13084 7528
rect 11204 7488 11210 7500
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 15749 7531 15807 7537
rect 15749 7497 15761 7531
rect 15795 7528 15807 7531
rect 16114 7528 16120 7540
rect 15795 7500 16120 7528
rect 15795 7497 15807 7500
rect 15749 7491 15807 7497
rect 16114 7488 16120 7500
rect 16172 7528 16178 7540
rect 16853 7531 16911 7537
rect 16853 7528 16865 7531
rect 16172 7500 16865 7528
rect 16172 7488 16178 7500
rect 16853 7497 16865 7500
rect 16899 7497 16911 7531
rect 18230 7528 18236 7540
rect 18191 7500 18236 7528
rect 16853 7491 16911 7497
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 24670 7528 24676 7540
rect 24631 7500 24676 7528
rect 24670 7488 24676 7500
rect 24728 7488 24734 7540
rect 2406 7420 2412 7472
rect 2464 7460 2470 7472
rect 2593 7463 2651 7469
rect 2593 7460 2605 7463
rect 2464 7432 2605 7460
rect 2464 7420 2470 7432
rect 2593 7429 2605 7432
rect 2639 7460 2651 7463
rect 6365 7463 6423 7469
rect 2639 7432 5488 7460
rect 2639 7429 2651 7432
rect 2593 7423 2651 7429
rect 5460 7404 5488 7432
rect 6365 7429 6377 7463
rect 6411 7460 6423 7463
rect 7561 7463 7619 7469
rect 7561 7460 7573 7463
rect 6411 7432 7573 7460
rect 6411 7429 6423 7432
rect 6365 7423 6423 7429
rect 7561 7429 7573 7432
rect 7607 7460 7619 7463
rect 7742 7460 7748 7472
rect 7607 7432 7748 7460
rect 7607 7429 7619 7432
rect 7561 7423 7619 7429
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5258 7392 5264 7404
rect 5215 7364 5264 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5442 7392 5448 7404
rect 5355 7364 5448 7392
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 8478 7392 8484 7404
rect 8439 7364 8484 7392
rect 8478 7352 8484 7364
rect 8536 7392 8542 7404
rect 9582 7392 9588 7404
rect 8536 7364 9588 7392
rect 8536 7352 8542 7364
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7392 10287 7395
rect 10962 7392 10968 7404
rect 10275 7364 10968 7392
rect 10275 7361 10287 7364
rect 10229 7355 10287 7361
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7392 12311 7395
rect 12437 7395 12495 7401
rect 12437 7392 12449 7395
rect 12299 7364 12449 7392
rect 12299 7361 12311 7364
rect 12253 7355 12311 7361
rect 12437 7361 12449 7364
rect 12483 7392 12495 7395
rect 12710 7392 12716 7404
rect 12483 7364 12716 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 16574 7392 16580 7404
rect 16535 7364 16580 7392
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 3421 7327 3479 7333
rect 3421 7293 3433 7327
rect 3467 7324 3479 7327
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 3467 7296 4169 7324
rect 3467 7293 3479 7296
rect 3421 7287 3479 7293
rect 4157 7293 4169 7296
rect 4203 7324 4215 7327
rect 4798 7324 4804 7336
rect 4203 7296 4804 7324
rect 4203 7293 4215 7296
rect 4157 7287 4215 7293
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 11756 7296 11897 7324
rect 11756 7284 11762 7296
rect 11885 7293 11897 7296
rect 11931 7324 11943 7327
rect 12529 7327 12587 7333
rect 12529 7324 12541 7327
rect 11931 7296 12541 7324
rect 11931 7293 11943 7296
rect 11885 7287 11943 7293
rect 12529 7293 12541 7296
rect 12575 7293 12587 7327
rect 16114 7324 16120 7336
rect 16075 7296 16120 7324
rect 12529 7287 12587 7293
rect 16114 7284 16120 7296
rect 16172 7284 16178 7336
rect 4246 7256 4252 7268
rect 4207 7228 4252 7256
rect 4246 7216 4252 7228
rect 4304 7216 4310 7268
rect 5261 7259 5319 7265
rect 5261 7225 5273 7259
rect 5307 7225 5319 7259
rect 5261 7219 5319 7225
rect 7009 7259 7067 7265
rect 7009 7225 7021 7259
rect 7055 7256 7067 7259
rect 8110 7256 8116 7268
rect 7055 7228 8116 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 2372 7160 4537 7188
rect 2372 7148 2378 7160
rect 4525 7157 4537 7160
rect 4571 7188 4583 7191
rect 4614 7188 4620 7200
rect 4571 7160 4620 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 4890 7188 4896 7200
rect 4851 7160 4896 7188
rect 4890 7148 4896 7160
rect 4948 7188 4954 7200
rect 5276 7188 5304 7219
rect 8110 7216 8116 7228
rect 8168 7216 8174 7268
rect 8202 7216 8208 7268
rect 8260 7256 8266 7268
rect 8260 7228 8305 7256
rect 8260 7216 8266 7228
rect 10042 7216 10048 7268
rect 10100 7256 10106 7268
rect 10321 7259 10379 7265
rect 10321 7256 10333 7259
rect 10100 7228 10333 7256
rect 10100 7216 10106 7228
rect 10321 7225 10333 7228
rect 10367 7225 10379 7259
rect 10870 7256 10876 7268
rect 10831 7228 10876 7256
rect 10321 7219 10379 7225
rect 10870 7216 10876 7228
rect 10928 7216 10934 7268
rect 17310 7188 17316 7200
rect 4948 7160 5304 7188
rect 17271 7160 17316 7188
rect 4948 7148 4954 7160
rect 17310 7148 17316 7160
rect 17368 7148 17374 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 4154 6944 4160 6996
rect 4212 6984 4218 6996
rect 4249 6987 4307 6993
rect 4249 6984 4261 6987
rect 4212 6956 4261 6984
rect 4212 6944 4218 6956
rect 4249 6953 4261 6956
rect 4295 6953 4307 6987
rect 8110 6984 8116 6996
rect 8071 6956 8116 6984
rect 4249 6947 4307 6953
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8389 6987 8447 6993
rect 8389 6984 8401 6987
rect 8352 6956 8401 6984
rect 8352 6944 8358 6956
rect 8389 6953 8401 6956
rect 8435 6953 8447 6987
rect 10778 6984 10784 6996
rect 10739 6956 10784 6984
rect 8389 6947 8447 6953
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 12529 6987 12587 6993
rect 12529 6984 12541 6987
rect 12492 6956 12541 6984
rect 12492 6944 12498 6956
rect 12529 6953 12541 6956
rect 12575 6953 12587 6987
rect 12529 6947 12587 6953
rect 4798 6876 4804 6928
rect 4856 6916 4862 6928
rect 5169 6919 5227 6925
rect 5169 6916 5181 6919
rect 4856 6888 5181 6916
rect 4856 6876 4862 6888
rect 5169 6885 5181 6888
rect 5215 6885 5227 6919
rect 6730 6916 6736 6928
rect 6691 6888 6736 6916
rect 5169 6879 5227 6885
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 9950 6916 9956 6928
rect 9911 6888 9956 6916
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 11609 6919 11667 6925
rect 11609 6885 11621 6919
rect 11655 6916 11667 6919
rect 11698 6916 11704 6928
rect 11655 6888 11704 6916
rect 11655 6885 11667 6888
rect 11609 6879 11667 6885
rect 11698 6876 11704 6888
rect 11756 6876 11762 6928
rect 12158 6916 12164 6928
rect 12119 6888 12164 6916
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 24581 6851 24639 6857
rect 24581 6817 24593 6851
rect 24627 6848 24639 6851
rect 24762 6848 24768 6860
rect 24627 6820 24768 6848
rect 24627 6817 24639 6820
rect 24581 6811 24639 6817
rect 24762 6808 24768 6820
rect 24820 6808 24826 6860
rect 4522 6740 4528 6792
rect 4580 6780 4586 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4580 6752 5089 6780
rect 4580 6740 4586 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5534 6780 5540 6792
rect 5495 6752 5540 6780
rect 5077 6743 5135 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 7006 6780 7012 6792
rect 6687 6752 7012 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 9858 6780 9864 6792
rect 9819 6752 9864 6780
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 10870 6780 10876 6792
rect 10551 6752 10876 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 10870 6740 10876 6752
rect 10928 6780 10934 6792
rect 11514 6780 11520 6792
rect 10928 6752 11520 6780
rect 10928 6740 10934 6752
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 5258 6672 5264 6724
rect 5316 6712 5322 6724
rect 7193 6715 7251 6721
rect 7193 6712 7205 6715
rect 5316 6684 7205 6712
rect 5316 6672 5322 6684
rect 7193 6681 7205 6684
rect 7239 6681 7251 6715
rect 7193 6675 7251 6681
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 2958 6644 2964 6656
rect 2915 6616 2964 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3099 6647 3157 6653
rect 3099 6613 3111 6647
rect 3145 6644 3157 6647
rect 4154 6644 4160 6656
rect 3145 6616 4160 6644
rect 3145 6613 3157 6616
rect 3099 6607 3157 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 24765 6647 24823 6653
rect 24765 6613 24777 6647
rect 24811 6644 24823 6647
rect 27614 6644 27620 6656
rect 24811 6616 27620 6644
rect 24811 6613 24823 6616
rect 24765 6607 24823 6613
rect 27614 6604 27620 6616
rect 27672 6604 27678 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 4304 6412 6561 6440
rect 4304 6400 4310 6412
rect 6549 6409 6561 6412
rect 6595 6440 6607 6443
rect 6730 6440 6736 6452
rect 6595 6412 6736 6440
rect 6595 6409 6607 6412
rect 6549 6403 6607 6409
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 11514 6400 11520 6452
rect 11572 6440 11578 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11572 6412 11805 6440
rect 11572 6400 11578 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 24673 6443 24731 6449
rect 24673 6409 24685 6443
rect 24719 6440 24731 6443
rect 24762 6440 24768 6452
rect 24719 6412 24768 6440
rect 24719 6409 24731 6412
rect 24673 6403 24731 6409
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 5166 6372 5172 6384
rect 4080 6344 5172 6372
rect 4080 6245 4108 6344
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 19889 6375 19947 6381
rect 19889 6341 19901 6375
rect 19935 6372 19947 6375
rect 21358 6372 21364 6384
rect 19935 6344 21364 6372
rect 19935 6341 19947 6344
rect 19889 6335 19947 6341
rect 21358 6332 21364 6344
rect 21416 6332 21422 6384
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4890 6304 4896 6316
rect 4203 6276 4896 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 5442 6304 5448 6316
rect 5403 6276 5448 6304
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6304 9643 6307
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9631 6276 9689 6304
rect 9631 6273 9643 6276
rect 9585 6267 9643 6273
rect 9677 6273 9689 6276
rect 9723 6304 9735 6307
rect 9950 6304 9956 6316
rect 9723 6276 9956 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6304 11575 6307
rect 11698 6304 11704 6316
rect 11563 6276 11704 6304
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 9217 6239 9275 6245
rect 9217 6205 9229 6239
rect 9263 6236 9275 6239
rect 10042 6236 10048 6248
rect 9263 6208 10048 6236
rect 9263 6205 9275 6208
rect 9217 6199 9275 6205
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 16390 6196 16396 6248
rect 16448 6236 16454 6248
rect 19705 6239 19763 6245
rect 19705 6236 19717 6239
rect 16448 6208 19717 6236
rect 16448 6196 16454 6208
rect 19705 6205 19717 6208
rect 19751 6236 19763 6239
rect 20257 6239 20315 6245
rect 20257 6236 20269 6239
rect 19751 6208 20269 6236
rect 19751 6205 19763 6208
rect 19705 6199 19763 6205
rect 20257 6205 20269 6208
rect 20303 6205 20315 6239
rect 20257 6199 20315 6205
rect 5074 6168 5080 6180
rect 5035 6140 5080 6168
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 5166 6128 5172 6180
rect 5224 6168 5230 6180
rect 5224 6140 5269 6168
rect 5224 6128 5230 6140
rect 2958 6100 2964 6112
rect 2919 6072 2964 6100
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 4890 6100 4896 6112
rect 4851 6072 4896 6100
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 5092 6100 5120 6128
rect 5534 6100 5540 6112
rect 5092 6072 5540 6100
rect 5534 6060 5540 6072
rect 5592 6100 5598 6112
rect 5997 6103 6055 6109
rect 5997 6100 6009 6103
rect 5592 6072 6009 6100
rect 5592 6060 5598 6072
rect 5997 6069 6009 6072
rect 6043 6069 6055 6103
rect 7006 6100 7012 6112
rect 6967 6072 7012 6100
rect 5997 6063 6055 6069
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5896 4307 5899
rect 7006 5896 7012 5908
rect 4295 5868 7012 5896
rect 4295 5865 4307 5868
rect 4249 5859 4307 5865
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 24578 5856 24584 5908
rect 24636 5896 24642 5908
rect 24719 5899 24777 5905
rect 24719 5896 24731 5899
rect 24636 5868 24731 5896
rect 24636 5856 24642 5868
rect 24719 5865 24731 5868
rect 24765 5865 24777 5899
rect 24719 5859 24777 5865
rect 3513 5831 3571 5837
rect 3513 5797 3525 5831
rect 3559 5828 3571 5831
rect 5077 5831 5135 5837
rect 5077 5828 5089 5831
rect 3559 5800 5089 5828
rect 3559 5797 3571 5800
rect 3513 5791 3571 5797
rect 5077 5797 5089 5800
rect 5123 5828 5135 5831
rect 5166 5828 5172 5840
rect 5123 5800 5172 5828
rect 5123 5797 5135 5800
rect 5077 5791 5135 5797
rect 5166 5788 5172 5800
rect 5224 5788 5230 5840
rect 5442 5828 5448 5840
rect 5403 5800 5448 5828
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 24648 5763 24706 5769
rect 24648 5729 24660 5763
rect 24694 5760 24706 5763
rect 25222 5760 25228 5772
rect 24694 5732 25228 5760
rect 24694 5729 24706 5732
rect 24648 5723 24706 5729
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 5350 5692 5356 5704
rect 5311 5664 5356 5692
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 5258 5584 5264 5636
rect 5316 5624 5322 5636
rect 5644 5624 5672 5655
rect 5316 5596 5672 5624
rect 5316 5584 5322 5596
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5442 5556 5448 5568
rect 4948 5528 5448 5556
rect 4948 5516 4954 5528
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 9858 5556 9864 5568
rect 8996 5528 9864 5556
rect 8996 5516 9002 5528
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4304 5324 4629 5352
rect 4304 5312 4310 5324
rect 4617 5321 4629 5324
rect 4663 5352 4675 5355
rect 4982 5352 4988 5364
rect 4663 5324 4988 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5500 5324 5825 5352
rect 5500 5312 5506 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 24762 5352 24768 5364
rect 24723 5324 24768 5352
rect 5813 5315 5871 5321
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4890 5216 4896 5228
rect 4212 5188 4896 5216
rect 4212 5176 4218 5188
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 5132 5188 5181 5216
rect 5132 5176 5138 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 24397 5151 24455 5157
rect 24397 5148 24409 5151
rect 19484 5120 24409 5148
rect 19484 5108 19490 5120
rect 24397 5117 24409 5120
rect 24443 5148 24455 5151
rect 24581 5151 24639 5157
rect 24581 5148 24593 5151
rect 24443 5120 24593 5148
rect 24443 5117 24455 5120
rect 24397 5111 24455 5117
rect 24581 5117 24593 5120
rect 24627 5117 24639 5151
rect 24581 5111 24639 5117
rect 4982 5080 4988 5092
rect 4943 5052 4988 5080
rect 4982 5040 4988 5052
rect 5040 5040 5046 5092
rect 25222 5012 25228 5024
rect 25183 4984 25228 5012
rect 25222 4972 25228 4984
rect 25280 4972 25286 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 4890 4808 4896 4820
rect 4851 4780 4896 4808
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5350 4808 5356 4820
rect 5311 4780 5356 4808
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 1210 4632 1216 4684
rect 1268 4672 1274 4684
rect 1397 4675 1455 4681
rect 1397 4672 1409 4675
rect 1268 4644 1409 4672
rect 1268 4632 1274 4644
rect 1397 4641 1409 4644
rect 1443 4672 1455 4675
rect 1670 4672 1676 4684
rect 1443 4644 1676 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1670 4632 1676 4644
rect 1728 4632 1734 4684
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 24029 4199 24087 4205
rect 24029 4165 24041 4199
rect 24075 4196 24087 4199
rect 27614 4196 27620 4208
rect 24075 4168 27620 4196
rect 24075 4165 24087 4168
rect 24029 4159 24087 4165
rect 27614 4156 27620 4168
rect 27672 4156 27678 4208
rect 1670 4060 1676 4072
rect 1631 4032 1676 4060
rect 1670 4020 1676 4032
rect 1728 4020 1734 4072
rect 23842 4060 23848 4072
rect 23755 4032 23848 4060
rect 23842 4020 23848 4032
rect 23900 4060 23906 4072
rect 24397 4063 24455 4069
rect 24397 4060 24409 4063
rect 23900 4032 24409 4060
rect 23900 4020 23906 4032
rect 24397 4029 24409 4032
rect 24443 4029 24455 4063
rect 24397 4023 24455 4029
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 10459 3179 10517 3185
rect 10459 3145 10471 3179
rect 10505 3176 10517 3179
rect 11422 3176 11428 3188
rect 10505 3148 11428 3176
rect 10505 3145 10517 3148
rect 10459 3139 10517 3145
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 24719 3179 24777 3185
rect 24719 3145 24731 3179
rect 24765 3176 24777 3179
rect 24854 3176 24860 3188
rect 24765 3148 24860 3176
rect 24765 3145 24777 3148
rect 24719 3139 24777 3145
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 10388 2975 10446 2981
rect 10388 2941 10400 2975
rect 10434 2972 10446 2975
rect 24648 2975 24706 2981
rect 10434 2944 10916 2972
rect 10434 2941 10446 2944
rect 10388 2935 10446 2941
rect 10888 2848 10916 2944
rect 24648 2941 24660 2975
rect 24694 2972 24706 2975
rect 24694 2944 25176 2972
rect 24694 2941 24706 2944
rect 24648 2935 24706 2941
rect 25148 2848 25176 2944
rect 10870 2836 10876 2848
rect 10831 2808 10876 2836
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 25130 2836 25136 2848
rect 25091 2808 25136 2836
rect 25130 2796 25136 2808
rect 25188 2796 25194 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 4522 2592 4528 2644
rect 4580 2632 4586 2644
rect 5031 2635 5089 2641
rect 5031 2632 5043 2635
rect 4580 2604 5043 2632
rect 4580 2592 4586 2604
rect 5031 2601 5043 2604
rect 5077 2601 5089 2635
rect 5031 2595 5089 2601
rect 8803 2635 8861 2641
rect 8803 2601 8815 2635
rect 8849 2632 8861 2635
rect 8938 2632 8944 2644
rect 8849 2604 8944 2632
rect 8849 2601 8861 2604
rect 8803 2595 8861 2601
rect 8938 2592 8944 2604
rect 8996 2592 9002 2644
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11287 2604 13814 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 4960 2499 5018 2505
rect 4960 2465 4972 2499
rect 5006 2496 5018 2499
rect 8732 2499 8790 2505
rect 5006 2468 5488 2496
rect 5006 2465 5018 2468
rect 4960 2459 5018 2465
rect 5460 2301 5488 2468
rect 8732 2465 8744 2499
rect 8778 2496 8790 2499
rect 9122 2496 9128 2508
rect 8778 2468 9128 2496
rect 8778 2465 8790 2468
rect 8732 2459 8790 2465
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2496 10655 2499
rect 11256 2496 11284 2595
rect 13786 2564 13814 2604
rect 16390 2592 16396 2644
rect 16448 2632 16454 2644
rect 23063 2635 23121 2641
rect 23063 2632 23075 2635
rect 16448 2604 23075 2632
rect 16448 2592 16454 2604
rect 23063 2601 23075 2604
rect 23109 2601 23121 2635
rect 24719 2635 24777 2641
rect 24719 2632 24731 2635
rect 23063 2595 23121 2601
rect 23216 2604 24731 2632
rect 17862 2564 17868 2576
rect 13786 2536 17868 2564
rect 17862 2524 17868 2536
rect 17920 2524 17926 2576
rect 23216 2564 23244 2604
rect 24719 2601 24731 2604
rect 24765 2601 24777 2635
rect 24719 2595 24777 2601
rect 25406 2564 25412 2576
rect 17972 2536 23244 2564
rect 23860 2536 25412 2564
rect 10643 2468 11284 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 11388 2468 12633 2496
rect 11388 2456 11394 2468
rect 12621 2465 12633 2468
rect 12667 2496 12679 2499
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12667 2468 13185 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 13173 2459 13231 2465
rect 15470 2456 15476 2468
rect 15528 2496 15534 2508
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15528 2468 16037 2496
rect 15528 2456 15534 2468
rect 16025 2465 16037 2468
rect 16071 2465 16083 2499
rect 16025 2459 16083 2465
rect 17678 2456 17684 2508
rect 17736 2496 17742 2508
rect 17972 2496 18000 2536
rect 17736 2468 18000 2496
rect 22992 2499 23050 2505
rect 17736 2456 17742 2468
rect 22992 2465 23004 2499
rect 23038 2496 23050 2499
rect 23477 2499 23535 2505
rect 23477 2496 23489 2499
rect 23038 2468 23489 2496
rect 23038 2465 23050 2468
rect 22992 2459 23050 2465
rect 23477 2465 23489 2468
rect 23523 2496 23535 2499
rect 23860 2496 23888 2536
rect 25406 2524 25412 2536
rect 25464 2524 25470 2576
rect 23523 2468 23888 2496
rect 24648 2499 24706 2505
rect 23523 2465 23535 2468
rect 23477 2459 23535 2465
rect 24648 2465 24660 2499
rect 24694 2496 24706 2499
rect 24694 2468 25176 2496
rect 24694 2465 24706 2468
rect 24648 2459 24706 2465
rect 10781 2363 10839 2369
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 11882 2360 11888 2372
rect 10827 2332 11888 2360
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 15657 2363 15715 2369
rect 15657 2329 15669 2363
rect 15703 2360 15715 2363
rect 17126 2360 17132 2372
rect 15703 2332 17132 2360
rect 15703 2329 15715 2332
rect 15657 2323 15715 2329
rect 17126 2320 17132 2332
rect 17184 2320 17190 2372
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 5994 2292 6000 2304
rect 5491 2264 6000 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 9122 2292 9128 2304
rect 9083 2264 9128 2292
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2292 12863 2295
rect 12986 2292 12992 2304
rect 12851 2264 12992 2292
rect 12851 2261 12863 2264
rect 12805 2255 12863 2261
rect 12986 2252 12992 2264
rect 13044 2252 13050 2304
rect 25148 2301 25176 2468
rect 25133 2295 25191 2301
rect 25133 2261 25145 2295
rect 25179 2292 25191 2295
rect 26878 2292 26884 2304
rect 25179 2264 26884 2292
rect 25179 2261 25191 2264
rect 25133 2255 25191 2261
rect 26878 2252 26884 2264
rect 26936 2252 26942 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 17218 184 17224 196
rect 14660 156 17224 184
rect 14660 128 14688 156
rect 17218 144 17224 156
rect 17276 144 17282 196
rect 658 76 664 128
rect 716 116 722 128
rect 1302 116 1308 128
rect 716 88 1308 116
rect 716 76 722 88
rect 1302 76 1308 88
rect 1360 76 1366 128
rect 4246 76 4252 128
rect 4304 116 4310 128
rect 4798 116 4804 128
rect 4304 88 4804 116
rect 4304 76 4310 88
rect 4798 76 4804 88
rect 4856 76 4862 128
rect 9674 76 9680 128
rect 9732 116 9738 128
rect 10410 116 10416 128
rect 9732 88 10416 116
rect 9732 76 9738 88
rect 10410 76 10416 88
rect 10468 76 10474 128
rect 14642 76 14648 128
rect 14700 76 14706 128
rect 17954 76 17960 128
rect 18012 116 18018 128
rect 18782 116 18788 128
rect 18012 88 18788 116
rect 18012 76 18018 88
rect 18782 76 18788 88
rect 18840 76 18846 128
rect 19518 76 19524 128
rect 19576 116 19582 128
rect 20162 116 20168 128
rect 19576 88 20168 116
rect 19576 76 19582 88
rect 20162 76 20168 88
rect 20220 76 20226 128
rect 23566 76 23572 128
rect 23624 116 23630 128
rect 24394 116 24400 128
rect 23624 88 24400 116
rect 23624 76 23630 88
rect 24394 76 24400 88
rect 24452 76 24458 128
<< via1 >>
rect 3240 27480 3292 27532
rect 3976 27480 4028 27532
rect 11244 27480 11296 27532
rect 12256 27480 12308 27532
rect 26240 27480 26292 27532
rect 27068 27480 27120 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 13912 24352 13964 24404
rect 5540 24216 5592 24268
rect 13360 24259 13412 24268
rect 13360 24225 13369 24259
rect 13369 24225 13403 24259
rect 13403 24225 13412 24259
rect 13360 24216 13412 24225
rect 4620 24012 4672 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 5540 23808 5592 23860
rect 13360 23851 13412 23860
rect 13360 23817 13369 23851
rect 13369 23817 13403 23851
rect 13403 23817 13412 23851
rect 13360 23808 13412 23817
rect 15476 23808 15528 23860
rect 20444 23808 20496 23860
rect 22100 23808 22152 23860
rect 5264 23604 5316 23656
rect 18052 23647 18104 23656
rect 5724 23468 5776 23520
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 21272 23647 21324 23656
rect 21272 23613 21281 23647
rect 21281 23613 21315 23647
rect 21315 23613 21324 23647
rect 21272 23604 21324 23613
rect 14648 23468 14700 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5724 23264 5776 23316
rect 6920 23264 6972 23316
rect 13360 23264 13412 23316
rect 18052 23264 18104 23316
rect 14556 23128 14608 23180
rect 16120 23171 16172 23180
rect 16120 23137 16129 23171
rect 16129 23137 16163 23171
rect 16163 23137 16172 23171
rect 16120 23128 16172 23137
rect 25136 23128 25188 23180
rect 13176 22924 13228 22976
rect 13820 22924 13872 22976
rect 21456 22924 21508 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1860 22763 1912 22772
rect 1860 22729 1869 22763
rect 1869 22729 1903 22763
rect 1903 22729 1912 22763
rect 1860 22720 1912 22729
rect 14556 22763 14608 22772
rect 14556 22729 14565 22763
rect 14565 22729 14599 22763
rect 14599 22729 14608 22763
rect 14556 22720 14608 22729
rect 15384 22720 15436 22772
rect 21272 22720 21324 22772
rect 25504 22763 25556 22772
rect 25504 22729 25513 22763
rect 25513 22729 25547 22763
rect 25547 22729 25556 22763
rect 25504 22720 25556 22729
rect 7012 22652 7064 22704
rect 25136 22695 25188 22704
rect 25136 22661 25145 22695
rect 25145 22661 25179 22695
rect 25179 22661 25188 22695
rect 25136 22652 25188 22661
rect 27620 22652 27672 22704
rect 6920 22627 6972 22636
rect 6920 22593 6929 22627
rect 6929 22593 6963 22627
rect 6963 22593 6972 22627
rect 6920 22584 6972 22593
rect 1860 22516 1912 22568
rect 7012 22491 7064 22500
rect 7012 22457 7021 22491
rect 7021 22457 7055 22491
rect 7055 22457 7064 22491
rect 7564 22491 7616 22500
rect 7012 22448 7064 22457
rect 7564 22457 7573 22491
rect 7573 22457 7607 22491
rect 7607 22457 7616 22491
rect 7564 22448 7616 22457
rect 8576 22448 8628 22500
rect 8668 22380 8720 22432
rect 8944 22380 8996 22432
rect 9772 22380 9824 22432
rect 11060 22380 11112 22432
rect 13820 22516 13872 22568
rect 14280 22491 14332 22500
rect 14280 22457 14289 22491
rect 14289 22457 14323 22491
rect 14323 22457 14332 22491
rect 14280 22448 14332 22457
rect 25504 22516 25556 22568
rect 14832 22380 14884 22432
rect 16120 22380 16172 22432
rect 20352 22380 20404 22432
rect 21640 22380 21692 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 8944 22219 8996 22228
rect 8944 22185 8953 22219
rect 8953 22185 8987 22219
rect 8987 22185 8996 22219
rect 8944 22176 8996 22185
rect 6460 22151 6512 22160
rect 6460 22117 6469 22151
rect 6469 22117 6503 22151
rect 6503 22117 6512 22151
rect 6460 22108 6512 22117
rect 7564 22108 7616 22160
rect 8024 22151 8076 22160
rect 8024 22117 8033 22151
rect 8033 22117 8067 22151
rect 8067 22117 8076 22151
rect 8024 22108 8076 22117
rect 8668 22108 8720 22160
rect 12532 22108 12584 22160
rect 1492 22040 1544 22092
rect 9772 22083 9824 22092
rect 9772 22049 9790 22083
rect 9790 22049 9824 22083
rect 18788 22176 18840 22228
rect 21456 22219 21508 22228
rect 21456 22185 21465 22219
rect 21465 22185 21499 22219
rect 21499 22185 21508 22219
rect 21456 22176 21508 22185
rect 12992 22151 13044 22160
rect 12992 22117 13001 22151
rect 13001 22117 13035 22151
rect 13035 22117 13044 22151
rect 12992 22108 13044 22117
rect 17408 22108 17460 22160
rect 9772 22040 9824 22049
rect 19156 22040 19208 22092
rect 22376 22040 22428 22092
rect 23940 22108 23992 22160
rect 25412 22108 25464 22160
rect 24676 22083 24728 22092
rect 24676 22049 24694 22083
rect 24694 22049 24728 22083
rect 24676 22040 24728 22049
rect 25228 22040 25280 22092
rect 5540 21972 5592 22024
rect 7932 22015 7984 22024
rect 7932 21981 7941 22015
rect 7941 21981 7975 22015
rect 7975 21981 7984 22015
rect 7932 21972 7984 21981
rect 8668 21972 8720 22024
rect 12900 22015 12952 22024
rect 12900 21981 12909 22015
rect 12909 21981 12943 22015
rect 12943 21981 12952 22015
rect 12900 21972 12952 21981
rect 13820 21972 13872 22024
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 17040 22015 17092 22024
rect 10968 21904 11020 21956
rect 15844 21904 15896 21956
rect 15936 21904 15988 21956
rect 17040 21981 17049 22015
rect 17049 21981 17083 22015
rect 17083 21981 17092 22015
rect 17040 21972 17092 21981
rect 20904 22015 20956 22024
rect 20904 21981 20913 22015
rect 20913 21981 20947 22015
rect 20947 21981 20956 22015
rect 20904 21972 20956 21981
rect 5540 21836 5592 21888
rect 9956 21836 10008 21888
rect 14188 21836 14240 21888
rect 16488 21836 16540 21888
rect 22192 21836 22244 21888
rect 24032 21836 24084 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1492 21632 1544 21684
rect 5540 21675 5592 21684
rect 5540 21641 5549 21675
rect 5549 21641 5583 21675
rect 5583 21641 5592 21675
rect 5540 21632 5592 21641
rect 7012 21632 7064 21684
rect 7748 21632 7800 21684
rect 8024 21607 8076 21616
rect 8024 21573 8033 21607
rect 8033 21573 8067 21607
rect 8067 21573 8076 21607
rect 8024 21564 8076 21573
rect 4160 21360 4212 21412
rect 7104 21403 7156 21412
rect 7104 21369 7113 21403
rect 7113 21369 7147 21403
rect 7147 21369 7156 21403
rect 7104 21360 7156 21369
rect 7840 21360 7892 21412
rect 9036 21632 9088 21684
rect 12900 21632 12952 21684
rect 15936 21675 15988 21684
rect 9772 21607 9824 21616
rect 9772 21573 9781 21607
rect 9781 21573 9815 21607
rect 9815 21573 9824 21607
rect 9772 21564 9824 21573
rect 15936 21641 15945 21675
rect 15945 21641 15979 21675
rect 15979 21641 15988 21675
rect 15936 21632 15988 21641
rect 22376 21675 22428 21684
rect 22376 21641 22385 21675
rect 22385 21641 22419 21675
rect 22419 21641 22428 21675
rect 22376 21632 22428 21641
rect 23756 21632 23808 21684
rect 23940 21675 23992 21684
rect 23940 21641 23949 21675
rect 23949 21641 23983 21675
rect 23983 21641 23992 21675
rect 23940 21632 23992 21641
rect 24676 21675 24728 21684
rect 24676 21641 24685 21675
rect 24685 21641 24719 21675
rect 24719 21641 24728 21675
rect 24676 21632 24728 21641
rect 8944 21496 8996 21548
rect 12532 21539 12584 21548
rect 12532 21505 12541 21539
rect 12541 21505 12575 21539
rect 12575 21505 12584 21539
rect 12532 21496 12584 21505
rect 12900 21539 12952 21548
rect 12900 21505 12909 21539
rect 12909 21505 12943 21539
rect 12943 21505 12952 21539
rect 12900 21496 12952 21505
rect 13636 21496 13688 21548
rect 16488 21539 16540 21548
rect 10048 21471 10100 21480
rect 10048 21437 10057 21471
rect 10057 21437 10091 21471
rect 10091 21437 10100 21471
rect 10048 21428 10100 21437
rect 16488 21505 16497 21539
rect 16497 21505 16531 21539
rect 16531 21505 16540 21539
rect 16488 21496 16540 21505
rect 17040 21564 17092 21616
rect 17132 21496 17184 21548
rect 19156 21539 19208 21548
rect 9220 21403 9272 21412
rect 9220 21369 9229 21403
rect 9229 21369 9263 21403
rect 9263 21369 9272 21403
rect 9220 21360 9272 21369
rect 6460 21292 6512 21344
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 14188 21360 14240 21412
rect 15292 21360 15344 21412
rect 12256 21292 12308 21301
rect 12808 21292 12860 21344
rect 12992 21292 13044 21344
rect 15936 21292 15988 21344
rect 16856 21360 16908 21412
rect 18144 21428 18196 21480
rect 19156 21505 19165 21539
rect 19165 21505 19199 21539
rect 19199 21505 19208 21539
rect 19156 21496 19208 21505
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 21548 21496 21600 21548
rect 18788 21403 18840 21412
rect 18788 21369 18797 21403
rect 18797 21369 18831 21403
rect 18831 21369 18840 21403
rect 18788 21360 18840 21369
rect 17408 21335 17460 21344
rect 17408 21301 17417 21335
rect 17417 21301 17451 21335
rect 17451 21301 17460 21335
rect 17408 21292 17460 21301
rect 19984 21292 20036 21344
rect 20628 21292 20680 21344
rect 22836 21292 22888 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 7012 21088 7064 21140
rect 10048 21088 10100 21140
rect 6368 21020 6420 21072
rect 6644 21063 6696 21072
rect 6644 21029 6653 21063
rect 6653 21029 6687 21063
rect 6687 21029 6696 21063
rect 6644 21020 6696 21029
rect 16488 21131 16540 21140
rect 16488 21097 16497 21131
rect 16497 21097 16531 21131
rect 16531 21097 16540 21131
rect 16488 21088 16540 21097
rect 18788 21088 18840 21140
rect 22192 21131 22244 21140
rect 22192 21097 22201 21131
rect 22201 21097 22235 21131
rect 22235 21097 22244 21131
rect 22192 21088 22244 21097
rect 12256 21063 12308 21072
rect 12256 21029 12265 21063
rect 12265 21029 12299 21063
rect 12299 21029 12308 21063
rect 12256 21020 12308 21029
rect 7380 20952 7432 21004
rect 8484 20952 8536 21004
rect 10692 20995 10744 21004
rect 10692 20961 10701 20995
rect 10701 20961 10735 20995
rect 10735 20961 10744 20995
rect 10692 20952 10744 20961
rect 11060 20995 11112 21004
rect 11060 20961 11069 20995
rect 11069 20961 11103 20995
rect 11103 20961 11112 20995
rect 11060 20952 11112 20961
rect 12900 21020 12952 21072
rect 13360 21020 13412 21072
rect 16764 21063 16816 21072
rect 16764 21029 16773 21063
rect 16773 21029 16807 21063
rect 16807 21029 16816 21063
rect 16764 21020 16816 21029
rect 17408 21020 17460 21072
rect 19524 21020 19576 21072
rect 20904 21020 20956 21072
rect 21364 21020 21416 21072
rect 22836 21063 22888 21072
rect 22836 21029 22845 21063
rect 22845 21029 22879 21063
rect 22879 21029 22888 21063
rect 22836 21020 22888 21029
rect 14648 20952 14700 21004
rect 18236 20995 18288 21004
rect 18236 20961 18245 20995
rect 18245 20961 18279 20995
rect 18279 20961 18288 20995
rect 18236 20952 18288 20961
rect 25504 20952 25556 21004
rect 12348 20884 12400 20936
rect 13452 20884 13504 20936
rect 13728 20927 13780 20936
rect 13728 20893 13737 20927
rect 13737 20893 13771 20927
rect 13771 20893 13780 20927
rect 13728 20884 13780 20893
rect 16672 20927 16724 20936
rect 16672 20893 16681 20927
rect 16681 20893 16715 20927
rect 16715 20893 16724 20927
rect 16672 20884 16724 20893
rect 14096 20816 14148 20868
rect 17592 20884 17644 20936
rect 19984 20884 20036 20936
rect 21456 20927 21508 20936
rect 21456 20893 21465 20927
rect 21465 20893 21499 20927
rect 21499 20893 21508 20927
rect 21456 20884 21508 20893
rect 22744 20927 22796 20936
rect 22744 20893 22753 20927
rect 22753 20893 22787 20927
rect 22787 20893 22796 20927
rect 22744 20884 22796 20893
rect 19800 20816 19852 20868
rect 20812 20816 20864 20868
rect 22008 20816 22060 20868
rect 5540 20748 5592 20800
rect 6184 20791 6236 20800
rect 6184 20757 6193 20791
rect 6193 20757 6227 20791
rect 6227 20757 6236 20791
rect 6184 20748 6236 20757
rect 7288 20791 7340 20800
rect 7288 20757 7297 20791
rect 7297 20757 7331 20791
rect 7331 20757 7340 20791
rect 7288 20748 7340 20757
rect 7932 20791 7984 20800
rect 7932 20757 7941 20791
rect 7941 20757 7975 20791
rect 7975 20757 7984 20791
rect 7932 20748 7984 20757
rect 15660 20748 15712 20800
rect 18052 20791 18104 20800
rect 18052 20757 18061 20791
rect 18061 20757 18095 20791
rect 18095 20757 18104 20791
rect 18052 20748 18104 20757
rect 18696 20791 18748 20800
rect 18696 20757 18705 20791
rect 18705 20757 18739 20791
rect 18739 20757 18748 20791
rect 18696 20748 18748 20757
rect 18880 20748 18932 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 7288 20544 7340 20596
rect 8760 20544 8812 20596
rect 13360 20587 13412 20596
rect 13360 20553 13369 20587
rect 13369 20553 13403 20587
rect 13403 20553 13412 20587
rect 13360 20544 13412 20553
rect 14648 20544 14700 20596
rect 16672 20544 16724 20596
rect 20904 20544 20956 20596
rect 22744 20544 22796 20596
rect 23388 20587 23440 20596
rect 23388 20553 23397 20587
rect 23397 20553 23431 20587
rect 23431 20553 23440 20587
rect 23388 20544 23440 20553
rect 25136 20587 25188 20596
rect 25136 20553 25145 20587
rect 25145 20553 25179 20587
rect 25179 20553 25188 20587
rect 25136 20544 25188 20553
rect 25504 20587 25556 20596
rect 25504 20553 25513 20587
rect 25513 20553 25547 20587
rect 25547 20553 25556 20587
rect 25504 20544 25556 20553
rect 7748 20519 7800 20528
rect 7748 20485 7757 20519
rect 7757 20485 7791 20519
rect 7791 20485 7800 20519
rect 7748 20476 7800 20485
rect 4160 20451 4212 20460
rect 4160 20417 4169 20451
rect 4169 20417 4203 20451
rect 4203 20417 4212 20451
rect 4160 20408 4212 20417
rect 6184 20408 6236 20460
rect 8852 20408 8904 20460
rect 3884 20272 3936 20324
rect 5540 20340 5592 20392
rect 7656 20340 7708 20392
rect 6644 20315 6696 20324
rect 6644 20281 6653 20315
rect 6653 20281 6687 20315
rect 6687 20281 6696 20315
rect 6644 20272 6696 20281
rect 7288 20272 7340 20324
rect 8668 20315 8720 20324
rect 8668 20281 8677 20315
rect 8677 20281 8711 20315
rect 8711 20281 8720 20315
rect 8668 20272 8720 20281
rect 8760 20315 8812 20324
rect 8760 20281 8769 20315
rect 8769 20281 8803 20315
rect 8803 20281 8812 20315
rect 8760 20272 8812 20281
rect 2044 20247 2096 20256
rect 2044 20213 2053 20247
rect 2053 20213 2087 20247
rect 2087 20213 2096 20247
rect 2044 20204 2096 20213
rect 6368 20204 6420 20256
rect 7472 20204 7524 20256
rect 10692 20408 10744 20460
rect 12256 20408 12308 20460
rect 11060 20383 11112 20392
rect 11060 20349 11069 20383
rect 11069 20349 11103 20383
rect 11103 20349 11112 20383
rect 11060 20340 11112 20349
rect 12440 20383 12492 20392
rect 10784 20272 10836 20324
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 12440 20340 12492 20349
rect 12624 20272 12676 20324
rect 12900 20408 12952 20460
rect 15292 20408 15344 20460
rect 21548 20476 21600 20528
rect 16764 20408 16816 20460
rect 17132 20408 17184 20460
rect 18788 20408 18840 20460
rect 19800 20408 19852 20460
rect 20536 20451 20588 20460
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 20812 20451 20864 20460
rect 20812 20417 20821 20451
rect 20821 20417 20855 20451
rect 20855 20417 20864 20451
rect 20812 20408 20864 20417
rect 22192 20408 22244 20460
rect 22836 20476 22888 20528
rect 17408 20383 17460 20392
rect 17408 20349 17417 20383
rect 17417 20349 17451 20383
rect 17451 20349 17460 20383
rect 17408 20340 17460 20349
rect 10692 20204 10744 20256
rect 11980 20204 12032 20256
rect 12256 20247 12308 20256
rect 12256 20213 12265 20247
rect 12265 20213 12299 20247
rect 12299 20213 12308 20247
rect 12256 20204 12308 20213
rect 13728 20272 13780 20324
rect 15660 20272 15712 20324
rect 18696 20272 18748 20324
rect 25136 20340 25188 20392
rect 20628 20315 20680 20324
rect 20628 20281 20637 20315
rect 20637 20281 20671 20315
rect 20671 20281 20680 20315
rect 20628 20272 20680 20281
rect 22284 20272 22336 20324
rect 14464 20204 14516 20256
rect 15844 20204 15896 20256
rect 17316 20204 17368 20256
rect 18236 20247 18288 20256
rect 18236 20213 18245 20247
rect 18245 20213 18279 20247
rect 18279 20213 18288 20247
rect 18236 20204 18288 20213
rect 19524 20204 19576 20256
rect 21364 20204 21416 20256
rect 23112 20204 23164 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 7656 20043 7708 20052
rect 7656 20009 7665 20043
rect 7665 20009 7699 20043
rect 7699 20009 7708 20043
rect 7656 20000 7708 20009
rect 8484 20000 8536 20052
rect 1952 19864 2004 19916
rect 4988 19864 5040 19916
rect 7748 19932 7800 19984
rect 8668 20000 8720 20052
rect 12164 20000 12216 20052
rect 12808 20043 12860 20052
rect 12808 20009 12817 20043
rect 12817 20009 12851 20043
rect 12851 20009 12860 20043
rect 12808 20000 12860 20009
rect 13728 20000 13780 20052
rect 15292 20000 15344 20052
rect 16672 20000 16724 20052
rect 19524 20043 19576 20052
rect 19524 20009 19533 20043
rect 19533 20009 19567 20043
rect 19567 20009 19576 20043
rect 19524 20000 19576 20009
rect 19984 20000 20036 20052
rect 20536 20043 20588 20052
rect 20536 20009 20545 20043
rect 20545 20009 20579 20043
rect 20579 20009 20588 20043
rect 20536 20000 20588 20009
rect 23388 20000 23440 20052
rect 11980 19932 12032 19984
rect 13912 19932 13964 19984
rect 15476 19932 15528 19984
rect 15660 19932 15712 19984
rect 16028 19932 16080 19984
rect 16764 19932 16816 19984
rect 17224 19975 17276 19984
rect 17224 19941 17233 19975
rect 17233 19941 17267 19975
rect 17267 19941 17276 19975
rect 17224 19932 17276 19941
rect 18696 19932 18748 19984
rect 21364 19932 21416 19984
rect 22100 19932 22152 19984
rect 7288 19864 7340 19916
rect 7932 19864 7984 19916
rect 10324 19907 10376 19916
rect 6000 19796 6052 19848
rect 7196 19796 7248 19848
rect 10324 19873 10333 19907
rect 10333 19873 10367 19907
rect 10367 19873 10376 19907
rect 10324 19864 10376 19873
rect 10784 19864 10836 19916
rect 4068 19728 4120 19780
rect 7104 19728 7156 19780
rect 8392 19728 8444 19780
rect 13544 19864 13596 19916
rect 22008 19907 22060 19916
rect 22008 19873 22017 19907
rect 22017 19873 22051 19907
rect 22051 19873 22060 19907
rect 22836 19907 22888 19916
rect 22008 19864 22060 19873
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 24216 19864 24268 19916
rect 11888 19839 11940 19848
rect 11888 19805 11897 19839
rect 11897 19805 11931 19839
rect 11931 19805 11940 19839
rect 11888 19796 11940 19805
rect 13452 19796 13504 19848
rect 14004 19796 14056 19848
rect 15292 19839 15344 19848
rect 15292 19805 15301 19839
rect 15301 19805 15335 19839
rect 15335 19805 15344 19839
rect 15292 19796 15344 19805
rect 17500 19796 17552 19848
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 18604 19839 18656 19848
rect 17592 19796 17644 19805
rect 18604 19805 18613 19839
rect 18613 19805 18647 19839
rect 18647 19805 18656 19839
rect 18604 19796 18656 19805
rect 20628 19796 20680 19848
rect 23112 19796 23164 19848
rect 11336 19728 11388 19780
rect 3608 19703 3660 19712
rect 3608 19669 3617 19703
rect 3617 19669 3651 19703
rect 3651 19669 3660 19703
rect 3608 19660 3660 19669
rect 5448 19660 5500 19712
rect 5540 19660 5592 19712
rect 11520 19660 11572 19712
rect 12440 19660 12492 19712
rect 14188 19728 14240 19780
rect 14740 19728 14792 19780
rect 18880 19728 18932 19780
rect 13728 19660 13780 19712
rect 15936 19660 15988 19712
rect 19340 19660 19392 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2044 19456 2096 19508
rect 3976 19320 4028 19372
rect 4988 19456 5040 19508
rect 8208 19456 8260 19508
rect 10324 19499 10376 19508
rect 10324 19465 10333 19499
rect 10333 19465 10367 19499
rect 10367 19465 10376 19499
rect 10324 19456 10376 19465
rect 11704 19456 11756 19508
rect 13820 19456 13872 19508
rect 14464 19456 14516 19508
rect 15476 19456 15528 19508
rect 15568 19456 15620 19508
rect 6276 19388 6328 19440
rect 6000 19320 6052 19372
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 7840 19363 7892 19372
rect 7840 19329 7849 19363
rect 7849 19329 7883 19363
rect 7883 19329 7892 19363
rect 7840 19320 7892 19329
rect 8300 19320 8352 19372
rect 9220 19363 9272 19372
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 1676 19252 1728 19304
rect 3424 19252 3476 19304
rect 3608 19295 3660 19304
rect 3608 19261 3617 19295
rect 3617 19261 3651 19295
rect 3651 19261 3660 19295
rect 3608 19252 3660 19261
rect 3700 19295 3752 19304
rect 3700 19261 3709 19295
rect 3709 19261 3743 19295
rect 3743 19261 3752 19295
rect 3700 19252 3752 19261
rect 4068 19252 4120 19304
rect 5172 19295 5224 19304
rect 5172 19261 5181 19295
rect 5181 19261 5215 19295
rect 5215 19261 5224 19295
rect 5172 19252 5224 19261
rect 5264 19252 5316 19304
rect 5540 19252 5592 19304
rect 7196 19252 7248 19304
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 11336 19295 11388 19304
rect 11336 19261 11345 19295
rect 11345 19261 11379 19295
rect 11379 19261 11388 19295
rect 11336 19252 11388 19261
rect 12256 19252 12308 19304
rect 15936 19456 15988 19508
rect 17224 19456 17276 19508
rect 18604 19456 18656 19508
rect 20628 19499 20680 19508
rect 20628 19465 20637 19499
rect 20637 19465 20671 19499
rect 20671 19465 20680 19499
rect 20628 19456 20680 19465
rect 22100 19499 22152 19508
rect 22100 19465 22109 19499
rect 22109 19465 22143 19499
rect 22143 19465 22152 19499
rect 22100 19456 22152 19465
rect 17408 19388 17460 19440
rect 24216 19388 24268 19440
rect 4344 19227 4396 19236
rect 112 19116 164 19168
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 3056 19116 3108 19168
rect 4344 19193 4353 19227
rect 4353 19193 4387 19227
rect 4387 19193 4396 19227
rect 4344 19184 4396 19193
rect 7748 19184 7800 19236
rect 8944 19227 8996 19236
rect 8944 19193 8953 19227
rect 8953 19193 8987 19227
rect 8987 19193 8996 19227
rect 8944 19184 8996 19193
rect 12716 19227 12768 19236
rect 6460 19116 6512 19168
rect 7288 19116 7340 19168
rect 7932 19116 7984 19168
rect 8392 19116 8444 19168
rect 12716 19193 12725 19227
rect 12725 19193 12759 19227
rect 12759 19193 12768 19227
rect 12716 19184 12768 19193
rect 12164 19159 12216 19168
rect 12164 19125 12173 19159
rect 12173 19125 12207 19159
rect 12207 19125 12216 19159
rect 12164 19116 12216 19125
rect 14096 19184 14148 19236
rect 16028 19227 16080 19236
rect 16028 19193 16037 19227
rect 16037 19193 16071 19227
rect 16071 19193 16080 19227
rect 16028 19184 16080 19193
rect 16580 19227 16632 19236
rect 16580 19193 16589 19227
rect 16589 19193 16623 19227
rect 16623 19193 16632 19227
rect 16580 19184 16632 19193
rect 15476 19116 15528 19168
rect 18696 19320 18748 19372
rect 19984 19320 20036 19372
rect 22008 19320 22060 19372
rect 18696 19184 18748 19236
rect 21272 19227 21324 19236
rect 21272 19193 21281 19227
rect 21281 19193 21315 19227
rect 21315 19193 21324 19227
rect 21272 19184 21324 19193
rect 22008 19184 22060 19236
rect 17500 19159 17552 19168
rect 17500 19125 17509 19159
rect 17509 19125 17543 19159
rect 17543 19125 17552 19159
rect 17500 19116 17552 19125
rect 18236 19159 18288 19168
rect 18236 19125 18245 19159
rect 18245 19125 18279 19159
rect 18279 19125 18288 19159
rect 18236 19116 18288 19125
rect 19432 19116 19484 19168
rect 20536 19116 20588 19168
rect 22836 19159 22888 19168
rect 22836 19125 22845 19159
rect 22845 19125 22879 19159
rect 22879 19125 22888 19159
rect 22836 19116 22888 19125
rect 24216 19116 24268 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1676 18955 1728 18964
rect 1676 18921 1685 18955
rect 1685 18921 1719 18955
rect 1719 18921 1728 18955
rect 1676 18912 1728 18921
rect 7380 18912 7432 18964
rect 8944 18955 8996 18964
rect 8944 18921 8953 18955
rect 8953 18921 8987 18955
rect 8987 18921 8996 18955
rect 8944 18912 8996 18921
rect 11888 18955 11940 18964
rect 11888 18921 11897 18955
rect 11897 18921 11931 18955
rect 11931 18921 11940 18955
rect 11888 18912 11940 18921
rect 12164 18912 12216 18964
rect 6460 18844 6512 18896
rect 12256 18844 12308 18896
rect 12716 18912 12768 18964
rect 13544 18912 13596 18964
rect 14004 18955 14056 18964
rect 14004 18921 14013 18955
rect 14013 18921 14047 18955
rect 14047 18921 14056 18955
rect 14004 18912 14056 18921
rect 14096 18844 14148 18896
rect 15936 18887 15988 18896
rect 15936 18853 15945 18887
rect 15945 18853 15979 18887
rect 15979 18853 15988 18887
rect 15936 18844 15988 18853
rect 16580 18912 16632 18964
rect 18696 18912 18748 18964
rect 18604 18844 18656 18896
rect 19432 18887 19484 18896
rect 19432 18853 19441 18887
rect 19441 18853 19475 18887
rect 19475 18853 19484 18887
rect 19432 18844 19484 18853
rect 19984 18887 20036 18896
rect 19984 18853 19993 18887
rect 19993 18853 20027 18887
rect 20027 18853 20036 18887
rect 19984 18844 20036 18853
rect 22192 18844 22244 18896
rect 22284 18844 22336 18896
rect 23112 18887 23164 18896
rect 23112 18853 23121 18887
rect 23121 18853 23155 18887
rect 23155 18853 23164 18887
rect 23112 18844 23164 18853
rect 2964 18819 3016 18828
rect 2964 18785 2973 18819
rect 2973 18785 3007 18819
rect 3007 18785 3016 18819
rect 2964 18776 3016 18785
rect 4896 18819 4948 18828
rect 4896 18785 4905 18819
rect 4905 18785 4939 18819
rect 4939 18785 4948 18819
rect 4896 18776 4948 18785
rect 4988 18776 5040 18828
rect 5264 18819 5316 18828
rect 5264 18785 5273 18819
rect 5273 18785 5307 18819
rect 5307 18785 5316 18819
rect 5264 18776 5316 18785
rect 5356 18776 5408 18828
rect 8024 18776 8076 18828
rect 8116 18819 8168 18828
rect 8116 18785 8125 18819
rect 8125 18785 8159 18819
rect 8159 18785 8168 18819
rect 10784 18819 10836 18828
rect 8116 18776 8168 18785
rect 10784 18785 10793 18819
rect 10793 18785 10827 18819
rect 10827 18785 10836 18819
rect 10784 18776 10836 18785
rect 11336 18776 11388 18828
rect 14372 18776 14424 18828
rect 17684 18819 17736 18828
rect 17684 18785 17693 18819
rect 17693 18785 17727 18819
rect 17727 18785 17736 18819
rect 17684 18776 17736 18785
rect 17960 18776 18012 18828
rect 12532 18708 12584 18760
rect 19340 18751 19392 18760
rect 19340 18717 19349 18751
rect 19349 18717 19383 18751
rect 19383 18717 19392 18751
rect 19340 18708 19392 18717
rect 20720 18708 20772 18760
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 22652 18708 22704 18760
rect 20812 18640 20864 18692
rect 22008 18683 22060 18692
rect 1768 18572 1820 18624
rect 2228 18572 2280 18624
rect 2688 18615 2740 18624
rect 2688 18581 2697 18615
rect 2697 18581 2731 18615
rect 2731 18581 2740 18615
rect 2688 18572 2740 18581
rect 3700 18615 3752 18624
rect 3700 18581 3709 18615
rect 3709 18581 3743 18615
rect 3743 18581 3752 18615
rect 3700 18572 3752 18581
rect 7380 18572 7432 18624
rect 15292 18572 15344 18624
rect 16488 18572 16540 18624
rect 21180 18615 21232 18624
rect 21180 18581 21189 18615
rect 21189 18581 21223 18615
rect 21223 18581 21232 18615
rect 21180 18572 21232 18581
rect 22008 18649 22017 18683
rect 22017 18649 22051 18683
rect 22051 18649 22060 18683
rect 22008 18640 22060 18649
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2780 18368 2832 18420
rect 3976 18368 4028 18420
rect 8944 18368 8996 18420
rect 10140 18368 10192 18420
rect 13636 18368 13688 18420
rect 14372 18368 14424 18420
rect 15936 18411 15988 18420
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 16856 18368 16908 18420
rect 17500 18368 17552 18420
rect 18696 18368 18748 18420
rect 19064 18411 19116 18420
rect 19064 18377 19073 18411
rect 19073 18377 19107 18411
rect 19107 18377 19116 18411
rect 19064 18368 19116 18377
rect 21272 18368 21324 18420
rect 23112 18368 23164 18420
rect 3148 18300 3200 18352
rect 4436 18300 4488 18352
rect 3424 18275 3476 18284
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 3424 18232 3476 18241
rect 3516 18232 3568 18284
rect 5540 18232 5592 18284
rect 7840 18232 7892 18284
rect 3148 18139 3200 18148
rect 3148 18105 3157 18139
rect 3157 18105 3191 18139
rect 3191 18105 3200 18139
rect 3148 18096 3200 18105
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 2964 18071 3016 18080
rect 2964 18037 2973 18071
rect 2973 18037 3007 18071
rect 3007 18037 3016 18071
rect 3792 18096 3844 18148
rect 4988 18096 5040 18148
rect 5356 18139 5408 18148
rect 5356 18105 5365 18139
rect 5365 18105 5399 18139
rect 5399 18105 5408 18139
rect 5356 18096 5408 18105
rect 7104 18139 7156 18148
rect 7104 18105 7113 18139
rect 7113 18105 7147 18139
rect 7147 18105 7156 18139
rect 7104 18096 7156 18105
rect 11336 18300 11388 18352
rect 13268 18300 13320 18352
rect 13728 18300 13780 18352
rect 16396 18300 16448 18352
rect 20536 18343 20588 18352
rect 20536 18309 20545 18343
rect 20545 18309 20579 18343
rect 20579 18309 20588 18343
rect 20536 18300 20588 18309
rect 22284 18300 22336 18352
rect 9956 18232 10008 18284
rect 12532 18232 12584 18284
rect 10692 18164 10744 18216
rect 11704 18164 11756 18216
rect 12072 18164 12124 18216
rect 12716 18164 12768 18216
rect 8852 18096 8904 18148
rect 9588 18139 9640 18148
rect 9588 18105 9597 18139
rect 9597 18105 9631 18139
rect 9631 18105 9640 18139
rect 9588 18096 9640 18105
rect 10784 18139 10836 18148
rect 10784 18105 10793 18139
rect 10793 18105 10827 18139
rect 10827 18105 10836 18139
rect 10784 18096 10836 18105
rect 13176 18096 13228 18148
rect 14924 18139 14976 18148
rect 14924 18105 14933 18139
rect 14933 18105 14967 18139
rect 14967 18105 14976 18139
rect 14924 18096 14976 18105
rect 4896 18071 4948 18080
rect 2964 18028 3016 18037
rect 4896 18037 4905 18071
rect 4905 18037 4939 18071
rect 4939 18037 4948 18071
rect 4896 18028 4948 18037
rect 6276 18028 6328 18080
rect 6460 18071 6512 18080
rect 6460 18037 6469 18071
rect 6469 18037 6503 18071
rect 6503 18037 6512 18071
rect 6460 18028 6512 18037
rect 7748 18028 7800 18080
rect 8116 18071 8168 18080
rect 8116 18037 8125 18071
rect 8125 18037 8159 18071
rect 8159 18037 8168 18071
rect 8116 18028 8168 18037
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 12164 18028 12216 18037
rect 12532 18071 12584 18080
rect 12532 18037 12541 18071
rect 12541 18037 12575 18071
rect 12575 18037 12584 18071
rect 12532 18028 12584 18037
rect 13268 18028 13320 18080
rect 13544 18028 13596 18080
rect 14372 18028 14424 18080
rect 14648 18071 14700 18080
rect 14648 18037 14657 18071
rect 14657 18037 14691 18071
rect 14691 18037 14700 18071
rect 15384 18096 15436 18148
rect 15660 18096 15712 18148
rect 16764 18164 16816 18216
rect 17776 18232 17828 18284
rect 19248 18207 19300 18216
rect 17684 18139 17736 18148
rect 17684 18105 17693 18139
rect 17693 18105 17727 18139
rect 17727 18105 17736 18139
rect 17684 18096 17736 18105
rect 16488 18071 16540 18080
rect 14648 18028 14700 18037
rect 16488 18037 16497 18071
rect 16497 18037 16531 18071
rect 16531 18037 16540 18071
rect 16488 18028 16540 18037
rect 19248 18173 19257 18207
rect 19257 18173 19291 18207
rect 19291 18173 19300 18207
rect 19248 18164 19300 18173
rect 21180 18164 21232 18216
rect 22560 18164 22612 18216
rect 19064 18096 19116 18148
rect 24032 18164 24084 18216
rect 18696 18028 18748 18080
rect 21088 18028 21140 18080
rect 22192 18071 22244 18080
rect 22192 18037 22201 18071
rect 22201 18037 22235 18071
rect 22235 18037 22244 18071
rect 22192 18028 22244 18037
rect 22652 18071 22704 18080
rect 22652 18037 22661 18071
rect 22661 18037 22695 18071
rect 22695 18037 22704 18071
rect 22652 18028 22704 18037
rect 23756 18071 23808 18080
rect 23756 18037 23765 18071
rect 23765 18037 23799 18071
rect 23799 18037 23808 18071
rect 23756 18028 23808 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1952 17824 2004 17876
rect 5356 17824 5408 17876
rect 6460 17867 6512 17876
rect 6460 17833 6469 17867
rect 6469 17833 6503 17867
rect 6503 17833 6512 17867
rect 6460 17824 6512 17833
rect 7104 17824 7156 17876
rect 7840 17824 7892 17876
rect 9956 17867 10008 17876
rect 9956 17833 9965 17867
rect 9965 17833 9999 17867
rect 9999 17833 10008 17867
rect 9956 17824 10008 17833
rect 11704 17824 11756 17876
rect 12624 17824 12676 17876
rect 14648 17824 14700 17876
rect 14924 17867 14976 17876
rect 14924 17833 14933 17867
rect 14933 17833 14967 17867
rect 14967 17833 14976 17867
rect 14924 17824 14976 17833
rect 16212 17824 16264 17876
rect 16396 17867 16448 17876
rect 16396 17833 16405 17867
rect 16405 17833 16439 17867
rect 16439 17833 16448 17867
rect 16396 17824 16448 17833
rect 19340 17824 19392 17876
rect 20720 17867 20772 17876
rect 20720 17833 20729 17867
rect 20729 17833 20763 17867
rect 20763 17833 20772 17867
rect 20720 17824 20772 17833
rect 22560 17867 22612 17876
rect 22560 17833 22569 17867
rect 22569 17833 22603 17867
rect 22603 17833 22612 17867
rect 22560 17824 22612 17833
rect 22652 17824 22704 17876
rect 2044 17756 2096 17808
rect 2688 17756 2740 17808
rect 3424 17756 3476 17808
rect 4160 17756 4212 17808
rect 8024 17799 8076 17808
rect 8024 17765 8033 17799
rect 8033 17765 8067 17799
rect 8067 17765 8076 17799
rect 8024 17756 8076 17765
rect 8852 17756 8904 17808
rect 10600 17756 10652 17808
rect 11796 17799 11848 17808
rect 11796 17765 11805 17799
rect 11805 17765 11839 17799
rect 11839 17765 11848 17799
rect 11796 17756 11848 17765
rect 12716 17799 12768 17808
rect 12716 17765 12725 17799
rect 12725 17765 12759 17799
rect 12759 17765 12768 17799
rect 12716 17756 12768 17765
rect 2320 17688 2372 17740
rect 1584 17620 1636 17672
rect 3516 17620 3568 17672
rect 4160 17663 4212 17672
rect 4160 17629 4169 17663
rect 4169 17629 4203 17663
rect 4203 17629 4212 17663
rect 4436 17663 4488 17672
rect 4160 17620 4212 17629
rect 4436 17629 4445 17663
rect 4445 17629 4479 17663
rect 4479 17629 4488 17663
rect 4436 17620 4488 17629
rect 20 17552 72 17604
rect 7748 17688 7800 17740
rect 12348 17688 12400 17740
rect 13544 17688 13596 17740
rect 14464 17756 14516 17808
rect 15476 17799 15528 17808
rect 15476 17765 15485 17799
rect 15485 17765 15519 17799
rect 15519 17765 15528 17799
rect 15476 17756 15528 17765
rect 18236 17799 18288 17808
rect 18236 17765 18245 17799
rect 18245 17765 18279 17799
rect 18279 17765 18288 17799
rect 18236 17756 18288 17765
rect 21088 17799 21140 17808
rect 17500 17731 17552 17740
rect 2964 17484 3016 17536
rect 5540 17527 5592 17536
rect 5540 17493 5549 17527
rect 5549 17493 5583 17527
rect 5583 17493 5592 17527
rect 5540 17484 5592 17493
rect 6000 17527 6052 17536
rect 6000 17493 6009 17527
rect 6009 17493 6043 17527
rect 6043 17493 6052 17527
rect 8300 17620 8352 17672
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 10692 17595 10744 17604
rect 10692 17561 10701 17595
rect 10701 17561 10735 17595
rect 10735 17561 10744 17595
rect 10692 17552 10744 17561
rect 11336 17552 11388 17604
rect 13636 17552 13688 17604
rect 17500 17697 17509 17731
rect 17509 17697 17543 17731
rect 17543 17697 17552 17731
rect 17500 17688 17552 17697
rect 17960 17731 18012 17740
rect 17960 17697 17969 17731
rect 17969 17697 18003 17731
rect 18003 17697 18012 17731
rect 21088 17765 21097 17799
rect 21097 17765 21131 17799
rect 21131 17765 21140 17799
rect 21088 17756 21140 17765
rect 17960 17688 18012 17697
rect 19524 17731 19576 17740
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 19524 17697 19533 17731
rect 19533 17697 19567 17731
rect 19567 17697 19576 17731
rect 19524 17688 19576 17697
rect 22468 17731 22520 17740
rect 22468 17697 22477 17731
rect 22477 17697 22511 17731
rect 22511 17697 22520 17731
rect 22468 17688 22520 17697
rect 22928 17731 22980 17740
rect 22928 17697 22937 17731
rect 22937 17697 22971 17731
rect 22971 17697 22980 17731
rect 22928 17688 22980 17697
rect 24032 17688 24084 17740
rect 25228 17688 25280 17740
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 20812 17620 20864 17672
rect 17408 17552 17460 17604
rect 19064 17552 19116 17604
rect 19248 17552 19300 17604
rect 23756 17620 23808 17672
rect 23848 17620 23900 17672
rect 22008 17552 22060 17604
rect 16764 17527 16816 17536
rect 6000 17484 6052 17493
rect 16764 17493 16773 17527
rect 16773 17493 16807 17527
rect 16807 17493 16816 17527
rect 16764 17484 16816 17493
rect 21916 17527 21968 17536
rect 21916 17493 21925 17527
rect 21925 17493 21959 17527
rect 21959 17493 21968 17527
rect 21916 17484 21968 17493
rect 24032 17484 24084 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2688 17280 2740 17332
rect 3792 17323 3844 17332
rect 3792 17289 3801 17323
rect 3801 17289 3835 17323
rect 3835 17289 3844 17323
rect 3792 17280 3844 17289
rect 4068 17323 4120 17332
rect 4068 17289 4077 17323
rect 4077 17289 4111 17323
rect 4111 17289 4120 17323
rect 4068 17280 4120 17289
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 10140 17280 10192 17332
rect 14740 17280 14792 17332
rect 15476 17323 15528 17332
rect 15476 17289 15485 17323
rect 15485 17289 15519 17323
rect 15519 17289 15528 17323
rect 15476 17280 15528 17289
rect 17500 17323 17552 17332
rect 17500 17289 17509 17323
rect 17509 17289 17543 17323
rect 17543 17289 17552 17323
rect 17500 17280 17552 17289
rect 17684 17280 17736 17332
rect 19064 17323 19116 17332
rect 10048 17212 10100 17264
rect 11796 17212 11848 17264
rect 14464 17255 14516 17264
rect 4160 17144 4212 17196
rect 12624 17144 12676 17196
rect 1032 17076 1084 17128
rect 2964 17076 3016 17128
rect 3332 17076 3384 17128
rect 5632 17076 5684 17128
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 9404 17119 9456 17128
rect 9404 17085 9413 17119
rect 9413 17085 9447 17119
rect 9447 17085 9456 17119
rect 9404 17076 9456 17085
rect 10600 17119 10652 17128
rect 10600 17085 10609 17119
rect 10609 17085 10643 17119
rect 10643 17085 10652 17119
rect 10600 17076 10652 17085
rect 10784 17076 10836 17128
rect 11244 17119 11296 17128
rect 11244 17085 11262 17119
rect 11262 17085 11296 17119
rect 11244 17076 11296 17085
rect 2780 16983 2832 16992
rect 2780 16949 2789 16983
rect 2789 16949 2823 16983
rect 2823 16949 2832 16983
rect 2780 16940 2832 16949
rect 6092 17008 6144 17060
rect 6460 16940 6512 16992
rect 10140 17008 10192 17060
rect 12164 17008 12216 17060
rect 13636 17008 13688 17060
rect 14464 17221 14473 17255
rect 14473 17221 14507 17255
rect 14507 17221 14516 17255
rect 14464 17212 14516 17221
rect 14280 17144 14332 17196
rect 16764 17144 16816 17196
rect 19064 17289 19073 17323
rect 19073 17289 19107 17323
rect 19107 17289 19116 17323
rect 19064 17280 19116 17289
rect 19524 17280 19576 17332
rect 22928 17280 22980 17332
rect 24032 17323 24084 17332
rect 24032 17289 24041 17323
rect 24041 17289 24075 17323
rect 24075 17289 24084 17323
rect 24032 17280 24084 17289
rect 22192 17212 22244 17264
rect 19616 17187 19668 17196
rect 19616 17153 19625 17187
rect 19625 17153 19659 17187
rect 19659 17153 19668 17187
rect 19616 17144 19668 17153
rect 20260 17144 20312 17196
rect 20444 17144 20496 17196
rect 20996 17144 21048 17196
rect 18236 17076 18288 17128
rect 22468 17119 22520 17128
rect 22468 17085 22477 17119
rect 22477 17085 22511 17119
rect 22511 17085 22520 17119
rect 22468 17076 22520 17085
rect 26240 17280 26292 17332
rect 16580 17008 16632 17060
rect 18788 17051 18840 17060
rect 18788 17017 18797 17051
rect 18797 17017 18831 17051
rect 18831 17017 18840 17051
rect 18788 17008 18840 17017
rect 8300 16940 8352 16992
rect 13820 16940 13872 16992
rect 16304 16940 16356 16992
rect 18880 16940 18932 16992
rect 21088 17008 21140 17060
rect 20720 16940 20772 16992
rect 21916 17008 21968 17060
rect 21640 16940 21692 16992
rect 24032 16940 24084 16992
rect 25228 16940 25280 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2044 16736 2096 16788
rect 5632 16736 5684 16788
rect 6000 16736 6052 16788
rect 6828 16779 6880 16788
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 10784 16736 10836 16788
rect 14280 16736 14332 16788
rect 1676 16668 1728 16720
rect 2872 16668 2924 16720
rect 3148 16711 3200 16720
rect 3148 16677 3157 16711
rect 3157 16677 3191 16711
rect 3191 16677 3200 16711
rect 3148 16668 3200 16677
rect 4068 16711 4120 16720
rect 4068 16677 4077 16711
rect 4077 16677 4111 16711
rect 4111 16677 4120 16711
rect 4068 16668 4120 16677
rect 1584 16600 1636 16652
rect 4160 16643 4212 16652
rect 4160 16609 4169 16643
rect 4169 16609 4203 16643
rect 4203 16609 4212 16643
rect 4160 16600 4212 16609
rect 4344 16600 4396 16652
rect 5908 16600 5960 16652
rect 6092 16643 6144 16652
rect 6092 16609 6101 16643
rect 6101 16609 6135 16643
rect 6135 16609 6144 16643
rect 6092 16600 6144 16609
rect 8392 16668 8444 16720
rect 9404 16711 9456 16720
rect 9404 16677 9413 16711
rect 9413 16677 9447 16711
rect 9447 16677 9456 16711
rect 9404 16668 9456 16677
rect 10140 16668 10192 16720
rect 13544 16711 13596 16720
rect 13544 16677 13553 16711
rect 13553 16677 13587 16711
rect 13587 16677 13596 16711
rect 13544 16668 13596 16677
rect 13820 16711 13872 16720
rect 13820 16677 13829 16711
rect 13829 16677 13863 16711
rect 13863 16677 13872 16711
rect 13820 16668 13872 16677
rect 15476 16668 15528 16720
rect 16120 16668 16172 16720
rect 8484 16643 8536 16652
rect 8484 16609 8493 16643
rect 8493 16609 8527 16643
rect 8527 16609 8536 16643
rect 8484 16600 8536 16609
rect 12348 16643 12400 16652
rect 2504 16575 2556 16584
rect 2504 16541 2513 16575
rect 2513 16541 2547 16575
rect 2547 16541 2556 16575
rect 2504 16532 2556 16541
rect 5448 16532 5500 16584
rect 9036 16575 9088 16584
rect 9036 16541 9045 16575
rect 9045 16541 9079 16575
rect 9079 16541 9088 16575
rect 9036 16532 9088 16541
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 17960 16736 18012 16788
rect 20260 16779 20312 16788
rect 20260 16745 20269 16779
rect 20269 16745 20303 16779
rect 20303 16745 20312 16779
rect 20260 16736 20312 16745
rect 20720 16779 20772 16788
rect 20720 16745 20729 16779
rect 20729 16745 20763 16779
rect 20763 16745 20772 16779
rect 20720 16736 20772 16745
rect 17316 16668 17368 16720
rect 19432 16711 19484 16720
rect 19432 16677 19441 16711
rect 19441 16677 19475 16711
rect 19475 16677 19484 16711
rect 19432 16668 19484 16677
rect 20444 16668 20496 16720
rect 12256 16532 12308 16584
rect 3884 16464 3936 16516
rect 12624 16464 12676 16516
rect 14188 16532 14240 16584
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 17776 16532 17828 16584
rect 19984 16532 20036 16584
rect 20904 16668 20956 16720
rect 21640 16668 21692 16720
rect 23020 16600 23072 16652
rect 23940 16643 23992 16652
rect 23940 16609 23949 16643
rect 23949 16609 23983 16643
rect 23983 16609 23992 16643
rect 23940 16600 23992 16609
rect 15384 16464 15436 16516
rect 16580 16464 16632 16516
rect 17040 16464 17092 16516
rect 21548 16464 21600 16516
rect 2320 16396 2372 16448
rect 2688 16396 2740 16448
rect 4988 16396 5040 16448
rect 6092 16396 6144 16448
rect 11336 16439 11388 16448
rect 11336 16405 11345 16439
rect 11345 16405 11379 16439
rect 11379 16405 11388 16439
rect 11336 16396 11388 16405
rect 11428 16396 11480 16448
rect 16304 16396 16356 16448
rect 18236 16396 18288 16448
rect 22376 16396 22428 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1676 16235 1728 16244
rect 1676 16201 1685 16235
rect 1685 16201 1719 16235
rect 1719 16201 1728 16235
rect 1676 16192 1728 16201
rect 1952 16192 2004 16244
rect 2504 16192 2556 16244
rect 2872 16192 2924 16244
rect 4160 16192 4212 16244
rect 5356 16192 5408 16244
rect 6000 16192 6052 16244
rect 7472 16192 7524 16244
rect 7748 16192 7800 16244
rect 8392 16192 8444 16244
rect 10876 16192 10928 16244
rect 12348 16192 12400 16244
rect 16764 16192 16816 16244
rect 18788 16192 18840 16244
rect 5172 16124 5224 16176
rect 7840 16124 7892 16176
rect 11244 16124 11296 16176
rect 8300 16056 8352 16108
rect 9680 16056 9732 16108
rect 10692 16056 10744 16108
rect 11428 16056 11480 16108
rect 15292 16124 15344 16176
rect 16120 16167 16172 16176
rect 16120 16133 16129 16167
rect 16129 16133 16163 16167
rect 16163 16133 16172 16167
rect 18880 16167 18932 16176
rect 16120 16124 16172 16133
rect 18880 16133 18889 16167
rect 18889 16133 18923 16167
rect 18923 16133 18932 16167
rect 18880 16124 18932 16133
rect 1216 15988 1268 16040
rect 2688 15988 2740 16040
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 5264 15963 5316 15972
rect 5264 15929 5273 15963
rect 5273 15929 5307 15963
rect 5307 15929 5316 15963
rect 5264 15920 5316 15929
rect 5356 15963 5408 15972
rect 5356 15929 5365 15963
rect 5365 15929 5399 15963
rect 5399 15929 5408 15963
rect 8484 15988 8536 16040
rect 11060 16031 11112 16040
rect 11060 15997 11069 16031
rect 11069 15997 11103 16031
rect 11103 15997 11112 16031
rect 11060 15988 11112 15997
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 5356 15920 5408 15929
rect 9036 15920 9088 15972
rect 9404 15963 9456 15972
rect 9404 15929 9413 15963
rect 9413 15929 9447 15963
rect 9447 15929 9456 15963
rect 9404 15920 9456 15929
rect 10048 15920 10100 15972
rect 17040 16099 17092 16108
rect 14280 16031 14332 16040
rect 14280 15997 14289 16031
rect 14289 15997 14323 16031
rect 14323 15997 14332 16031
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 17776 16099 17828 16108
rect 17776 16065 17785 16099
rect 17785 16065 17819 16099
rect 17819 16065 17828 16099
rect 17776 16056 17828 16065
rect 21916 16192 21968 16244
rect 22376 16235 22428 16244
rect 22376 16201 22385 16235
rect 22385 16201 22419 16235
rect 22419 16201 22428 16235
rect 22376 16192 22428 16201
rect 23020 16235 23072 16244
rect 23020 16201 23029 16235
rect 23029 16201 23063 16235
rect 23063 16201 23072 16235
rect 23020 16192 23072 16201
rect 23940 16235 23992 16244
rect 23940 16201 23949 16235
rect 23949 16201 23983 16235
rect 23983 16201 23992 16235
rect 23940 16192 23992 16201
rect 14280 15988 14332 15997
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 18972 16031 19024 16040
rect 18972 15997 18981 16031
rect 18981 15997 19015 16031
rect 19015 15997 19024 16031
rect 18972 15988 19024 15997
rect 19432 15988 19484 16040
rect 21640 15988 21692 16040
rect 13728 15963 13780 15972
rect 13728 15929 13737 15963
rect 13737 15929 13771 15963
rect 13771 15929 13780 15963
rect 13728 15920 13780 15929
rect 16396 15963 16448 15972
rect 16396 15929 16405 15963
rect 16405 15929 16439 15963
rect 16439 15929 16448 15963
rect 16396 15920 16448 15929
rect 2780 15852 2832 15904
rect 4988 15895 5040 15904
rect 4988 15861 4997 15895
rect 4997 15861 5031 15895
rect 5031 15861 5040 15895
rect 4988 15852 5040 15861
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 10140 15852 10192 15904
rect 10692 15852 10744 15904
rect 12624 15852 12676 15904
rect 15660 15852 15712 15904
rect 16304 15852 16356 15904
rect 18880 15920 18932 15972
rect 21180 15920 21232 15972
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 21640 15852 21692 15904
rect 23020 15852 23072 15904
rect 24032 15852 24084 15904
rect 27620 15852 27672 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 5264 15648 5316 15700
rect 7380 15648 7432 15700
rect 9680 15648 9732 15700
rect 11244 15648 11296 15700
rect 13268 15691 13320 15700
rect 13268 15657 13277 15691
rect 13277 15657 13311 15691
rect 13311 15657 13320 15691
rect 13268 15648 13320 15657
rect 13820 15691 13872 15700
rect 13820 15657 13829 15691
rect 13829 15657 13863 15691
rect 13863 15657 13872 15691
rect 14280 15691 14332 15700
rect 13820 15648 13872 15657
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 19984 15648 20036 15700
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 3332 15580 3384 15632
rect 7196 15580 7248 15632
rect 8852 15580 8904 15632
rect 10784 15580 10836 15632
rect 11428 15623 11480 15632
rect 11428 15589 11437 15623
rect 11437 15589 11471 15623
rect 11471 15589 11480 15623
rect 11428 15580 11480 15589
rect 11980 15623 12032 15632
rect 11980 15589 11989 15623
rect 11989 15589 12023 15623
rect 12023 15589 12032 15623
rect 11980 15580 12032 15589
rect 15660 15580 15712 15632
rect 21180 15623 21232 15632
rect 21180 15589 21189 15623
rect 21189 15589 21223 15623
rect 21223 15589 21232 15623
rect 21180 15580 21232 15589
rect 21916 15580 21968 15632
rect 2412 15555 2464 15564
rect 2412 15521 2421 15555
rect 2421 15521 2455 15555
rect 2455 15521 2464 15555
rect 2412 15512 2464 15521
rect 2596 15512 2648 15564
rect 3056 15512 3108 15564
rect 4068 15512 4120 15564
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 6460 15555 6512 15564
rect 6460 15521 6469 15555
rect 6469 15521 6503 15555
rect 6503 15521 6512 15555
rect 6460 15512 6512 15521
rect 8024 15555 8076 15564
rect 3792 15444 3844 15496
rect 2504 15419 2556 15428
rect 2504 15385 2513 15419
rect 2513 15385 2547 15419
rect 2547 15385 2556 15419
rect 2504 15376 2556 15385
rect 3700 15376 3752 15428
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8024 15512 8076 15521
rect 8208 15512 8260 15564
rect 8484 15555 8536 15564
rect 8484 15521 8493 15555
rect 8493 15521 8527 15555
rect 8527 15521 8536 15555
rect 8484 15512 8536 15521
rect 12532 15512 12584 15564
rect 13084 15555 13136 15564
rect 13084 15521 13093 15555
rect 13093 15521 13127 15555
rect 13127 15521 13136 15555
rect 13084 15512 13136 15521
rect 17684 15512 17736 15564
rect 18236 15555 18288 15564
rect 18236 15521 18245 15555
rect 18245 15521 18279 15555
rect 18279 15521 18288 15555
rect 18236 15512 18288 15521
rect 5080 15376 5132 15428
rect 7840 15444 7892 15496
rect 9404 15444 9456 15496
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 11336 15487 11388 15496
rect 10048 15444 10100 15453
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 15844 15444 15896 15496
rect 21824 15512 21876 15564
rect 23296 15512 23348 15564
rect 24124 15512 24176 15564
rect 18512 15487 18564 15496
rect 18512 15453 18521 15487
rect 18521 15453 18555 15487
rect 18555 15453 18564 15487
rect 18512 15444 18564 15453
rect 21548 15487 21600 15496
rect 21548 15453 21557 15487
rect 21557 15453 21591 15487
rect 21591 15453 21600 15487
rect 21548 15444 21600 15453
rect 23112 15487 23164 15496
rect 23112 15453 23121 15487
rect 23121 15453 23155 15487
rect 23155 15453 23164 15487
rect 23112 15444 23164 15453
rect 6552 15419 6604 15428
rect 6552 15385 6561 15419
rect 6561 15385 6595 15419
rect 6595 15385 6604 15419
rect 6552 15376 6604 15385
rect 12992 15376 13044 15428
rect 16212 15419 16264 15428
rect 16212 15385 16221 15419
rect 16221 15385 16255 15419
rect 16255 15385 16264 15419
rect 16212 15376 16264 15385
rect 22928 15376 22980 15428
rect 2872 15308 2924 15360
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 12256 15351 12308 15360
rect 12256 15317 12265 15351
rect 12265 15317 12299 15351
rect 12299 15317 12308 15351
rect 12256 15308 12308 15317
rect 16396 15308 16448 15360
rect 17684 15308 17736 15360
rect 18972 15351 19024 15360
rect 18972 15317 18981 15351
rect 18981 15317 19015 15351
rect 19015 15317 19024 15351
rect 18972 15308 19024 15317
rect 20444 15351 20496 15360
rect 20444 15317 20453 15351
rect 20453 15317 20487 15351
rect 20487 15317 20496 15351
rect 20444 15308 20496 15317
rect 22192 15351 22244 15360
rect 22192 15317 22201 15351
rect 22201 15317 22235 15351
rect 22235 15317 22244 15351
rect 22192 15308 22244 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2596 15104 2648 15156
rect 8484 15104 8536 15156
rect 10784 15104 10836 15156
rect 11428 15036 11480 15088
rect 2412 14968 2464 15020
rect 8392 15011 8444 15020
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 2872 14900 2924 14909
rect 3700 14900 3752 14952
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 9036 14968 9088 15020
rect 16488 15104 16540 15156
rect 16856 15104 16908 15156
rect 17592 15104 17644 15156
rect 21180 15104 21232 15156
rect 21732 15147 21784 15156
rect 21732 15113 21741 15147
rect 21741 15113 21775 15147
rect 21775 15113 21784 15147
rect 21732 15104 21784 15113
rect 16396 15036 16448 15088
rect 17316 15036 17368 15088
rect 22836 15036 22888 15088
rect 18972 14968 19024 15020
rect 20444 15011 20496 15020
rect 20444 14977 20453 15011
rect 20453 14977 20487 15011
rect 20487 14977 20496 15011
rect 20444 14968 20496 14977
rect 22192 14968 22244 15020
rect 4068 14900 4120 14952
rect 5908 14900 5960 14952
rect 6092 14943 6144 14952
rect 6092 14909 6101 14943
rect 6101 14909 6135 14943
rect 6135 14909 6144 14943
rect 6460 14943 6512 14952
rect 6092 14900 6144 14909
rect 6460 14909 6469 14943
rect 6469 14909 6503 14943
rect 6503 14909 6512 14943
rect 6460 14900 6512 14909
rect 9404 14900 9456 14952
rect 11060 14900 11112 14952
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 14648 14943 14700 14952
rect 14648 14909 14657 14943
rect 14657 14909 14691 14943
rect 14691 14909 14700 14943
rect 14648 14900 14700 14909
rect 16488 14943 16540 14952
rect 16488 14909 16497 14943
rect 16497 14909 16531 14943
rect 16531 14909 16540 14943
rect 16488 14900 16540 14909
rect 3516 14832 3568 14884
rect 5080 14875 5132 14884
rect 5080 14841 5089 14875
rect 5089 14841 5123 14875
rect 5123 14841 5132 14875
rect 5080 14832 5132 14841
rect 5356 14832 5408 14884
rect 8300 14875 8352 14884
rect 8300 14841 8309 14875
rect 8309 14841 8343 14875
rect 8343 14841 8352 14875
rect 8300 14832 8352 14841
rect 2688 14807 2740 14816
rect 2688 14773 2697 14807
rect 2697 14773 2731 14807
rect 2731 14773 2740 14807
rect 2688 14764 2740 14773
rect 5448 14764 5500 14816
rect 6000 14764 6052 14816
rect 8024 14764 8076 14816
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 10140 14764 10192 14816
rect 12992 14764 13044 14816
rect 13636 14764 13688 14816
rect 14740 14764 14792 14816
rect 17592 14832 17644 14884
rect 18236 14832 18288 14884
rect 19248 14900 19300 14952
rect 18788 14875 18840 14884
rect 18788 14841 18797 14875
rect 18797 14841 18831 14875
rect 18831 14841 18840 14875
rect 18788 14832 18840 14841
rect 20536 14875 20588 14884
rect 20536 14841 20545 14875
rect 20545 14841 20579 14875
rect 20579 14841 20588 14875
rect 20536 14832 20588 14841
rect 21272 14832 21324 14884
rect 17776 14764 17828 14816
rect 22008 14832 22060 14884
rect 22744 14832 22796 14884
rect 24124 14900 24176 14952
rect 22928 14807 22980 14816
rect 22928 14773 22937 14807
rect 22937 14773 22971 14807
rect 22971 14773 22980 14807
rect 22928 14764 22980 14773
rect 23296 14807 23348 14816
rect 23296 14773 23305 14807
rect 23305 14773 23339 14807
rect 23339 14773 23348 14807
rect 23296 14764 23348 14773
rect 27620 14764 27672 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2504 14560 2556 14612
rect 3240 14560 3292 14612
rect 5080 14492 5132 14544
rect 5540 14560 5592 14612
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 9956 14560 10008 14612
rect 11428 14560 11480 14612
rect 10784 14492 10836 14544
rect 13084 14560 13136 14612
rect 13636 14603 13688 14612
rect 13636 14569 13645 14603
rect 13645 14569 13679 14603
rect 13679 14569 13688 14603
rect 13636 14560 13688 14569
rect 13728 14560 13780 14612
rect 14372 14560 14424 14612
rect 14648 14603 14700 14612
rect 14648 14569 14657 14603
rect 14657 14569 14691 14603
rect 14691 14569 14700 14603
rect 14648 14560 14700 14569
rect 15660 14560 15712 14612
rect 18788 14603 18840 14612
rect 18788 14569 18797 14603
rect 18797 14569 18831 14603
rect 18831 14569 18840 14603
rect 18788 14560 18840 14569
rect 20536 14560 20588 14612
rect 21916 14603 21968 14612
rect 21916 14569 21925 14603
rect 21925 14569 21959 14603
rect 21959 14569 21968 14603
rect 21916 14560 21968 14569
rect 15752 14535 15804 14544
rect 15752 14501 15761 14535
rect 15761 14501 15795 14535
rect 15795 14501 15804 14535
rect 15752 14492 15804 14501
rect 18880 14492 18932 14544
rect 20260 14492 20312 14544
rect 21088 14535 21140 14544
rect 21088 14501 21097 14535
rect 21097 14501 21131 14535
rect 21131 14501 21140 14535
rect 21088 14492 21140 14501
rect 23020 14492 23072 14544
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 2504 14331 2556 14340
rect 2504 14297 2513 14331
rect 2513 14297 2547 14331
rect 2547 14297 2556 14331
rect 2504 14288 2556 14297
rect 3700 14424 3752 14476
rect 4436 14424 4488 14476
rect 5356 14467 5408 14476
rect 5356 14433 5365 14467
rect 5365 14433 5399 14467
rect 5399 14433 5408 14467
rect 5356 14424 5408 14433
rect 5540 14424 5592 14476
rect 5908 14424 5960 14476
rect 7196 14424 7248 14476
rect 7748 14424 7800 14476
rect 8484 14467 8536 14476
rect 8484 14433 8493 14467
rect 8493 14433 8527 14467
rect 8527 14433 8536 14467
rect 8484 14424 8536 14433
rect 8852 14424 8904 14476
rect 17408 14467 17460 14476
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 17592 14424 17644 14476
rect 18512 14424 18564 14476
rect 19892 14424 19944 14476
rect 3976 14356 4028 14408
rect 6000 14356 6052 14408
rect 7840 14356 7892 14408
rect 9496 14356 9548 14408
rect 11152 14356 11204 14408
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 13176 14356 13228 14408
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 16488 14356 16540 14408
rect 20444 14356 20496 14408
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 22100 14356 22152 14408
rect 22836 14399 22888 14408
rect 22836 14365 22845 14399
rect 22845 14365 22879 14399
rect 22879 14365 22888 14399
rect 22836 14356 22888 14365
rect 3516 14331 3568 14340
rect 3516 14297 3525 14331
rect 3525 14297 3559 14331
rect 3559 14297 3568 14331
rect 3516 14288 3568 14297
rect 5448 14331 5500 14340
rect 5448 14297 5457 14331
rect 5457 14297 5491 14331
rect 5491 14297 5500 14331
rect 5448 14288 5500 14297
rect 6552 14288 6604 14340
rect 20168 14288 20220 14340
rect 3608 14220 3660 14272
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4252 14220 4304 14229
rect 5356 14220 5408 14272
rect 7012 14220 7064 14272
rect 9036 14263 9088 14272
rect 9036 14229 9045 14263
rect 9045 14229 9079 14263
rect 9079 14229 9088 14263
rect 9036 14220 9088 14229
rect 14372 14220 14424 14272
rect 16304 14220 16356 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 7748 14016 7800 14068
rect 9588 14059 9640 14068
rect 9588 14025 9597 14059
rect 9597 14025 9631 14059
rect 9631 14025 9640 14059
rect 9588 14016 9640 14025
rect 11428 14059 11480 14068
rect 11428 14025 11437 14059
rect 11437 14025 11471 14059
rect 11471 14025 11480 14059
rect 11428 14016 11480 14025
rect 12348 14016 12400 14068
rect 12532 14059 12584 14068
rect 12532 14025 12541 14059
rect 12541 14025 12575 14059
rect 12575 14025 12584 14059
rect 12532 14016 12584 14025
rect 13360 14016 13412 14068
rect 13636 14016 13688 14068
rect 14372 14016 14424 14068
rect 15752 14016 15804 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 17592 14016 17644 14068
rect 21088 14016 21140 14068
rect 22744 14059 22796 14068
rect 22744 14025 22753 14059
rect 22753 14025 22787 14059
rect 22787 14025 22796 14059
rect 22744 14016 22796 14025
rect 23020 14059 23072 14068
rect 23020 14025 23029 14059
rect 23029 14025 23063 14059
rect 23063 14025 23072 14059
rect 23020 14016 23072 14025
rect 3516 13948 3568 14000
rect 2872 13880 2924 13932
rect 1676 13812 1728 13864
rect 3792 13880 3844 13932
rect 1492 13744 1544 13796
rect 2504 13744 2556 13796
rect 1124 13676 1176 13728
rect 2964 13719 3016 13728
rect 2964 13685 2973 13719
rect 2973 13685 3007 13719
rect 3007 13685 3016 13719
rect 2964 13676 3016 13685
rect 3516 13744 3568 13796
rect 3700 13855 3752 13864
rect 3700 13821 3709 13855
rect 3709 13821 3743 13855
rect 3743 13821 3752 13855
rect 3700 13812 3752 13821
rect 5172 13948 5224 14000
rect 4988 13880 5040 13932
rect 7472 13880 7524 13932
rect 8484 13880 8536 13932
rect 9036 13880 9088 13932
rect 5356 13812 5408 13864
rect 5540 13812 5592 13864
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 4436 13744 4488 13796
rect 8300 13744 8352 13796
rect 10784 13948 10836 14000
rect 15844 13948 15896 14000
rect 19892 13991 19944 14000
rect 19892 13957 19901 13991
rect 19901 13957 19935 13991
rect 19935 13957 19944 13991
rect 19892 13948 19944 13957
rect 20260 13991 20312 14000
rect 20260 13957 20269 13991
rect 20269 13957 20303 13991
rect 20303 13957 20312 13991
rect 20260 13948 20312 13957
rect 10692 13880 10744 13932
rect 11152 13923 11204 13932
rect 11152 13889 11161 13923
rect 11161 13889 11195 13923
rect 11195 13889 11204 13923
rect 11152 13880 11204 13889
rect 12532 13880 12584 13932
rect 14740 13880 14792 13932
rect 16212 13880 16264 13932
rect 16488 13923 16540 13932
rect 16488 13889 16497 13923
rect 16497 13889 16531 13923
rect 16531 13889 16540 13923
rect 16488 13880 16540 13889
rect 18788 13880 18840 13932
rect 5448 13676 5500 13728
rect 6000 13676 6052 13728
rect 7196 13676 7248 13728
rect 9956 13719 10008 13728
rect 9956 13685 9965 13719
rect 9965 13685 9999 13719
rect 9999 13685 10008 13719
rect 9956 13676 10008 13685
rect 12624 13676 12676 13728
rect 15844 13812 15896 13864
rect 14648 13787 14700 13796
rect 14648 13753 14657 13787
rect 14657 13753 14691 13787
rect 14691 13753 14700 13787
rect 14648 13744 14700 13753
rect 16212 13787 16264 13796
rect 14372 13676 14424 13728
rect 16212 13753 16221 13787
rect 16221 13753 16255 13787
rect 16255 13753 16264 13787
rect 16212 13744 16264 13753
rect 16396 13744 16448 13796
rect 18420 13676 18472 13728
rect 18880 13676 18932 13728
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 22744 13812 22796 13864
rect 23388 13812 23440 13864
rect 20536 13744 20588 13796
rect 21364 13719 21416 13728
rect 21364 13685 21373 13719
rect 21373 13685 21407 13719
rect 21407 13685 21416 13719
rect 21364 13676 21416 13685
rect 22100 13719 22152 13728
rect 22100 13685 22109 13719
rect 22109 13685 22143 13719
rect 22143 13685 22152 13719
rect 22100 13676 22152 13685
rect 22192 13676 22244 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1676 13515 1728 13524
rect 1676 13481 1685 13515
rect 1685 13481 1719 13515
rect 1719 13481 1728 13515
rect 9496 13515 9548 13524
rect 1676 13472 1728 13481
rect 2780 13404 2832 13456
rect 4252 13447 4304 13456
rect 2688 13336 2740 13388
rect 4252 13413 4261 13447
rect 4261 13413 4295 13447
rect 4295 13413 4304 13447
rect 4252 13404 4304 13413
rect 5448 13404 5500 13456
rect 9496 13481 9505 13515
rect 9505 13481 9539 13515
rect 9539 13481 9548 13515
rect 9496 13472 9548 13481
rect 13176 13515 13228 13524
rect 11796 13404 11848 13456
rect 12624 13404 12676 13456
rect 13176 13481 13185 13515
rect 13185 13481 13219 13515
rect 13219 13481 13228 13515
rect 13176 13472 13228 13481
rect 15568 13472 15620 13524
rect 13452 13404 13504 13456
rect 16028 13472 16080 13524
rect 16396 13472 16448 13524
rect 18420 13472 18472 13524
rect 20168 13515 20220 13524
rect 20168 13481 20177 13515
rect 20177 13481 20211 13515
rect 20211 13481 20220 13515
rect 20168 13472 20220 13481
rect 20444 13515 20496 13524
rect 20444 13481 20453 13515
rect 20453 13481 20487 13515
rect 20487 13481 20496 13515
rect 20444 13472 20496 13481
rect 22100 13472 22152 13524
rect 19432 13404 19484 13456
rect 20536 13404 20588 13456
rect 20720 13404 20772 13456
rect 21364 13404 21416 13456
rect 22652 13447 22704 13456
rect 22652 13413 22661 13447
rect 22661 13413 22695 13447
rect 22695 13413 22704 13447
rect 22652 13404 22704 13413
rect 3516 13268 3568 13320
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 4344 13268 4396 13320
rect 6000 13336 6052 13388
rect 7840 13379 7892 13388
rect 7840 13345 7849 13379
rect 7849 13345 7883 13379
rect 7883 13345 7892 13379
rect 7840 13336 7892 13345
rect 8484 13336 8536 13388
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 13268 13379 13320 13388
rect 13268 13345 13277 13379
rect 13277 13345 13311 13379
rect 13311 13345 13320 13379
rect 13268 13336 13320 13345
rect 13636 13379 13688 13388
rect 13636 13345 13645 13379
rect 13645 13345 13679 13379
rect 13679 13345 13688 13379
rect 13636 13336 13688 13345
rect 6092 13268 6144 13320
rect 6276 13268 6328 13320
rect 7380 13268 7432 13320
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 11888 13311 11940 13320
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 14372 13268 14424 13320
rect 15384 13336 15436 13388
rect 17040 13379 17092 13388
rect 17040 13345 17049 13379
rect 17049 13345 17083 13379
rect 17083 13345 17092 13379
rect 17040 13336 17092 13345
rect 24216 13336 24268 13388
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 17868 13268 17920 13320
rect 21456 13268 21508 13320
rect 22560 13311 22612 13320
rect 22560 13277 22569 13311
rect 22569 13277 22603 13311
rect 22603 13277 22612 13311
rect 22560 13268 22612 13277
rect 22836 13311 22888 13320
rect 22836 13277 22845 13311
rect 22845 13277 22879 13311
rect 22879 13277 22888 13311
rect 22836 13268 22888 13277
rect 3332 13132 3384 13184
rect 3792 13132 3844 13184
rect 3976 13132 4028 13184
rect 7288 13200 7340 13252
rect 14464 13200 14516 13252
rect 14648 13243 14700 13252
rect 14648 13209 14657 13243
rect 14657 13209 14691 13243
rect 14691 13209 14700 13243
rect 14648 13200 14700 13209
rect 21272 13200 21324 13252
rect 23940 13200 23992 13252
rect 5172 13175 5224 13184
rect 5172 13141 5181 13175
rect 5181 13141 5215 13175
rect 5215 13141 5224 13175
rect 5172 13132 5224 13141
rect 6736 13175 6788 13184
rect 6736 13141 6745 13175
rect 6745 13141 6779 13175
rect 6779 13141 6788 13175
rect 6736 13132 6788 13141
rect 7104 13132 7156 13184
rect 7472 13132 7524 13184
rect 10876 13132 10928 13184
rect 11244 13132 11296 13184
rect 12624 13175 12676 13184
rect 12624 13141 12633 13175
rect 12633 13141 12667 13175
rect 12667 13141 12676 13175
rect 12624 13132 12676 13141
rect 13176 13132 13228 13184
rect 17500 13132 17552 13184
rect 19064 13175 19116 13184
rect 19064 13141 19073 13175
rect 19073 13141 19107 13175
rect 19107 13141 19116 13175
rect 19064 13132 19116 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 3240 12928 3292 12980
rect 5448 12971 5500 12980
rect 5448 12937 5457 12971
rect 5457 12937 5491 12971
rect 5491 12937 5500 12971
rect 5448 12928 5500 12937
rect 7840 12971 7892 12980
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 14372 12971 14424 12980
rect 14372 12937 14381 12971
rect 14381 12937 14415 12971
rect 14415 12937 14424 12971
rect 14372 12928 14424 12937
rect 15568 12928 15620 12980
rect 16672 12928 16724 12980
rect 20720 12971 20772 12980
rect 20720 12937 20729 12971
rect 20729 12937 20763 12971
rect 20763 12937 20772 12971
rect 20720 12928 20772 12937
rect 21364 12928 21416 12980
rect 22652 12928 22704 12980
rect 24216 12928 24268 12980
rect 24952 12928 25004 12980
rect 2780 12903 2832 12912
rect 2780 12869 2789 12903
rect 2789 12869 2823 12903
rect 2823 12869 2832 12903
rect 2780 12860 2832 12869
rect 5540 12860 5592 12912
rect 6828 12860 6880 12912
rect 1400 12792 1452 12844
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 4344 12792 4396 12844
rect 6736 12792 6788 12844
rect 7380 12860 7432 12912
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 3700 12767 3752 12776
rect 3700 12733 3709 12767
rect 3709 12733 3743 12767
rect 3743 12733 3752 12767
rect 3700 12724 3752 12733
rect 4252 12767 4304 12776
rect 4252 12733 4261 12767
rect 4261 12733 4295 12767
rect 4295 12733 4304 12767
rect 4252 12724 4304 12733
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 6184 12724 6236 12776
rect 13636 12860 13688 12912
rect 16028 12903 16080 12912
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 11888 12792 11940 12844
rect 11980 12792 12032 12844
rect 14832 12792 14884 12844
rect 15660 12792 15712 12844
rect 8484 12724 8536 12776
rect 13176 12767 13228 12776
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 4712 12656 4764 12708
rect 6000 12656 6052 12708
rect 7012 12699 7064 12708
rect 7012 12665 7021 12699
rect 7021 12665 7055 12699
rect 7055 12665 7064 12699
rect 7012 12656 7064 12665
rect 10876 12699 10928 12708
rect 10876 12665 10885 12699
rect 10885 12665 10919 12699
rect 10919 12665 10928 12699
rect 10876 12656 10928 12665
rect 3516 12631 3568 12640
rect 3516 12597 3525 12631
rect 3525 12597 3559 12631
rect 3559 12597 3568 12631
rect 3516 12588 3568 12597
rect 6092 12631 6144 12640
rect 6092 12597 6101 12631
rect 6101 12597 6135 12631
rect 6135 12597 6144 12631
rect 6092 12588 6144 12597
rect 10140 12588 10192 12640
rect 11152 12656 11204 12708
rect 11888 12588 11940 12640
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 12624 12656 12676 12708
rect 14096 12724 14148 12776
rect 16028 12869 16037 12903
rect 16037 12869 16071 12903
rect 16071 12869 16080 12903
rect 16028 12860 16080 12869
rect 17408 12860 17460 12912
rect 18512 12860 18564 12912
rect 23388 12860 23440 12912
rect 19432 12835 19484 12844
rect 19432 12801 19441 12835
rect 19441 12801 19475 12835
rect 19475 12801 19484 12835
rect 19432 12792 19484 12801
rect 20168 12792 20220 12844
rect 16488 12767 16540 12776
rect 16488 12733 16532 12767
rect 16532 12733 16540 12767
rect 18236 12767 18288 12776
rect 16488 12724 16540 12733
rect 18236 12733 18245 12767
rect 18245 12733 18279 12767
rect 18279 12733 18288 12767
rect 18236 12724 18288 12733
rect 25136 12767 25188 12776
rect 25136 12733 25145 12767
rect 25145 12733 25179 12767
rect 25179 12733 25188 12767
rect 25136 12724 25188 12733
rect 14004 12699 14056 12708
rect 14004 12665 14013 12699
rect 14013 12665 14047 12699
rect 14047 12665 14056 12699
rect 14004 12656 14056 12665
rect 15016 12699 15068 12708
rect 15016 12665 15025 12699
rect 15025 12665 15059 12699
rect 15059 12665 15068 12699
rect 15016 12656 15068 12665
rect 13084 12588 13136 12640
rect 14648 12588 14700 12640
rect 17316 12656 17368 12708
rect 17776 12656 17828 12708
rect 21272 12699 21324 12708
rect 15936 12588 15988 12640
rect 17040 12631 17092 12640
rect 17040 12597 17049 12631
rect 17049 12597 17083 12631
rect 17083 12597 17092 12631
rect 17040 12588 17092 12597
rect 17868 12631 17920 12640
rect 17868 12597 17877 12631
rect 17877 12597 17911 12631
rect 17911 12597 17920 12631
rect 17868 12588 17920 12597
rect 18420 12588 18472 12640
rect 19064 12588 19116 12640
rect 21272 12665 21281 12699
rect 21281 12665 21315 12699
rect 21315 12665 21324 12699
rect 21272 12656 21324 12665
rect 21364 12699 21416 12708
rect 21364 12665 21373 12699
rect 21373 12665 21407 12699
rect 21407 12665 21416 12699
rect 21364 12656 21416 12665
rect 21548 12656 21600 12708
rect 21916 12699 21968 12708
rect 21916 12665 21925 12699
rect 21925 12665 21959 12699
rect 21959 12665 21968 12699
rect 21916 12656 21968 12665
rect 22008 12656 22060 12708
rect 23204 12656 23256 12708
rect 24216 12656 24268 12708
rect 22836 12631 22888 12640
rect 22836 12597 22845 12631
rect 22845 12597 22879 12631
rect 22879 12597 22888 12631
rect 22836 12588 22888 12597
rect 24032 12588 24084 12640
rect 24676 12588 24728 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 3332 12427 3384 12436
rect 3332 12393 3341 12427
rect 3341 12393 3375 12427
rect 3375 12393 3384 12427
rect 3332 12384 3384 12393
rect 3700 12427 3752 12436
rect 3700 12393 3709 12427
rect 3709 12393 3743 12427
rect 3743 12393 3752 12427
rect 3700 12384 3752 12393
rect 4344 12384 4396 12436
rect 4804 12384 4856 12436
rect 4988 12427 5040 12436
rect 4988 12393 4997 12427
rect 4997 12393 5031 12427
rect 5031 12393 5040 12427
rect 4988 12384 5040 12393
rect 7012 12384 7064 12436
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 8852 12384 8904 12436
rect 11152 12427 11204 12436
rect 11152 12393 11161 12427
rect 11161 12393 11195 12427
rect 11195 12393 11204 12427
rect 11152 12384 11204 12393
rect 12624 12384 12676 12436
rect 13820 12427 13872 12436
rect 13820 12393 13829 12427
rect 13829 12393 13863 12427
rect 13863 12393 13872 12427
rect 15016 12427 15068 12436
rect 13820 12384 13872 12393
rect 15016 12393 15025 12427
rect 15025 12393 15059 12427
rect 15059 12393 15068 12427
rect 15016 12384 15068 12393
rect 15292 12384 15344 12436
rect 16672 12427 16724 12436
rect 16672 12393 16681 12427
rect 16681 12393 16715 12427
rect 16715 12393 16724 12427
rect 16672 12384 16724 12393
rect 17868 12384 17920 12436
rect 21916 12384 21968 12436
rect 22560 12384 22612 12436
rect 22836 12384 22888 12436
rect 25136 12427 25188 12436
rect 25136 12393 25145 12427
rect 25145 12393 25179 12427
rect 25179 12393 25188 12427
rect 25136 12384 25188 12393
rect 4160 12316 4212 12368
rect 6828 12316 6880 12368
rect 7196 12359 7248 12368
rect 7196 12325 7205 12359
rect 7205 12325 7239 12359
rect 7239 12325 7248 12359
rect 7196 12316 7248 12325
rect 9956 12316 10008 12368
rect 11060 12316 11112 12368
rect 12164 12359 12216 12368
rect 12164 12325 12173 12359
rect 12173 12325 12207 12359
rect 12207 12325 12216 12359
rect 12164 12316 12216 12325
rect 13360 12316 13412 12368
rect 15476 12359 15528 12368
rect 15476 12325 15485 12359
rect 15485 12325 15519 12359
rect 15519 12325 15528 12359
rect 15476 12316 15528 12325
rect 17316 12359 17368 12368
rect 17316 12325 17325 12359
rect 17325 12325 17359 12359
rect 17359 12325 17368 12359
rect 17316 12316 17368 12325
rect 17500 12316 17552 12368
rect 1860 12248 1912 12300
rect 2688 12291 2740 12300
rect 2688 12257 2697 12291
rect 2697 12257 2731 12291
rect 2731 12257 2740 12291
rect 2688 12248 2740 12257
rect 3240 12248 3292 12300
rect 4620 12248 4672 12300
rect 4804 12248 4856 12300
rect 4252 12180 4304 12232
rect 5448 12248 5500 12300
rect 5356 12180 5408 12232
rect 6092 12248 6144 12300
rect 8116 12248 8168 12300
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 14372 12291 14424 12300
rect 14372 12257 14381 12291
rect 14381 12257 14415 12291
rect 14415 12257 14424 12291
rect 14372 12248 14424 12257
rect 18236 12316 18288 12368
rect 19064 12248 19116 12300
rect 19248 12291 19300 12300
rect 19248 12257 19257 12291
rect 19257 12257 19291 12291
rect 19291 12257 19300 12291
rect 19248 12248 19300 12257
rect 22284 12248 22336 12300
rect 23020 12248 23072 12300
rect 23940 12291 23992 12300
rect 23940 12257 23949 12291
rect 23949 12257 23983 12291
rect 23983 12257 23992 12291
rect 23940 12248 23992 12257
rect 25504 12248 25556 12300
rect 7840 12180 7892 12232
rect 10968 12180 11020 12232
rect 14004 12180 14056 12232
rect 14464 12180 14516 12232
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 15660 12223 15712 12232
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 16948 12180 17000 12232
rect 18788 12180 18840 12232
rect 20904 12223 20956 12232
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 112 12112 164 12164
rect 4068 12112 4120 12164
rect 6828 12112 6880 12164
rect 9220 12112 9272 12164
rect 11612 12112 11664 12164
rect 18604 12112 18656 12164
rect 21272 12112 21324 12164
rect 3332 12044 3384 12096
rect 3792 12044 3844 12096
rect 4436 12044 4488 12096
rect 7104 12044 7156 12096
rect 10232 12044 10284 12096
rect 13176 12044 13228 12096
rect 13544 12044 13596 12096
rect 13728 12044 13780 12096
rect 14372 12044 14424 12096
rect 16396 12087 16448 12096
rect 16396 12053 16405 12087
rect 16405 12053 16439 12087
rect 16439 12053 16448 12087
rect 16396 12044 16448 12053
rect 20352 12044 20404 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1308 11840 1360 11892
rect 1860 11840 1912 11892
rect 2596 11840 2648 11892
rect 4068 11883 4120 11892
rect 4068 11849 4077 11883
rect 4077 11849 4111 11883
rect 4111 11849 4120 11883
rect 4068 11840 4120 11849
rect 4804 11840 4856 11892
rect 7104 11840 7156 11892
rect 9496 11840 9548 11892
rect 11888 11840 11940 11892
rect 3148 11772 3200 11824
rect 4252 11772 4304 11824
rect 6368 11772 6420 11824
rect 12256 11772 12308 11824
rect 2504 11704 2556 11756
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 7196 11704 7248 11756
rect 7840 11704 7892 11756
rect 8852 11704 8904 11756
rect 2596 11679 2648 11688
rect 2596 11645 2605 11679
rect 2605 11645 2639 11679
rect 2639 11645 2648 11679
rect 2596 11636 2648 11645
rect 3884 11679 3936 11688
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 2412 11568 2464 11620
rect 5540 11568 5592 11620
rect 7012 11679 7064 11688
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 8116 11636 8168 11688
rect 9496 11679 9548 11688
rect 3424 11543 3476 11552
rect 3424 11509 3433 11543
rect 3433 11509 3467 11543
rect 3467 11509 3476 11543
rect 3424 11500 3476 11509
rect 5264 11500 5316 11552
rect 6644 11500 6696 11552
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 12072 11704 12124 11756
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 9680 11568 9732 11620
rect 11980 11636 12032 11688
rect 12808 11636 12860 11688
rect 14004 11840 14056 11892
rect 15476 11840 15528 11892
rect 19064 11883 19116 11892
rect 19064 11849 19073 11883
rect 19073 11849 19107 11883
rect 19107 11849 19116 11883
rect 19064 11840 19116 11849
rect 19248 11840 19300 11892
rect 23940 11883 23992 11892
rect 23940 11849 23949 11883
rect 23949 11849 23983 11883
rect 23983 11849 23992 11883
rect 23940 11840 23992 11849
rect 13820 11772 13872 11824
rect 14832 11772 14884 11824
rect 16948 11815 17000 11824
rect 16948 11781 16957 11815
rect 16957 11781 16991 11815
rect 16991 11781 17000 11815
rect 16948 11772 17000 11781
rect 17316 11772 17368 11824
rect 24768 11815 24820 11824
rect 15292 11704 15344 11756
rect 18788 11747 18840 11756
rect 18788 11713 18797 11747
rect 18797 11713 18831 11747
rect 18831 11713 18840 11747
rect 18788 11704 18840 11713
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 14096 11679 14148 11688
rect 13820 11636 13872 11645
rect 14096 11645 14105 11679
rect 14105 11645 14139 11679
rect 14139 11645 14148 11679
rect 14096 11636 14148 11645
rect 20352 11679 20404 11688
rect 20352 11645 20361 11679
rect 20361 11645 20395 11679
rect 20395 11645 20404 11679
rect 20352 11636 20404 11645
rect 24768 11781 24777 11815
rect 24777 11781 24811 11815
rect 24811 11781 24820 11815
rect 24768 11772 24820 11781
rect 25504 11747 25556 11756
rect 25504 11713 25513 11747
rect 25513 11713 25547 11747
rect 25547 11713 25556 11747
rect 25504 11704 25556 11713
rect 24124 11636 24176 11688
rect 10968 11611 11020 11620
rect 10968 11577 10977 11611
rect 10977 11577 11011 11611
rect 11011 11577 11020 11611
rect 10968 11568 11020 11577
rect 14372 11611 14424 11620
rect 8852 11500 8904 11552
rect 9496 11500 9548 11552
rect 10692 11500 10744 11552
rect 11704 11500 11756 11552
rect 14372 11577 14381 11611
rect 14381 11577 14415 11611
rect 14415 11577 14424 11611
rect 14372 11568 14424 11577
rect 16396 11611 16448 11620
rect 16396 11577 16405 11611
rect 16405 11577 16439 11611
rect 16439 11577 16448 11611
rect 16396 11568 16448 11577
rect 17776 11568 17828 11620
rect 18144 11611 18196 11620
rect 18144 11577 18153 11611
rect 18153 11577 18187 11611
rect 18187 11577 18196 11611
rect 18144 11568 18196 11577
rect 20168 11543 20220 11552
rect 20168 11509 20177 11543
rect 20177 11509 20211 11543
rect 20211 11509 20220 11543
rect 20168 11500 20220 11509
rect 22284 11543 22336 11552
rect 22284 11509 22293 11543
rect 22293 11509 22327 11543
rect 22327 11509 22336 11543
rect 22284 11500 22336 11509
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 23572 11500 23624 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1400 11296 1452 11348
rect 2688 11296 2740 11348
rect 3516 11339 3568 11348
rect 3516 11305 3525 11339
rect 3525 11305 3559 11339
rect 3559 11305 3568 11339
rect 3516 11296 3568 11305
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 4620 11296 4672 11348
rect 4896 11296 4948 11348
rect 6644 11296 6696 11348
rect 7012 11296 7064 11348
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 7840 11296 7892 11305
rect 10876 11296 10928 11348
rect 12164 11339 12216 11348
rect 12164 11305 12173 11339
rect 12173 11305 12207 11339
rect 12207 11305 12216 11339
rect 12164 11296 12216 11305
rect 12532 11339 12584 11348
rect 12532 11305 12541 11339
rect 12541 11305 12575 11339
rect 12575 11305 12584 11339
rect 12532 11296 12584 11305
rect 15384 11296 15436 11348
rect 16212 11296 16264 11348
rect 9220 11228 9272 11280
rect 9312 11228 9364 11280
rect 10232 11228 10284 11280
rect 10968 11228 11020 11280
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 2688 11203 2740 11212
rect 2504 11160 2556 11169
rect 2688 11169 2697 11203
rect 2697 11169 2731 11203
rect 2731 11169 2740 11203
rect 2688 11160 2740 11169
rect 4252 11203 4304 11212
rect 4252 11169 4261 11203
rect 4261 11169 4295 11203
rect 4295 11169 4304 11203
rect 4252 11160 4304 11169
rect 6368 11160 6420 11212
rect 8024 11160 8076 11212
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 10416 11160 10468 11212
rect 11336 11160 11388 11212
rect 14832 11228 14884 11280
rect 18420 11228 18472 11280
rect 20352 11228 20404 11280
rect 21456 11228 21508 11280
rect 12992 11160 13044 11212
rect 13360 11160 13412 11212
rect 13636 11160 13688 11212
rect 14096 11203 14148 11212
rect 14096 11169 14105 11203
rect 14105 11169 14139 11203
rect 14139 11169 14148 11203
rect 14096 11160 14148 11169
rect 14372 11160 14424 11212
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 17316 11160 17368 11212
rect 17500 11203 17552 11212
rect 17500 11169 17518 11203
rect 17518 11169 17552 11203
rect 17500 11160 17552 11169
rect 18512 11160 18564 11212
rect 22836 11160 22888 11212
rect 9128 11092 9180 11144
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 19156 11092 19208 11144
rect 21272 11092 21324 11144
rect 10876 11024 10928 11076
rect 11704 11024 11756 11076
rect 20444 11024 20496 11076
rect 21088 11024 21140 11076
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 6644 10956 6696 11008
rect 7104 10999 7156 11008
rect 7104 10965 7113 10999
rect 7113 10965 7147 10999
rect 7147 10965 7156 10999
rect 7104 10956 7156 10965
rect 9312 10999 9364 11008
rect 9312 10965 9321 10999
rect 9321 10965 9355 10999
rect 9355 10965 9364 10999
rect 9312 10956 9364 10965
rect 11060 10956 11112 11008
rect 11796 10999 11848 11008
rect 11796 10965 11805 10999
rect 11805 10965 11839 10999
rect 11839 10965 11848 10999
rect 11796 10956 11848 10965
rect 16948 10956 17000 11008
rect 18052 10999 18104 11008
rect 18052 10965 18061 10999
rect 18061 10965 18095 10999
rect 18095 10965 18104 10999
rect 18052 10956 18104 10965
rect 18144 10956 18196 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2228 10795 2280 10804
rect 2228 10761 2237 10795
rect 2237 10761 2271 10795
rect 2271 10761 2280 10795
rect 2228 10752 2280 10761
rect 2596 10752 2648 10804
rect 3424 10795 3476 10804
rect 3424 10761 3433 10795
rect 3433 10761 3467 10795
rect 3467 10761 3476 10795
rect 3424 10752 3476 10761
rect 4988 10752 5040 10804
rect 6368 10752 6420 10804
rect 9588 10752 9640 10804
rect 10232 10795 10284 10804
rect 10232 10761 10241 10795
rect 10241 10761 10275 10795
rect 10275 10761 10284 10795
rect 10232 10752 10284 10761
rect 2412 10684 2464 10736
rect 8576 10684 8628 10736
rect 10416 10684 10468 10736
rect 2596 10616 2648 10668
rect 3148 10659 3200 10668
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 2688 10548 2740 10557
rect 4252 10548 4304 10600
rect 4528 10548 4580 10600
rect 5172 10616 5224 10668
rect 6276 10616 6328 10668
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 7472 10616 7524 10668
rect 10048 10616 10100 10668
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 2320 10480 2372 10532
rect 4436 10523 4488 10532
rect 4436 10489 4445 10523
rect 4445 10489 4479 10523
rect 4479 10489 4488 10523
rect 4436 10480 4488 10489
rect 7472 10480 7524 10532
rect 9312 10523 9364 10532
rect 9312 10489 9321 10523
rect 9321 10489 9355 10523
rect 9355 10489 9364 10523
rect 9312 10480 9364 10489
rect 9588 10480 9640 10532
rect 14188 10752 14240 10804
rect 14832 10795 14884 10804
rect 14832 10761 14841 10795
rect 14841 10761 14875 10795
rect 14875 10761 14884 10795
rect 14832 10752 14884 10761
rect 16396 10752 16448 10804
rect 11796 10684 11848 10736
rect 20168 10752 20220 10804
rect 21456 10795 21508 10804
rect 21088 10727 21140 10736
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 18052 10616 18104 10668
rect 21088 10693 21097 10727
rect 21097 10693 21131 10727
rect 21131 10693 21140 10727
rect 21088 10684 21140 10693
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 22836 10795 22888 10804
rect 22836 10761 22845 10795
rect 22845 10761 22879 10795
rect 22879 10761 22888 10795
rect 22836 10752 22888 10761
rect 20536 10659 20588 10668
rect 20536 10625 20545 10659
rect 20545 10625 20579 10659
rect 20579 10625 20588 10659
rect 20536 10616 20588 10625
rect 20904 10616 20956 10668
rect 12532 10548 12584 10600
rect 12992 10548 13044 10600
rect 13636 10591 13688 10600
rect 13636 10557 13645 10591
rect 13645 10557 13679 10591
rect 13679 10557 13688 10591
rect 13636 10548 13688 10557
rect 15016 10591 15068 10600
rect 8024 10412 8076 10464
rect 10692 10412 10744 10464
rect 15016 10557 15025 10591
rect 15025 10557 15059 10591
rect 15059 10557 15068 10591
rect 15016 10548 15068 10557
rect 16396 10548 16448 10600
rect 17500 10591 17552 10600
rect 17500 10557 17509 10591
rect 17509 10557 17543 10591
rect 17543 10557 17552 10591
rect 17500 10548 17552 10557
rect 17960 10548 18012 10600
rect 22468 10591 22520 10600
rect 22468 10557 22477 10591
rect 22477 10557 22511 10591
rect 22511 10557 22520 10591
rect 22468 10548 22520 10557
rect 14832 10480 14884 10532
rect 15568 10480 15620 10532
rect 18420 10523 18472 10532
rect 18420 10489 18429 10523
rect 18429 10489 18463 10523
rect 18463 10489 18472 10523
rect 18420 10480 18472 10489
rect 14096 10412 14148 10464
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 20168 10412 20220 10464
rect 21272 10480 21324 10532
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2504 10208 2556 10260
rect 2320 10140 2372 10192
rect 3424 10208 3476 10260
rect 3608 10208 3660 10260
rect 4528 10251 4580 10260
rect 4528 10217 4537 10251
rect 4537 10217 4571 10251
rect 4571 10217 4580 10251
rect 4528 10208 4580 10217
rect 6828 10208 6880 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9312 10208 9364 10260
rect 12164 10208 12216 10260
rect 4068 10140 4120 10192
rect 4436 10140 4488 10192
rect 5448 10140 5500 10192
rect 1308 10072 1360 10124
rect 6276 10115 6328 10124
rect 6276 10081 6285 10115
rect 6285 10081 6319 10115
rect 6319 10081 6328 10115
rect 6276 10072 6328 10081
rect 6644 10140 6696 10192
rect 8024 10183 8076 10192
rect 8024 10149 8033 10183
rect 8033 10149 8067 10183
rect 8067 10149 8076 10183
rect 8024 10140 8076 10149
rect 9588 10140 9640 10192
rect 11152 10140 11204 10192
rect 6460 10072 6512 10124
rect 10876 10115 10928 10124
rect 10876 10081 10885 10115
rect 10885 10081 10919 10115
rect 10919 10081 10928 10115
rect 10876 10072 10928 10081
rect 11888 10072 11940 10124
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 7196 9936 7248 9988
rect 9220 9936 9272 9988
rect 10324 10004 10376 10056
rect 12532 10208 12584 10260
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 16028 10251 16080 10260
rect 16028 10217 16037 10251
rect 16037 10217 16071 10251
rect 16071 10217 16080 10251
rect 16028 10208 16080 10217
rect 18420 10208 18472 10260
rect 19156 10251 19208 10260
rect 19156 10217 19165 10251
rect 19165 10217 19199 10251
rect 19199 10217 19208 10251
rect 19156 10208 19208 10217
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 15016 10183 15068 10192
rect 15016 10149 15025 10183
rect 15025 10149 15059 10183
rect 15059 10149 15068 10183
rect 15016 10140 15068 10149
rect 16396 10183 16448 10192
rect 16396 10149 16405 10183
rect 16405 10149 16439 10183
rect 16439 10149 16448 10183
rect 16396 10140 16448 10149
rect 16948 10183 17000 10192
rect 16948 10149 16957 10183
rect 16957 10149 16991 10183
rect 16991 10149 17000 10183
rect 16948 10140 17000 10149
rect 17776 10183 17828 10192
rect 17776 10149 17785 10183
rect 17785 10149 17819 10183
rect 17819 10149 17828 10183
rect 17776 10140 17828 10149
rect 21088 10183 21140 10192
rect 12808 10072 12860 10124
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 13636 10072 13688 10081
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 14096 10115 14148 10124
rect 13820 10072 13872 10081
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 14096 10072 14148 10081
rect 17500 10072 17552 10124
rect 19432 10072 19484 10124
rect 21088 10149 21097 10183
rect 21097 10149 21131 10183
rect 21131 10149 21140 10183
rect 21088 10140 21140 10149
rect 24032 10208 24084 10260
rect 24768 10251 24820 10260
rect 24768 10217 24777 10251
rect 24777 10217 24811 10251
rect 24811 10217 24820 10251
rect 24768 10208 24820 10217
rect 25228 10140 25280 10192
rect 23388 10072 23440 10124
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 16304 10004 16356 10013
rect 20996 10047 21048 10056
rect 20996 10013 21005 10047
rect 21005 10013 21039 10047
rect 21039 10013 21048 10047
rect 20996 10004 21048 10013
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 21272 10004 21324 10013
rect 23296 10004 23348 10056
rect 25136 10072 25188 10124
rect 11428 9936 11480 9988
rect 2412 9911 2464 9920
rect 2412 9877 2421 9911
rect 2421 9877 2455 9911
rect 2455 9877 2464 9911
rect 2412 9868 2464 9877
rect 7380 9911 7432 9920
rect 7380 9877 7389 9911
rect 7389 9877 7423 9911
rect 7423 9877 7432 9911
rect 7380 9868 7432 9877
rect 9496 9868 9548 9920
rect 11336 9911 11388 9920
rect 11336 9877 11345 9911
rect 11345 9877 11379 9911
rect 11379 9877 11388 9911
rect 11336 9868 11388 9877
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 19984 9868 20036 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1860 9707 1912 9716
rect 1860 9673 1869 9707
rect 1869 9673 1903 9707
rect 1903 9673 1912 9707
rect 1860 9664 1912 9673
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 1860 9460 1912 9512
rect 2872 9392 2924 9444
rect 3516 9664 3568 9716
rect 5356 9664 5408 9716
rect 6460 9664 6512 9716
rect 12808 9664 12860 9716
rect 13636 9707 13688 9716
rect 13636 9673 13645 9707
rect 13645 9673 13679 9707
rect 13679 9673 13688 9707
rect 13636 9664 13688 9673
rect 16396 9664 16448 9716
rect 17500 9707 17552 9716
rect 17500 9673 17509 9707
rect 17509 9673 17543 9707
rect 17543 9673 17552 9707
rect 17500 9664 17552 9673
rect 18972 9664 19024 9716
rect 23388 9664 23440 9716
rect 24676 9664 24728 9716
rect 25136 9707 25188 9716
rect 25136 9673 25145 9707
rect 25145 9673 25179 9707
rect 25179 9673 25188 9707
rect 25136 9664 25188 9673
rect 3792 9596 3844 9648
rect 4252 9528 4304 9580
rect 4896 9528 4948 9580
rect 6276 9596 6328 9648
rect 7564 9596 7616 9648
rect 4068 9460 4120 9512
rect 4528 9460 4580 9512
rect 4712 9503 4764 9512
rect 4712 9469 4721 9503
rect 4721 9469 4755 9503
rect 4755 9469 4764 9503
rect 4712 9460 4764 9469
rect 7380 9528 7432 9580
rect 7196 9460 7248 9512
rect 7564 9503 7616 9512
rect 7564 9469 7573 9503
rect 7573 9469 7607 9503
rect 7607 9469 7616 9503
rect 7564 9460 7616 9469
rect 14188 9596 14240 9648
rect 16304 9596 16356 9648
rect 18144 9596 18196 9648
rect 21272 9596 21324 9648
rect 12716 9528 12768 9580
rect 14096 9528 14148 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 16028 9528 16080 9580
rect 19984 9571 20036 9580
rect 19984 9537 19993 9571
rect 19993 9537 20027 9571
rect 20027 9537 20036 9571
rect 19984 9528 20036 9537
rect 21088 9528 21140 9580
rect 21824 9528 21876 9580
rect 23296 9528 23348 9580
rect 9220 9503 9272 9512
rect 6644 9392 6696 9444
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 9956 9460 10008 9512
rect 10324 9503 10376 9512
rect 10324 9469 10333 9503
rect 10333 9469 10367 9503
rect 10367 9469 10376 9503
rect 10324 9460 10376 9469
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 11520 9460 11572 9512
rect 11888 9503 11940 9512
rect 11888 9469 11897 9503
rect 11897 9469 11931 9503
rect 11931 9469 11940 9503
rect 11888 9460 11940 9469
rect 13728 9460 13780 9512
rect 3516 9324 3568 9376
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 7564 9324 7616 9376
rect 10140 9324 10192 9376
rect 12348 9392 12400 9444
rect 10784 9324 10836 9376
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12440 9324 12492 9333
rect 17316 9392 17368 9444
rect 16120 9324 16172 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 18972 9392 19024 9444
rect 19524 9392 19576 9444
rect 19984 9392 20036 9444
rect 17776 9324 17828 9333
rect 19432 9324 19484 9376
rect 24400 9367 24452 9376
rect 24400 9333 24409 9367
rect 24409 9333 24443 9367
rect 24443 9333 24452 9367
rect 24400 9324 24452 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 3792 9163 3844 9172
rect 3792 9129 3801 9163
rect 3801 9129 3835 9163
rect 3835 9129 3844 9163
rect 3792 9120 3844 9129
rect 4160 9163 4212 9172
rect 4160 9129 4169 9163
rect 4169 9129 4203 9163
rect 4203 9129 4212 9163
rect 4160 9120 4212 9129
rect 6644 9120 6696 9172
rect 7932 9120 7984 9172
rect 9312 9120 9364 9172
rect 12348 9163 12400 9172
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 12808 9163 12860 9172
rect 12808 9129 12817 9163
rect 12817 9129 12851 9163
rect 12851 9129 12860 9163
rect 12808 9120 12860 9129
rect 15568 9120 15620 9172
rect 17776 9120 17828 9172
rect 19984 9163 20036 9172
rect 19984 9129 19993 9163
rect 19993 9129 20027 9163
rect 20027 9129 20036 9163
rect 19984 9120 20036 9129
rect 24400 9120 24452 9172
rect 3976 9052 4028 9104
rect 1584 8984 1636 9036
rect 4252 9027 4304 9036
rect 4252 8993 4261 9027
rect 4261 8993 4295 9027
rect 4295 8993 4304 9027
rect 4252 8984 4304 8993
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 4712 8984 4764 9036
rect 3792 8916 3844 8968
rect 5356 8984 5408 9036
rect 6736 9052 6788 9104
rect 7472 9052 7524 9104
rect 8024 9095 8076 9104
rect 8024 9061 8033 9095
rect 8033 9061 8067 9095
rect 8067 9061 8076 9095
rect 8024 9052 8076 9061
rect 11888 9052 11940 9104
rect 6920 8984 6972 9036
rect 8668 9027 8720 9036
rect 8668 8993 8686 9027
rect 8686 8993 8720 9027
rect 8668 8984 8720 8993
rect 9956 9027 10008 9036
rect 9956 8993 9965 9027
rect 9965 8993 9999 9027
rect 9999 8993 10008 9027
rect 9956 8984 10008 8993
rect 10140 9027 10192 9036
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10140 8984 10192 8993
rect 10692 9027 10744 9036
rect 10692 8993 10701 9027
rect 10701 8993 10735 9027
rect 10735 8993 10744 9027
rect 10692 8984 10744 8993
rect 10968 9027 11020 9036
rect 10968 8993 10977 9027
rect 10977 8993 11011 9027
rect 11011 8993 11020 9027
rect 10968 8984 11020 8993
rect 17224 9095 17276 9104
rect 17224 9061 17233 9095
rect 17233 9061 17267 9095
rect 17267 9061 17276 9095
rect 17224 9052 17276 9061
rect 18420 9052 18472 9104
rect 19064 9052 19116 9104
rect 12992 8984 13044 9036
rect 13728 9027 13780 9036
rect 13728 8993 13737 9027
rect 13737 8993 13771 9027
rect 13771 8993 13780 9027
rect 13728 8984 13780 8993
rect 14188 9027 14240 9036
rect 14188 8993 14197 9027
rect 14197 8993 14231 9027
rect 14231 8993 14240 9027
rect 14188 8984 14240 8993
rect 23756 8984 23808 9036
rect 24676 8984 24728 9036
rect 7196 8916 7248 8968
rect 14832 8916 14884 8968
rect 17132 8959 17184 8968
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 17316 8916 17368 8968
rect 18972 8959 19024 8968
rect 18972 8925 18981 8959
rect 18981 8925 19015 8959
rect 19015 8925 19024 8959
rect 18972 8916 19024 8925
rect 1308 8848 1360 8900
rect 20996 8848 21048 8900
rect 1768 8780 1820 8832
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 11428 8823 11480 8832
rect 11428 8789 11437 8823
rect 11437 8789 11471 8823
rect 11471 8789 11480 8823
rect 11428 8780 11480 8789
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 18880 8780 18932 8832
rect 22284 8780 22336 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 1860 8576 1912 8628
rect 4252 8576 4304 8628
rect 4620 8576 4672 8628
rect 8668 8619 8720 8628
rect 8668 8585 8677 8619
rect 8677 8585 8711 8619
rect 8711 8585 8720 8619
rect 8668 8576 8720 8585
rect 10140 8576 10192 8628
rect 10692 8576 10744 8628
rect 12992 8576 13044 8628
rect 13084 8576 13136 8628
rect 15568 8576 15620 8628
rect 16120 8619 16172 8628
rect 16120 8585 16129 8619
rect 16129 8585 16163 8619
rect 16163 8585 16172 8619
rect 16120 8576 16172 8585
rect 24676 8619 24728 8628
rect 24676 8585 24685 8619
rect 24685 8585 24719 8619
rect 24719 8585 24728 8619
rect 24676 8576 24728 8585
rect 1768 8508 1820 8560
rect 2320 8440 2372 8492
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3516 8440 3568 8492
rect 8208 8508 8260 8560
rect 9496 8508 9548 8560
rect 10968 8508 11020 8560
rect 12716 8551 12768 8560
rect 12716 8517 12725 8551
rect 12725 8517 12759 8551
rect 12759 8517 12768 8551
rect 12716 8508 12768 8517
rect 12808 8508 12860 8560
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 12348 8440 12400 8492
rect 15476 8440 15528 8492
rect 18052 8508 18104 8560
rect 21824 8508 21876 8560
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 1860 8304 1912 8356
rect 3792 8236 3844 8288
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 7104 8304 7156 8356
rect 9588 8347 9640 8356
rect 9588 8313 9597 8347
rect 9597 8313 9631 8347
rect 9631 8313 9640 8347
rect 9588 8304 9640 8313
rect 12808 8372 12860 8424
rect 12992 8372 13044 8424
rect 13544 8372 13596 8424
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 13728 8372 13780 8381
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 15200 8415 15252 8424
rect 15200 8381 15209 8415
rect 15209 8381 15243 8415
rect 15243 8381 15252 8415
rect 15200 8372 15252 8381
rect 15936 8372 15988 8424
rect 16948 8415 17000 8424
rect 16948 8381 16957 8415
rect 16957 8381 16991 8415
rect 16991 8381 17000 8415
rect 16948 8372 17000 8381
rect 17224 8372 17276 8424
rect 17132 8304 17184 8356
rect 17500 8304 17552 8356
rect 6736 8236 6788 8288
rect 10048 8236 10100 8288
rect 10968 8236 11020 8288
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 15568 8279 15620 8288
rect 15568 8245 15577 8279
rect 15577 8245 15611 8279
rect 15611 8245 15620 8279
rect 15568 8236 15620 8245
rect 16580 8236 16632 8288
rect 17592 8236 17644 8288
rect 19064 8279 19116 8288
rect 19064 8245 19073 8279
rect 19073 8245 19107 8279
rect 19107 8245 19116 8279
rect 19064 8236 19116 8245
rect 23756 8236 23808 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1676 8032 1728 8084
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 3516 8075 3568 8084
rect 3516 8041 3525 8075
rect 3525 8041 3559 8075
rect 3559 8041 3568 8075
rect 3516 8032 3568 8041
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 4620 8032 4672 8041
rect 6920 8032 6972 8084
rect 7472 8032 7524 8084
rect 9588 8032 9640 8084
rect 9956 8032 10008 8084
rect 10968 8032 11020 8084
rect 11152 8075 11204 8084
rect 11152 8041 11161 8075
rect 11161 8041 11195 8075
rect 11195 8041 11204 8075
rect 11152 8032 11204 8041
rect 11520 8032 11572 8084
rect 13544 8075 13596 8084
rect 13544 8041 13553 8075
rect 13553 8041 13587 8075
rect 13587 8041 13596 8075
rect 13544 8032 13596 8041
rect 14832 8032 14884 8084
rect 15200 8032 15252 8084
rect 17500 8075 17552 8084
rect 17500 8041 17509 8075
rect 17509 8041 17543 8075
rect 17543 8041 17552 8075
rect 17500 8032 17552 8041
rect 2872 7964 2924 8016
rect 2228 7896 2280 7948
rect 2412 7939 2464 7948
rect 2412 7905 2421 7939
rect 2421 7905 2455 7939
rect 2455 7905 2464 7939
rect 2412 7896 2464 7905
rect 4160 7896 4212 7948
rect 7748 7964 7800 8016
rect 12440 7964 12492 8016
rect 12716 8007 12768 8016
rect 12716 7973 12725 8007
rect 12725 7973 12759 8007
rect 12759 7973 12768 8007
rect 15476 8007 15528 8016
rect 12716 7964 12768 7973
rect 15476 7973 15485 8007
rect 15485 7973 15519 8007
rect 15519 7973 15528 8007
rect 15476 7964 15528 7973
rect 16120 7964 16172 8016
rect 18420 7964 18472 8016
rect 19064 7964 19116 8016
rect 9588 7896 9640 7948
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 8208 7828 8260 7880
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 12348 7896 12400 7948
rect 17776 7896 17828 7948
rect 18236 7896 18288 7948
rect 23204 7896 23256 7948
rect 24676 7896 24728 7948
rect 16396 7828 16448 7880
rect 17316 7828 17368 7880
rect 8484 7803 8536 7812
rect 8484 7769 8493 7803
rect 8493 7769 8527 7803
rect 8527 7769 8536 7803
rect 8484 7760 8536 7769
rect 12164 7760 12216 7812
rect 13452 7760 13504 7812
rect 2228 7692 2280 7744
rect 4804 7692 4856 7744
rect 5264 7692 5316 7744
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 27620 7692 27672 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2228 7488 2280 7540
rect 7012 7488 7064 7540
rect 8208 7488 8260 7540
rect 10048 7531 10100 7540
rect 10048 7497 10057 7531
rect 10057 7497 10091 7531
rect 10091 7497 10100 7531
rect 10048 7488 10100 7497
rect 11152 7531 11204 7540
rect 11152 7497 11161 7531
rect 11161 7497 11195 7531
rect 11195 7497 11204 7531
rect 11152 7488 11204 7497
rect 13084 7488 13136 7540
rect 16120 7488 16172 7540
rect 18236 7531 18288 7540
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 24676 7531 24728 7540
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 2412 7420 2464 7472
rect 7748 7420 7800 7472
rect 5264 7352 5316 7404
rect 5448 7395 5500 7404
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 5448 7352 5500 7361
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 9588 7395 9640 7404
rect 8484 7352 8536 7361
rect 9588 7361 9597 7395
rect 9597 7361 9631 7395
rect 9631 7361 9640 7395
rect 9588 7352 9640 7361
rect 10968 7352 11020 7404
rect 12716 7352 12768 7404
rect 16580 7395 16632 7404
rect 16580 7361 16589 7395
rect 16589 7361 16623 7395
rect 16623 7361 16632 7395
rect 16580 7352 16632 7361
rect 4804 7284 4856 7336
rect 11704 7284 11756 7336
rect 16120 7327 16172 7336
rect 16120 7293 16129 7327
rect 16129 7293 16163 7327
rect 16163 7293 16172 7327
rect 16120 7284 16172 7293
rect 4252 7259 4304 7268
rect 4252 7225 4261 7259
rect 4261 7225 4295 7259
rect 4295 7225 4304 7259
rect 4252 7216 4304 7225
rect 8116 7259 8168 7268
rect 2320 7148 2372 7200
rect 4620 7148 4672 7200
rect 4896 7191 4948 7200
rect 4896 7157 4905 7191
rect 4905 7157 4939 7191
rect 4939 7157 4948 7191
rect 8116 7225 8125 7259
rect 8125 7225 8159 7259
rect 8159 7225 8168 7259
rect 8116 7216 8168 7225
rect 8208 7259 8260 7268
rect 8208 7225 8217 7259
rect 8217 7225 8251 7259
rect 8251 7225 8260 7259
rect 8208 7216 8260 7225
rect 10048 7216 10100 7268
rect 10876 7259 10928 7268
rect 10876 7225 10885 7259
rect 10885 7225 10919 7259
rect 10919 7225 10928 7259
rect 10876 7216 10928 7225
rect 17316 7191 17368 7200
rect 4896 7148 4948 7157
rect 17316 7157 17325 7191
rect 17325 7157 17359 7191
rect 17359 7157 17368 7191
rect 17316 7148 17368 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 4160 6944 4212 6996
rect 8116 6987 8168 6996
rect 8116 6953 8125 6987
rect 8125 6953 8159 6987
rect 8159 6953 8168 6987
rect 8116 6944 8168 6953
rect 8300 6944 8352 6996
rect 10784 6987 10836 6996
rect 10784 6953 10793 6987
rect 10793 6953 10827 6987
rect 10827 6953 10836 6987
rect 10784 6944 10836 6953
rect 12440 6944 12492 6996
rect 4804 6876 4856 6928
rect 6736 6919 6788 6928
rect 6736 6885 6745 6919
rect 6745 6885 6779 6919
rect 6779 6885 6788 6919
rect 6736 6876 6788 6885
rect 9956 6919 10008 6928
rect 9956 6885 9965 6919
rect 9965 6885 9999 6919
rect 9999 6885 10008 6919
rect 9956 6876 10008 6885
rect 11704 6876 11756 6928
rect 12164 6919 12216 6928
rect 12164 6885 12173 6919
rect 12173 6885 12207 6919
rect 12207 6885 12216 6919
rect 12164 6876 12216 6885
rect 24768 6808 24820 6860
rect 4528 6740 4580 6792
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 7012 6740 7064 6792
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 10876 6740 10928 6792
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 5264 6672 5316 6724
rect 2964 6604 3016 6656
rect 4160 6604 4212 6656
rect 27620 6604 27672 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 4252 6400 4304 6452
rect 6736 6400 6788 6452
rect 11520 6400 11572 6452
rect 24768 6400 24820 6452
rect 5172 6332 5224 6384
rect 21364 6332 21416 6384
rect 4896 6264 4948 6316
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 9956 6264 10008 6316
rect 11704 6264 11756 6316
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 16396 6196 16448 6248
rect 5080 6171 5132 6180
rect 5080 6137 5089 6171
rect 5089 6137 5123 6171
rect 5123 6137 5132 6171
rect 5080 6128 5132 6137
rect 5172 6171 5224 6180
rect 5172 6137 5181 6171
rect 5181 6137 5215 6171
rect 5215 6137 5224 6171
rect 5172 6128 5224 6137
rect 2964 6103 3016 6112
rect 2964 6069 2973 6103
rect 2973 6069 3007 6103
rect 3007 6069 3016 6103
rect 2964 6060 3016 6069
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 5540 6060 5592 6112
rect 7012 6103 7064 6112
rect 7012 6069 7021 6103
rect 7021 6069 7055 6103
rect 7055 6069 7064 6103
rect 7012 6060 7064 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 7012 5856 7064 5908
rect 24584 5856 24636 5908
rect 5172 5788 5224 5840
rect 5448 5831 5500 5840
rect 5448 5797 5457 5831
rect 5457 5797 5491 5831
rect 5491 5797 5500 5831
rect 5448 5788 5500 5797
rect 25228 5720 25280 5772
rect 5356 5695 5408 5704
rect 5356 5661 5365 5695
rect 5365 5661 5399 5695
rect 5399 5661 5408 5695
rect 5356 5652 5408 5661
rect 5264 5584 5316 5636
rect 4896 5516 4948 5568
rect 5448 5516 5500 5568
rect 8944 5516 8996 5568
rect 9864 5559 9916 5568
rect 9864 5525 9873 5559
rect 9873 5525 9907 5559
rect 9907 5525 9916 5559
rect 9864 5516 9916 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 4252 5312 4304 5364
rect 4988 5312 5040 5364
rect 5448 5312 5500 5364
rect 24768 5355 24820 5364
rect 24768 5321 24777 5355
rect 24777 5321 24811 5355
rect 24811 5321 24820 5355
rect 24768 5312 24820 5321
rect 4160 5176 4212 5228
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 5080 5176 5132 5228
rect 19432 5108 19484 5160
rect 4988 5083 5040 5092
rect 4988 5049 4997 5083
rect 4997 5049 5031 5083
rect 5031 5049 5040 5083
rect 4988 5040 5040 5049
rect 25228 5015 25280 5024
rect 25228 4981 25237 5015
rect 25237 4981 25271 5015
rect 25271 4981 25280 5015
rect 25228 4972 25280 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 4896 4811 4948 4820
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 5356 4811 5408 4820
rect 5356 4777 5365 4811
rect 5365 4777 5399 4811
rect 5399 4777 5408 4811
rect 5356 4768 5408 4777
rect 1216 4632 1268 4684
rect 1676 4632 1728 4684
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 27620 4156 27672 4208
rect 1676 4063 1728 4072
rect 1676 4029 1685 4063
rect 1685 4029 1719 4063
rect 1719 4029 1728 4063
rect 1676 4020 1728 4029
rect 23848 4063 23900 4072
rect 23848 4029 23857 4063
rect 23857 4029 23891 4063
rect 23891 4029 23900 4063
rect 23848 4020 23900 4029
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 11428 3136 11480 3188
rect 24860 3136 24912 3188
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 25136 2839 25188 2848
rect 25136 2805 25145 2839
rect 25145 2805 25179 2839
rect 25179 2805 25188 2839
rect 25136 2796 25188 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 4528 2592 4580 2644
rect 8944 2592 8996 2644
rect 9128 2456 9180 2508
rect 16396 2592 16448 2644
rect 17868 2524 17920 2576
rect 11336 2456 11388 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 17684 2456 17736 2508
rect 25412 2524 25464 2576
rect 11888 2320 11940 2372
rect 17132 2320 17184 2372
rect 6000 2252 6052 2304
rect 9128 2295 9180 2304
rect 9128 2261 9137 2295
rect 9137 2261 9171 2295
rect 9171 2261 9180 2295
rect 9128 2252 9180 2261
rect 12992 2252 13044 2304
rect 26884 2252 26936 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 17224 144 17276 196
rect 664 76 716 128
rect 1308 76 1360 128
rect 4252 76 4304 128
rect 4804 76 4856 128
rect 9680 76 9732 128
rect 10416 76 10468 128
rect 14648 76 14700 128
rect 17960 76 18012 128
rect 18788 76 18840 128
rect 19524 76 19576 128
rect 20168 76 20220 128
rect 23572 76 23624 128
rect 24400 76 24452 128
<< metal2 >>
rect 754 27554 810 28000
rect 2318 27554 2374 28000
rect 754 27526 1164 27554
rect 754 27520 810 27526
rect 1030 22944 1086 22953
rect 1030 22879 1086 22888
rect 112 19168 164 19174
rect 112 19110 164 19116
rect 20 17604 72 17610
rect 20 17546 72 17552
rect 32 15881 60 17546
rect 18 15872 74 15881
rect 18 15807 74 15816
rect 124 14657 152 19110
rect 1044 17134 1072 22879
rect 1136 19334 1164 27526
rect 1964 27526 2374 27554
rect 1964 27418 1992 27526
rect 2318 27520 2374 27526
rect 3240 27532 3292 27538
rect 3974 27532 4030 28000
rect 5630 27554 5686 28000
rect 7286 27554 7342 28000
rect 3974 27520 3976 27532
rect 3240 27474 3292 27480
rect 4028 27520 4030 27532
rect 5552 27526 5686 27554
rect 3976 27474 4028 27480
rect 1780 27390 1992 27418
rect 1490 26888 1546 26897
rect 1490 26823 1546 26832
rect 1504 22098 1532 26823
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1504 21690 1532 22034
rect 1582 21720 1638 21729
rect 1492 21684 1544 21690
rect 1582 21655 1638 21664
rect 1492 21626 1544 21632
rect 1596 20602 1624 21655
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1582 20360 1638 20369
rect 1582 20295 1638 20304
rect 1596 20058 1624 20295
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1136 19306 1348 19334
rect 1032 17128 1084 17134
rect 1032 17070 1084 17076
rect 1216 16040 1268 16046
rect 1216 15982 1268 15988
rect 110 14648 166 14657
rect 110 14583 166 14592
rect 1124 13728 1176 13734
rect 1124 13670 1176 13676
rect 1136 13569 1164 13670
rect 1122 13560 1178 13569
rect 1122 13495 1178 13504
rect 112 12164 164 12170
rect 112 12106 164 12112
rect 124 12073 152 12106
rect 110 12064 166 12073
rect 110 11999 166 12008
rect 1228 4690 1256 15982
rect 1320 11898 1348 19306
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1688 19145 1716 19246
rect 1674 19136 1730 19145
rect 1674 19071 1730 19080
rect 1688 18970 1716 19071
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1780 18630 1808 27390
rect 1858 24440 1914 24449
rect 1858 24375 1914 24384
rect 1872 22778 1900 24375
rect 1860 22772 1912 22778
rect 1860 22714 1912 22720
rect 1872 22574 1900 22714
rect 1860 22568 1912 22574
rect 1860 22510 1912 22516
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 1952 19916 2004 19922
rect 1952 19858 2004 19864
rect 1858 19272 1914 19281
rect 1858 19207 1914 19216
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 16658 1624 17614
rect 1676 16720 1728 16726
rect 1676 16662 1728 16668
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1688 16250 1716 16662
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 12850 1440 14350
rect 1676 13864 1728 13870
rect 1872 13814 1900 19207
rect 1964 19174 1992 19858
rect 2056 19514 2084 20198
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 1964 17882 1992 19110
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 2056 17814 2084 18022
rect 2044 17808 2096 17814
rect 2044 17750 2096 17756
rect 2056 16794 2084 17750
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1964 15706 1992 16186
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1676 13806 1728 13812
rect 1492 13796 1544 13802
rect 1492 13738 1544 13744
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1308 11892 1360 11898
rect 1308 11834 1360 11840
rect 1412 11354 1440 12786
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1308 10124 1360 10130
rect 1308 10066 1360 10072
rect 1320 8906 1348 10066
rect 1308 8900 1360 8906
rect 1308 8842 1360 8848
rect 1216 4684 1268 4690
rect 1216 4626 1268 4632
rect 662 128 718 480
rect 1320 134 1348 8842
rect 1504 1193 1532 13738
rect 1688 13530 1716 13806
rect 1780 13786 1900 13814
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1582 10160 1638 10169
rect 1582 10095 1638 10104
rect 1596 9042 1624 10095
rect 1780 9364 1808 13786
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1872 12306 1900 12650
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1872 9722 1900 11834
rect 2240 10810 2268 18566
rect 2700 17814 2728 18566
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2688 17808 2740 17814
rect 2688 17750 2740 17756
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2332 16454 2360 17682
rect 2700 17338 2728 17750
rect 2792 17649 2820 18362
rect 2976 18086 3004 18770
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2778 17640 2834 17649
rect 2778 17575 2834 17584
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2976 17134 3004 17478
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 13814 2360 16390
rect 2516 16250 2544 16526
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2700 16046 2728 16390
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2424 15026 2452 15506
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2516 14618 2544 15370
rect 2608 15162 2636 15506
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2700 14822 2728 15982
rect 2792 15910 2820 16934
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2884 16250 2912 16662
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2884 14958 2912 15302
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2332 13786 2452 13814
rect 2516 13802 2544 14282
rect 2884 13938 2912 14894
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2424 12850 2452 13786
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 2976 13734 3004 17070
rect 3068 15570 3096 19110
rect 3148 18352 3200 18358
rect 3148 18294 3200 18300
rect 3160 18154 3188 18294
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 3160 16726 3188 18090
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3252 14618 3280 27474
rect 3988 27443 4016 27474
rect 5262 25528 5318 25537
rect 5262 25463 5318 25472
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4160 21412 4212 21418
rect 4160 21354 4212 21360
rect 4172 20466 4200 21354
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 3884 20324 3936 20330
rect 3884 20266 3936 20272
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3620 19310 3648 19654
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 3436 18290 3464 19246
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3436 17814 3464 18226
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 3528 17678 3556 18226
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3344 15638 3372 17070
rect 3332 15632 3384 15638
rect 3332 15574 3384 15580
rect 3516 14884 3568 14890
rect 3516 14826 3568 14832
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2700 12306 2728 13330
rect 2792 12918 2820 13398
rect 3252 12986 3280 14554
rect 3528 14346 3556 14826
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3528 14006 3556 14282
rect 3620 14278 3648 19246
rect 3712 18630 3740 19246
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3712 15434 3740 18566
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3804 17338 3832 18090
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3896 16640 3924 20266
rect 4068 19780 4120 19786
rect 4068 19722 4120 19728
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3988 18426 4016 19314
rect 4080 19310 4108 19722
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4344 19236 4396 19242
rect 4344 19178 4396 19184
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 4160 17808 4212 17814
rect 4080 17756 4160 17762
rect 4080 17750 4212 17756
rect 4080 17734 4200 17750
rect 4080 17338 4108 17734
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4080 16726 4108 17274
rect 4172 17202 4200 17614
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 4356 16658 4384 19178
rect 4436 18352 4488 18358
rect 4436 18294 4488 18300
rect 4448 17678 4476 18294
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4160 16652 4212 16658
rect 3896 16612 4016 16640
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3700 15428 3752 15434
rect 3700 15370 3752 15376
rect 3698 15056 3754 15065
rect 3804 15042 3832 15438
rect 3754 15014 3832 15042
rect 3698 14991 3754 15000
rect 3712 14958 3740 14991
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14482 3740 14894
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3528 13802 3556 13942
rect 3712 13870 3740 14418
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3700 13864 3752 13870
rect 3620 13824 3700 13852
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 3252 12782 3280 12922
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3252 12306 3280 12718
rect 3344 12442 3372 13126
rect 3528 12646 3556 13262
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2424 11218 2452 11562
rect 2516 11218 2544 11698
rect 2608 11694 2636 11834
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2700 11354 2728 12242
rect 3344 12102 3372 12378
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1872 9518 1900 9658
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1688 9336 1808 9364
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1596 8634 1624 8978
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1688 8090 1716 9336
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8566 1808 8774
rect 1872 8634 1900 9454
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 1872 8362 1900 8570
rect 2240 8430 2268 10746
rect 2424 10742 2452 11154
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 2332 10418 2360 10474
rect 2332 10390 2452 10418
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2332 9178 2360 10134
rect 2424 9926 2452 10390
rect 2516 10266 2544 11154
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2608 10674 2636 10746
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2700 10606 2728 11154
rect 3160 10674 3188 11766
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3436 10810 3464 11494
rect 3528 11354 3556 12582
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 3436 10266 3464 10746
rect 3620 10418 3648 13824
rect 3700 13806 3752 13812
rect 3804 13190 3832 13874
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3712 12442 3740 12718
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3528 10390 3648 10418
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 9722 2452 9862
rect 3528 9722 3556 10390
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2332 8498 2360 9114
rect 2884 8498 2912 9386
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 8498 3556 9318
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 2240 8090 2268 8366
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2884 8022 2912 8434
rect 3528 8090 3556 8434
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2240 7750 2268 7890
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2240 7546 2268 7686
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2424 7478 2452 7890
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1596 4826 1624 5063
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 4078 1716 4626
rect 1676 4072 1728 4078
rect 1674 4040 1676 4049
rect 1728 4040 1730 4049
rect 1674 3975 1730 3984
rect 1688 3949 1716 3975
rect 1490 1184 1546 1193
rect 1490 1119 1546 1128
rect 662 76 664 128
rect 716 76 718 128
rect 662 0 718 76
rect 1308 128 1360 134
rect 1308 70 1360 76
rect 2042 82 2098 480
rect 2332 82 2360 7142
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 6225 3004 6598
rect 2962 6216 3018 6225
rect 2962 6151 3018 6160
rect 2976 6118 3004 6151
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2976 5001 3004 6054
rect 2962 4992 3018 5001
rect 2962 4927 3018 4936
rect 3620 4154 3648 10202
rect 3804 9654 3832 12038
rect 3896 11694 3924 16458
rect 3988 14414 4016 16612
rect 4160 16594 4212 16600
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4172 16250 4200 16594
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4080 14958 4108 15506
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4264 13462 4292 14214
rect 4448 13802 4476 14418
rect 4632 13814 4660 24006
rect 5276 23662 5304 25463
rect 5552 24274 5580 27526
rect 5630 27520 5686 27526
rect 7116 27526 7342 27554
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 5552 23866 5580 24210
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5736 23322 5764 23462
rect 5724 23316 5776 23322
rect 5724 23258 5776 23264
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6932 22642 6960 23258
rect 7012 22704 7064 22710
rect 7012 22646 7064 22652
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 7024 22506 7052 22646
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 6460 22160 6512 22166
rect 6460 22102 6512 22108
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5552 21894 5580 21966
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5552 21690 5580 21830
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 6472 21350 6500 22102
rect 7024 21690 7052 22442
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 7116 21536 7144 27526
rect 7286 27520 7342 27526
rect 8942 27520 8998 28000
rect 10598 27520 10654 28000
rect 10704 27526 11008 27554
rect 10704 27520 10732 27526
rect 8956 23474 8984 27520
rect 10612 27492 10732 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 8956 23446 9076 23474
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 8576 22500 8628 22506
rect 8576 22442 8628 22448
rect 7576 22166 7604 22442
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 8024 22160 8076 22166
rect 8024 22102 8076 22108
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7024 21508 7144 21536
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 7024 21146 7052 21508
rect 7104 21412 7156 21418
rect 7104 21354 7156 21360
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 6368 21072 6420 21078
rect 6368 21014 6420 21020
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 5552 20398 5580 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6196 20466 6224 20742
rect 6184 20460 6236 20466
rect 6184 20402 6236 20408
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 5000 19514 5028 19858
rect 5552 19718 5580 20334
rect 6380 20262 6408 21014
rect 6656 20330 6684 21014
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 4908 18086 4936 18770
rect 5000 18154 5028 18770
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 5000 16454 5028 18090
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 5000 15910 5028 16390
rect 5184 16182 5212 19246
rect 5276 18834 5304 19246
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5368 18154 5396 18770
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5368 17882 5396 18090
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5368 16250 5396 17818
rect 5460 16590 5488 19654
rect 5552 19310 5580 19654
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6012 19378 6040 19790
rect 6276 19440 6328 19446
rect 6276 19382 6328 19388
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5552 17542 5580 18226
rect 6288 18086 6316 19382
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5172 16176 5224 16182
rect 5172 16118 5224 16124
rect 5368 15978 5396 16186
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5000 13938 5028 15846
rect 5276 15706 5304 15914
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5080 15428 5132 15434
rect 5080 15370 5132 15376
rect 5092 14890 5120 15370
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5092 14550 5120 14826
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 5368 14482 5396 14826
rect 5460 14822 5488 15506
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5460 14346 5488 14758
rect 5552 14618 5580 17478
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5644 16794 5672 17070
rect 6012 16794 6040 17478
rect 6092 17060 6144 17066
rect 6092 17002 6144 17008
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 6104 16658 6132 17002
rect 5908 16652 5960 16658
rect 6092 16652 6144 16658
rect 5960 16612 6040 16640
rect 5908 16594 5960 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16250 6040 16612
rect 6092 16594 6144 16600
rect 6104 16454 6132 16594
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5920 14482 5948 14894
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4436 13796 4488 13802
rect 4436 13738 4488 13744
rect 4540 13786 4660 13814
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3896 11354 3924 11630
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3804 9178 3832 9590
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3988 9110 4016 13126
rect 4172 12374 4200 13262
rect 4356 12850 4384 13262
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4448 12782 4476 13738
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4264 12238 4292 12718
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 4080 11898 4108 12106
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4264 11830 4292 12174
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4264 10606 4292 11154
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4356 10520 4384 12378
rect 4448 12102 4476 12718
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4540 10713 4568 13786
rect 5184 13190 5212 13942
rect 5368 13870 5396 14214
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4632 11354 4660 12242
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4526 10704 4582 10713
rect 4526 10639 4582 10648
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4436 10532 4488 10538
rect 4356 10492 4436 10520
rect 4436 10474 4488 10480
rect 4448 10198 4476 10474
rect 4540 10266 4568 10542
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4080 9518 4108 10134
rect 4724 9674 4752 12650
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 4816 12306 4844 12378
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4816 11898 4844 12242
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 5000 11762 5028 12378
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4356 9646 4752 9674
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3804 8294 3832 8910
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3528 4126 3648 4154
rect 3528 2417 3556 4126
rect 3514 2408 3570 2417
rect 3514 2343 3570 2352
rect 2042 54 2360 82
rect 3422 82 3478 480
rect 3804 82 3832 8230
rect 4172 7954 4200 9114
rect 4264 9042 4292 9522
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4264 8634 4292 8978
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4172 7002 4200 7890
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4172 5234 4200 6598
rect 4264 6458 4292 7210
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4264 5370 4292 6394
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4356 4154 4384 9646
rect 4908 9586 4936 11290
rect 5000 10810 5028 11698
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5184 10674 5212 13126
rect 5368 12322 5396 13806
rect 5460 13734 5488 14282
rect 5552 13870 5580 14418
rect 5920 14260 5948 14418
rect 6012 14414 6040 14758
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5920 14232 6040 14260
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 6012 13734 6040 14232
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5460 13462 5488 13670
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5460 12986 5488 13398
rect 6012 13394 6040 13670
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5368 12306 5488 12322
rect 5368 12300 5500 12306
rect 5368 12294 5448 12300
rect 5448 12242 5500 12248
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5264 11552 5316 11558
rect 5368 11540 5396 12174
rect 5316 11512 5396 11540
rect 5264 11494 5316 11500
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5368 9722 5396 11512
rect 5460 10198 5488 12242
rect 5552 11626 5580 12854
rect 6012 12714 6040 13330
rect 6104 13326 6132 14894
rect 6288 13326 6316 18022
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6104 12646 6132 13262
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6104 12306 6132 12582
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6196 11801 6224 12718
rect 6380 11830 6408 20198
rect 7116 19786 7144 21354
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7288 20800 7340 20806
rect 7288 20742 7340 20748
rect 7300 20602 7328 20742
rect 7288 20596 7340 20602
rect 7288 20538 7340 20544
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 7300 19922 7328 20266
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 7208 19310 7236 19790
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7300 19174 7328 19858
rect 7392 19378 7420 20946
rect 7760 20534 7788 21626
rect 7840 21412 7892 21418
rect 7840 21354 7892 21360
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 6472 18902 6500 19110
rect 7392 18970 7420 19314
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 6460 18896 6512 18902
rect 6460 18838 6512 18844
rect 6472 18086 6500 18838
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6472 17882 6500 18022
rect 7116 17882 7144 18090
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 6472 16998 6500 17818
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6840 16794 6868 17070
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15638 7236 15846
rect 7392 15706 7420 18566
rect 7484 16250 7512 20198
rect 7668 20058 7696 20334
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7760 19990 7788 20470
rect 7748 19984 7800 19990
rect 7748 19926 7800 19932
rect 7760 19242 7788 19926
rect 7852 19378 7880 21354
rect 7944 20806 7972 21966
rect 8036 21622 8064 22102
rect 8588 22012 8616 22442
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 8680 22166 8708 22374
rect 8956 22234 8984 22374
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 8668 22160 8720 22166
rect 8668 22102 8720 22108
rect 8668 22024 8720 22030
rect 8588 21984 8668 22012
rect 8668 21966 8720 21972
rect 8024 21616 8076 21622
rect 8024 21558 8076 21564
rect 7932 20800 7984 20806
rect 7932 20742 7984 20748
rect 7944 20369 7972 20742
rect 7930 20360 7986 20369
rect 7930 20295 7986 20304
rect 7932 19916 7984 19922
rect 7932 19858 7984 19864
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7852 18290 7880 19314
rect 7944 19174 7972 19858
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7760 17746 7788 18022
rect 7852 17882 7880 18226
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6472 14958 6500 15506
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6564 14346 6592 15370
rect 7760 14482 7788 16186
rect 7840 16176 7892 16182
rect 7840 16118 7892 16124
rect 7852 16046 7880 16118
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7852 15502 7880 15982
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 13870 7052 14214
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7208 13734 7236 14418
rect 7760 14074 7788 14418
rect 7840 14408 7892 14414
rect 7944 14396 7972 19110
rect 8036 18834 8064 21558
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8496 20058 8524 20946
rect 8680 20330 8708 21966
rect 8956 21554 8984 22170
rect 9048 21690 9076 23446
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9784 22098 9812 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9036 21684 9088 21690
rect 9036 21626 9088 21632
rect 9784 21622 9812 22034
rect 10980 21962 11008 27526
rect 11244 27532 11296 27538
rect 12254 27532 12310 28000
rect 12254 27520 12256 27532
rect 11244 27474 11296 27480
rect 12308 27520 12310 27532
rect 13910 27520 13966 28000
rect 15474 27520 15530 28000
rect 17130 27520 17186 28000
rect 18786 27520 18842 28000
rect 20442 27520 20498 28000
rect 22098 27520 22154 28000
rect 23754 27520 23810 28000
rect 25410 27520 25466 28000
rect 26240 27532 26292 27538
rect 12256 27474 12308 27480
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9772 21616 9824 21622
rect 9772 21558 9824 21564
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 9220 21412 9272 21418
rect 9220 21354 9272 21360
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8772 20330 8800 20538
rect 8852 20460 8904 20466
rect 8852 20402 8904 20408
rect 8668 20324 8720 20330
rect 8668 20266 8720 20272
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8680 20058 8708 20266
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8392 19780 8444 19786
rect 8392 19722 8444 19728
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 8128 18086 8156 18770
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 8036 17338 8064 17750
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8036 14822 8064 15506
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 7892 14368 7972 14396
rect 7840 14350 7892 14356
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7208 13138 7236 13670
rect 7300 13258 7328 13806
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 6748 12850 6776 13126
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6840 12374 6868 12854
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7024 12442 7052 12650
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6840 12170 6868 12310
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6368 11824 6420 11830
rect 6182 11792 6238 11801
rect 6368 11766 6420 11772
rect 6182 11727 6238 11736
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5552 11014 5580 11562
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4528 9512 4580 9518
rect 4712 9512 4764 9518
rect 4580 9472 4660 9500
rect 4528 9454 4580 9460
rect 4632 9042 4660 9472
rect 4712 9454 4764 9460
rect 4724 9042 4752 9454
rect 5368 9042 5396 9658
rect 6196 9217 6224 11727
rect 6380 11218 6408 11766
rect 7024 11694 7052 12378
rect 7116 12102 7144 13126
rect 7208 13110 7328 13138
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11898 7144 12038
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7208 11762 7236 12310
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6656 11354 6684 11494
rect 7024 11354 7052 11630
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6380 10810 6408 11154
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6656 10674 6684 10950
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6288 10130 6316 10610
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 10266 6868 10542
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6288 9654 6316 10066
rect 6472 9722 6500 10066
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6656 9450 6684 10134
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6182 9208 6238 9217
rect 6656 9178 6684 9386
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6182 9143 6238 9152
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 4632 8634 4660 8978
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 6748 8294 6776 9046
rect 6932 9042 6960 9318
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 4632 8090 4660 8230
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4632 7206 4660 8026
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 7342 4844 7686
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4816 6934 4844 7278
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6118 4568 6734
rect 4710 6352 4766 6361
rect 4710 6287 4766 6296
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4264 4126 4384 4154
rect 4264 134 4292 4126
rect 4540 2650 4568 6054
rect 4724 5681 4752 6287
rect 4816 6100 4844 6870
rect 4908 6322 4936 7142
rect 5184 6390 5212 8230
rect 6932 8090 6960 8978
rect 7116 8362 7144 10950
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7208 9518 7236 9930
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7208 8974 7236 9454
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7300 7993 7328 13110
rect 7392 12918 7420 13262
rect 7484 13190 7512 13874
rect 7852 13433 7880 14350
rect 7838 13424 7894 13433
rect 7838 13359 7840 13368
rect 7892 13359 7894 13368
rect 7840 13330 7892 13336
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7852 12986 7880 13330
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 8128 12306 8156 18022
rect 8220 16561 8248 19450
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8312 17678 8340 19314
rect 8404 19174 8432 19722
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8864 18154 8892 20402
rect 9232 19378 9260 21354
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 8956 18970 8984 19178
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 8956 18426 8984 18906
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 9968 18290 9996 21830
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 10060 21146 10088 21422
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 11072 21010 11100 22374
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 10704 20466 10732 20946
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10704 20262 10732 20402
rect 11072 20398 11100 20946
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 10784 20324 10836 20330
rect 10784 20266 10836 20272
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10796 19922 10824 20266
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10336 19514 10364 19858
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10138 19136 10194 19145
rect 10138 19071 10194 19080
rect 10152 18426 10180 19071
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 8864 17814 8892 18090
rect 8942 17912 8998 17921
rect 8942 17847 8998 17856
rect 8852 17808 8904 17814
rect 8852 17750 8904 17756
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8312 16998 8340 17614
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8206 16552 8262 16561
rect 8206 16487 8262 16496
rect 8220 15570 8248 16487
rect 8312 16114 8340 16934
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8404 16250 8432 16662
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8496 16046 8524 16594
rect 8956 16289 8984 17847
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9416 16726 9444 17070
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 8942 16280 8998 16289
rect 8942 16215 8998 16224
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 9048 15978 9076 16526
rect 9036 15972 9088 15978
rect 9404 15972 9456 15978
rect 9036 15914 9088 15920
rect 9324 15932 9404 15960
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8496 15162 8524 15506
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 8312 13802 8340 14826
rect 8300 13796 8352 13802
rect 8300 13738 8352 13744
rect 8404 13326 8432 14962
rect 8496 14482 8524 15098
rect 8864 14482 8892 15574
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9048 15026 9076 15302
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9324 14822 9352 15932
rect 9404 15914 9456 15920
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 14958 9444 15438
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8496 13938 8524 14418
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 8496 13394 8524 13874
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8496 12782 8524 13330
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8496 12442 8524 12718
rect 8864 12442 8892 14418
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13938 9076 14214
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9048 12850 9076 13874
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7852 11762 7880 12174
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11354 7880 11698
rect 8128 11694 8156 12242
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8864 11558 8892 11698
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 9232 11286 9260 12106
rect 9324 11286 9352 14758
rect 9416 14618 9444 14894
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9508 13530 9536 14350
rect 9600 14074 9628 18090
rect 9968 17882 9996 18226
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10152 17338 10180 17614
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10048 17264 10100 17270
rect 10048 17206 10100 17212
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16114 9720 16526
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9692 15706 9720 16050
rect 10060 15978 10088 17206
rect 10612 17134 10640 17750
rect 10704 17610 10732 18158
rect 10796 18154 10824 18770
rect 10784 18148 10836 18154
rect 10836 18108 10916 18136
rect 10784 18090 10836 18096
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 10152 16726 10180 17002
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10152 15910 10180 16662
rect 10704 16114 10732 17546
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10796 16794 10824 17070
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9508 11694 9536 11834
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7484 10538 7512 10610
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9586 7420 9862
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7484 9110 7512 10474
rect 8036 10470 8064 11154
rect 8588 10742 8616 11154
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 10198 8064 10406
rect 8024 10192 8076 10198
rect 8024 10134 8076 10140
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7576 9518 7604 9590
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7576 9382 7604 9454
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7944 9178 7972 9998
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 8036 9110 8064 10134
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7484 8090 7512 9046
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7760 8022 7788 8774
rect 8220 8566 8248 9998
rect 8208 8560 8260 8566
rect 8588 8537 8616 10678
rect 9140 10266 9168 11086
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10538 9352 10950
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9324 10266 9352 10474
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9232 9518 9260 9930
rect 9508 9926 9536 11494
rect 9600 10810 9628 14010
rect 9968 13734 9996 14554
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9968 12374 9996 13670
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9600 10538 9628 10746
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9600 10198 9628 10474
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8680 8634 8708 8978
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8208 8502 8260 8508
rect 8574 8528 8630 8537
rect 7748 8016 7800 8022
rect 7286 7984 7342 7993
rect 7748 7958 7800 7964
rect 7286 7919 7342 7928
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5276 7410 5304 7686
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 7024 7546 7052 7822
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5276 6730 5304 7346
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 5184 6186 5212 6326
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 4896 6112 4948 6118
rect 4816 6072 4896 6100
rect 4896 6054 4948 6060
rect 4710 5672 4766 5681
rect 4710 5607 4766 5616
rect 4908 5574 4936 6054
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4908 4826 4936 5170
rect 5000 5098 5028 5306
rect 5092 5234 5120 6122
rect 5184 5846 5212 6122
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 5276 5642 5304 6666
rect 5460 6322 5488 7346
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5552 6118 5580 6734
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6748 6458 6776 6870
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 7024 6118 7052 6734
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7024 5914 7052 6054
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 5448 5840 5500 5846
rect 5354 5808 5410 5817
rect 5448 5782 5500 5788
rect 5354 5743 5410 5752
rect 5368 5710 5396 5743
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 5368 4826 5396 5646
rect 5460 5574 5488 5782
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 5370 5488 5510
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 3422 54 3832 82
rect 4252 128 4304 134
rect 4252 70 4304 76
rect 4802 128 4858 480
rect 4802 76 4804 128
rect 4856 76 4858 128
rect 2042 0 2098 54
rect 3422 0 3478 54
rect 4802 0 4858 76
rect 6012 82 6040 2246
rect 6182 82 6238 480
rect 6012 54 6238 82
rect 7300 82 7328 7919
rect 7760 7478 7788 7958
rect 8220 7886 8248 8502
rect 9324 8498 9352 9114
rect 9508 8566 9536 9862
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 8574 8463 8630 8472
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9600 8090 9628 8298
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 8208 7880 8260 7886
rect 8260 7840 8340 7868
rect 8208 7822 8260 7828
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 8220 7274 8248 7482
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 8128 7002 8156 7210
rect 8312 7002 8340 7840
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8496 7410 8524 7754
rect 9600 7410 9628 7890
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 2650 8984 5510
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9140 2310 9168 2450
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 7654 82 7710 480
rect 7300 54 7710 82
rect 6182 0 6238 54
rect 7654 0 7710 54
rect 9034 82 9090 480
rect 9140 82 9168 2246
rect 9692 134 9720 11562
rect 10060 11150 10088 15438
rect 10152 14822 10180 15846
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 13938 10732 15846
rect 10796 15638 10824 16730
rect 10888 16250 10916 18108
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 11072 16046 11100 20334
rect 11256 17134 11284 27474
rect 12268 27443 12296 27474
rect 13924 24410 13952 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 13912 24404 13964 24410
rect 13912 24346 13964 24352
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 13372 23866 13400 24210
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15488 23866 15516 27520
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 13372 23322 13400 23802
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 13360 23316 13412 23322
rect 13360 23258 13412 23264
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13820 22976 13872 22982
rect 13820 22918 13872 22924
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 12992 22160 13044 22166
rect 12992 22102 13044 22108
rect 12544 21554 12572 22102
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12912 21690 12940 21966
rect 12900 21684 12952 21690
rect 12900 21626 12952 21632
rect 12912 21554 12940 21626
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12268 21078 12296 21286
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12268 20262 12296 20402
rect 11980 20256 12032 20262
rect 12256 20256 12308 20262
rect 12032 20216 12112 20244
rect 11980 20198 12032 20204
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 11348 19310 11376 19722
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 11532 19378 11560 19654
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11348 18834 11376 19246
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11348 18358 11376 18770
rect 11336 18352 11388 18358
rect 11336 18294 11388 18300
rect 11716 18222 11744 19450
rect 11900 18970 11928 19790
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11716 17882 11744 18158
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11348 16980 11376 17546
rect 11808 17270 11836 17750
rect 11992 17678 12020 19926
rect 12084 18222 12112 20216
rect 12176 20216 12256 20244
rect 12176 20058 12204 20216
rect 12256 20198 12308 20204
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12176 19174 12204 19994
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12176 18970 12204 19110
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12176 18086 12204 18906
rect 12268 18902 12296 19246
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11256 16952 11376 16980
rect 11256 16182 11284 16952
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11256 16046 11284 16118
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10796 15162 10824 15574
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10796 14550 10824 15098
rect 11072 14958 11100 15982
rect 11256 15706 11284 15982
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11348 15502 11376 16390
rect 11440 16114 11468 16390
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11992 15638 12020 17614
rect 12176 17066 12204 18022
rect 12360 17746 12388 20878
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12452 19718 12480 20334
rect 12624 20324 12676 20330
rect 12624 20266 12676 20272
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12544 18290 12572 18702
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12544 18086 12572 18226
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12636 17882 12664 20266
rect 12820 20058 12848 21286
rect 12912 21078 12940 21490
rect 13004 21350 13032 22102
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 12900 21072 12952 21078
rect 12900 21014 12952 21020
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12728 18970 12756 19178
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12636 17202 12664 17818
rect 12728 17814 12756 18158
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11440 15094 11468 15574
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10796 14006 10824 14486
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 11164 13938 11192 14350
rect 11440 14074 11468 14554
rect 11992 14414 12020 15574
rect 12268 15366 12296 16526
rect 12360 16250 12388 16594
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 15065 12296 15302
rect 12254 15056 12310 15065
rect 12254 14991 12310 15000
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 12360 14074 12388 16186
rect 12636 15910 12664 16458
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12544 14074 12572 15506
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11164 13814 11192 13874
rect 12360 13814 12388 14010
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12544 13814 12572 13874
rect 11164 13786 11284 13814
rect 12360 13786 12572 13814
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10152 12646 10180 13330
rect 11256 13190 11284 13786
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 10888 12714 10916 13126
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10244 11694 10272 12038
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11558 10732 11630
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10888 11354 10916 12650
rect 11164 12442 11192 12650
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10980 11626 11008 12174
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10980 11286 11008 11562
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10060 10674 10088 11086
rect 10244 10810 10272 11222
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10428 10742 10456 11154
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10324 10056 10376 10062
rect 10704 10044 10732 10406
rect 10888 10130 10916 11018
rect 11072 11014 11100 12310
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10324 9998 10376 10004
rect 10612 10016 10732 10044
rect 10336 9518 10364 9998
rect 10612 9518 10640 10016
rect 10888 9518 10916 10066
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10600 9512 10652 9518
rect 10876 9512 10928 9518
rect 10600 9454 10652 9460
rect 10704 9472 10876 9500
rect 9968 9042 9996 9454
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 9042 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9042 10732 9472
rect 10876 9454 10928 9460
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 9968 8090 9996 8978
rect 10152 8634 10180 8978
rect 10704 8634 10732 8978
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10060 7546 10088 8230
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10796 7886 10824 9318
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10980 8566 11008 8978
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 8090 11008 8230
rect 10968 8084 11020 8090
rect 11072 8072 11100 10950
rect 11152 10668 11204 10674
rect 11256 10656 11284 13126
rect 11624 12170 11652 13262
rect 11808 12986 11836 13398
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11900 12850 11928 13262
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11900 11898 11928 12582
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11992 11694 12020 12786
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12072 11756 12124 11762
rect 12176 11744 12204 12310
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12268 11830 12296 12242
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 12124 11716 12204 11744
rect 12072 11698 12124 11704
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11204 10628 11284 10656
rect 11152 10610 11204 10616
rect 11164 10198 11192 10610
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11348 9926 11376 11154
rect 11716 11082 11744 11494
rect 12176 11354 12204 11716
rect 12544 11354 12572 13786
rect 12636 13734 12664 15846
rect 12912 13784 12940 20402
rect 13188 18154 13216 22918
rect 13832 22574 13860 22918
rect 14568 22778 14596 23122
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 14280 22500 14332 22506
rect 14280 22442 14332 22448
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 13372 20602 13400 21014
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13464 19854 13492 20878
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13556 18970 13584 19858
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13648 18426 13676 21490
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13740 20330 13768 20878
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13740 20058 13768 20266
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13832 19972 13860 21966
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14200 21418 14228 21830
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 13912 19984 13964 19990
rect 13832 19944 13912 19972
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13188 17241 13216 18090
rect 13280 18086 13308 18294
rect 13268 18080 13320 18086
rect 13544 18080 13596 18086
rect 13268 18022 13320 18028
rect 13464 18040 13544 18068
rect 13174 17232 13230 17241
rect 13174 17167 13230 17176
rect 13280 15706 13308 18022
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 13004 14929 13032 15370
rect 12990 14920 13046 14929
rect 12990 14855 13046 14864
rect 13004 14822 13032 14855
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12728 13756 12940 13784
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 13462 12664 13670
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12636 12714 12664 13126
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12636 12442 12664 12650
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12728 12322 12756 13756
rect 12636 12294 12756 12322
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11808 10742 11836 10950
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11152 8084 11204 8090
rect 11072 8044 11152 8072
rect 10968 8026 11020 8032
rect 11152 8026 11204 8032
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10060 7274 10088 7482
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 5574 9904 6734
rect 9968 6322 9996 6870
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 10060 6254 10088 7210
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10796 7002 10824 7822
rect 10980 7410 11008 8026
rect 11164 7546 11192 8026
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10888 6798 10916 7210
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10888 1873 10916 2790
rect 11348 2514 11376 9862
rect 11440 8838 11468 9930
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11440 3194 11468 8774
rect 11532 8090 11560 9454
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11532 6458 11560 6734
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11624 2961 11652 8230
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11716 7342 11744 7686
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11716 6934 11744 7278
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11716 6322 11744 6870
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11610 2952 11666 2961
rect 11610 2887 11666 2896
rect 11808 2553 11836 10678
rect 12176 10266 12204 11290
rect 12544 10606 12572 11290
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12544 10266 12572 10542
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11900 9625 11928 10066
rect 11886 9616 11942 9625
rect 11886 9551 11942 9560
rect 11900 9518 11928 9551
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11900 9110 11928 9454
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12360 9178 12388 9386
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 12360 8498 12388 9114
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12360 7954 12388 8434
rect 12452 8022 12480 9318
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12176 6934 12204 7754
rect 12452 7002 12480 7958
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12636 6225 12664 12294
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12820 10130 12848 11630
rect 13004 11218 13032 14758
rect 13096 14618 13124 15506
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13096 14385 13124 14554
rect 13176 14408 13228 14414
rect 13082 14376 13138 14385
rect 13176 14350 13228 14356
rect 13082 14311 13138 14320
rect 13096 12646 13124 14311
rect 13188 13530 13216 14350
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13280 13394 13308 14894
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12782 13216 13126
rect 13372 12782 13400 14010
rect 13464 13462 13492 18040
rect 13544 18022 13596 18028
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13556 16726 13584 17682
rect 13648 17610 13676 18362
rect 13740 18358 13768 19654
rect 13832 19514 13860 19944
rect 13912 19926 13964 19932
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 14016 18970 14044 19790
rect 14108 19242 14136 20810
rect 14200 19786 14228 21354
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 14108 18902 14136 19178
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 14292 17202 14320 22442
rect 14660 21010 14688 23462
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14660 20602 14688 20946
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14476 19514 14504 20198
rect 14740 19780 14792 19786
rect 14740 19722 14792 19728
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14384 18426 14412 18770
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14384 18086 14412 18362
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14660 17882 14688 18022
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14476 17270 14504 17750
rect 14752 17338 14780 19722
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13452 13456 13504 13462
rect 13556 13433 13584 14894
rect 13648 14822 13676 17002
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16726 13860 16934
rect 14292 16794 14320 17138
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13648 14618 13676 14758
rect 13740 14618 13768 15914
rect 13832 15706 13860 16662
rect 14188 16584 14240 16590
rect 14240 16544 14320 16572
rect 14188 16526 14240 16532
rect 14292 16046 14320 16544
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15706 14320 15982
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14660 14618 14688 14894
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 13648 14074 13676 14554
rect 14384 14278 14412 14554
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 14074 14412 14214
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14384 13734 14412 14010
rect 14752 13938 14780 14758
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 13452 13398 13504 13404
rect 13542 13424 13598 13433
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13188 12102 13216 12718
rect 13372 12374 13400 12718
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13372 11218 13400 12310
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13004 10606 13032 11154
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12728 9586 12756 9862
rect 12820 9722 12848 10066
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12728 8566 12756 9522
rect 12820 9178 12848 9658
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12820 8566 12848 9114
rect 13004 9042 13032 10542
rect 13464 10033 13492 13398
rect 13542 13359 13598 13368
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 12918 13676 13330
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14384 12986 14412 13262
rect 14660 13258 14688 13738
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13556 11694 13584 12038
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13556 10112 13584 11630
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13648 10606 13676 11154
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13636 10124 13688 10130
rect 13556 10084 13636 10112
rect 13636 10066 13688 10072
rect 13450 10024 13506 10033
rect 13450 9959 13506 9968
rect 13648 9722 13676 10066
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13740 9518 13768 12038
rect 13832 11830 13860 12378
rect 14016 12238 14044 12650
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14016 11898 14044 12174
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 14108 11694 14136 12718
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14384 12102 14412 12242
rect 14476 12238 14504 13194
rect 14844 12850 14872 22374
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20466 15332 21354
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15304 20058 15332 20402
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 18630 15332 19790
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15396 18154 15424 22714
rect 16132 22438 16160 23122
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 15476 19984 15528 19990
rect 15476 19926 15528 19932
rect 15488 19514 15516 19926
rect 15580 19514 15608 21966
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15672 20330 15700 20742
rect 15660 20324 15712 20330
rect 15660 20266 15712 20272
rect 15672 19990 15700 20266
rect 15856 20262 15884 21898
rect 15948 21690 15976 21898
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 16500 21554 16528 21830
rect 17052 21622 17080 21966
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 17144 21554 17172 27520
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18064 23322 18092 23598
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 18800 22234 18828 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20456 23866 20484 27520
rect 22112 23866 22140 27520
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 22100 23860 22152 23866
rect 22100 23802 22152 23808
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 21284 22778 21312 23598
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15948 19718 15976 21286
rect 16500 21146 16528 21490
rect 16856 21412 16908 21418
rect 16856 21354 16908 21360
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 16684 20602 16712 20878
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 16684 20058 16712 20538
rect 16776 20466 16804 21014
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16776 19990 16804 20402
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 15948 19514 15976 19654
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15488 19174 15516 19450
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15948 18902 15976 19450
rect 16040 19242 16068 19926
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16592 18970 16620 19178
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 15948 18426 15976 18838
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 14924 18148 14976 18154
rect 14924 18090 14976 18096
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15660 18148 15712 18154
rect 15660 18090 15712 18096
rect 14936 17882 14964 18090
rect 14924 17876 14976 17882
rect 14924 17818 14976 17824
rect 15476 17808 15528 17814
rect 15476 17750 15528 17756
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16182 15332 16526
rect 15396 16522 15424 17614
rect 15488 17338 15516 17750
rect 15672 17678 15700 18090
rect 16408 17882 16436 18294
rect 16500 18086 16528 18566
rect 16868 18426 16896 21354
rect 17144 20466 17172 21490
rect 17420 21350 17448 22102
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 19168 21554 19196 22034
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 18144 21480 18196 21486
rect 19168 21457 19196 21490
rect 18144 21422 18196 21428
rect 19154 21448 19210 21457
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17420 21078 17448 21286
rect 17408 21072 17460 21078
rect 17408 21014 17460 21020
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 17224 19984 17276 19990
rect 17224 19926 17276 19932
rect 17236 19514 17264 19926
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17328 19394 17356 20198
rect 17420 19446 17448 20334
rect 17604 19854 17632 20878
rect 18052 20800 18104 20806
rect 18156 20788 18184 21422
rect 18788 21412 18840 21418
rect 19154 21383 19210 21392
rect 18788 21354 18840 21360
rect 18800 21146 18828 21354
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 18788 21140 18840 21146
rect 18788 21082 18840 21088
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18104 20760 18184 20788
rect 18052 20742 18104 20748
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17236 19366 17356 19394
rect 17408 19440 17460 19446
rect 17408 19382 17460 19388
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16764 18216 16816 18222
rect 16868 18204 16896 18362
rect 16816 18176 16896 18204
rect 16764 18158 16816 18164
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15476 16720 15528 16726
rect 15672 16708 15700 17614
rect 15528 16680 15700 16708
rect 16120 16720 16172 16726
rect 15476 16662 15528 16668
rect 16120 16662 16172 16668
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 16132 16182 16160 16662
rect 15292 16176 15344 16182
rect 16120 16176 16172 16182
rect 15292 16118 15344 16124
rect 15842 16144 15898 16153
rect 16120 16118 16172 16124
rect 15842 16079 15898 16088
rect 15856 16046 15884 16079
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15638 15700 15846
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15672 14618 15700 15574
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15568 13524 15620 13530
rect 15672 13512 15700 14350
rect 15764 14074 15792 14486
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15856 14006 15884 15438
rect 16224 15434 16252 17818
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16776 17202 16804 17478
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16316 16454 16344 16934
rect 16592 16522 16620 17002
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16316 15910 16344 16390
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 16224 13938 16252 15370
rect 16408 15366 16436 15914
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 15844 13864 15896 13870
rect 16316 13814 16344 14214
rect 15844 13806 15896 13812
rect 15620 13484 15700 13512
rect 15568 13466 15620 13472
rect 15672 13433 15700 13484
rect 15658 13424 15714 13433
rect 15384 13388 15436 13394
rect 15658 13359 15714 13368
rect 15384 13330 15436 13336
rect 15396 13297 15424 13330
rect 15856 13326 15884 13806
rect 16224 13802 16344 13814
rect 16408 13802 16436 15030
rect 16500 14958 16528 15098
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16488 14408 16540 14414
rect 16592 14396 16620 16458
rect 16776 16250 16804 17138
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16868 15162 16896 18176
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 17052 16114 17080 16458
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16540 14368 16620 14396
rect 16488 14350 16540 14356
rect 16500 13938 16528 14350
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 17236 13814 17264 19366
rect 17512 19174 17540 19790
rect 18064 19334 18092 20742
rect 18248 20262 18276 20946
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20330 18736 20742
rect 18800 20466 18828 21082
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18696 20324 18748 20330
rect 18696 20266 18748 20272
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18708 19990 18736 20266
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18616 19514 18644 19790
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 17972 19306 18092 19334
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17512 18426 17540 19110
rect 17972 18834 18000 19306
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17696 18154 17724 18770
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17328 15910 17356 16662
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 15094 17356 15846
rect 17316 15088 17368 15094
rect 17316 15030 17368 15036
rect 17420 14482 17448 17546
rect 17512 17338 17540 17682
rect 17696 17338 17724 18090
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17420 14074 17448 14418
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 16212 13796 16344 13802
rect 16264 13786 16344 13796
rect 16396 13796 16448 13802
rect 16212 13738 16264 13744
rect 17236 13786 17356 13814
rect 16396 13738 16448 13744
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15568 13320 15620 13326
rect 15382 13288 15438 13297
rect 15568 13262 15620 13268
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15382 13223 15438 13232
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15580 12986 15608 13262
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 16040 12918 16068 13466
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 13832 10130 13860 11630
rect 14108 11218 14136 11630
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14384 11218 14412 11562
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14108 10792 14136 11154
rect 14188 10804 14240 10810
rect 14108 10764 14188 10792
rect 14188 10746 14240 10752
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10130 14136 10406
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14108 9586 14136 10066
rect 14200 9654 14228 10746
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13004 8634 13032 8978
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12820 8430 12848 8502
rect 13004 8430 13032 8570
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12728 7410 12756 7958
rect 13096 7546 13124 8570
rect 13740 8430 13768 8978
rect 14108 8430 14136 9522
rect 14200 9042 14228 9590
rect 14660 9586 14688 12582
rect 15028 12442 15056 12650
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14844 11286 14872 11766
rect 15304 11762 15332 12378
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15396 11354 15424 12174
rect 15488 11898 15516 12310
rect 15672 12238 15700 12786
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14844 10810 14872 11222
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14844 10538 14872 10746
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 15028 10198 15056 10542
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15016 10192 15068 10198
rect 15016 10134 15068 10140
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 15580 9178 15608 10474
rect 15672 10266 15700 11154
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 13556 8090 13584 8366
rect 14844 8090 14872 8910
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15580 8634 15608 9114
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15212 8090 15240 8366
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15488 8022 15516 8434
rect 15580 8294 15608 8570
rect 15948 8430 15976 12582
rect 16224 11354 16252 13738
rect 16408 13530 16436 13738
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16396 12096 16448 12102
rect 16500 12073 16528 12718
rect 16684 12442 16712 12922
rect 17052 12646 17080 13330
rect 17328 12714 17356 13786
rect 17512 13190 17540 17274
rect 17590 17232 17646 17241
rect 17788 17218 17816 18226
rect 17972 17746 18000 18770
rect 18248 17814 18276 19110
rect 18616 18902 18644 19450
rect 18708 19378 18736 19926
rect 18892 19786 18920 20742
rect 19536 20262 19564 21014
rect 19996 20942 20024 21286
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 19812 20466 19840 20810
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19536 20058 19564 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19996 20058 20024 20878
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18708 19242 18736 19314
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18708 18970 18736 19178
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 18708 18426 18736 18906
rect 19352 18766 19380 19654
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19444 18902 19472 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19996 18902 20024 19314
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 19076 18154 19104 18362
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18236 17808 18288 17814
rect 18708 17785 18736 18022
rect 18236 17750 18288 17756
rect 18694 17776 18750 17785
rect 17960 17740 18012 17746
rect 18694 17711 18750 17720
rect 17960 17682 18012 17688
rect 17590 17167 17646 17176
rect 17696 17190 17816 17218
rect 17604 15162 17632 17167
rect 17696 16561 17724 17190
rect 17972 16794 18000 17682
rect 19260 17610 19288 18158
rect 19352 17882 19380 18702
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 19064 17604 19116 17610
rect 19064 17546 19116 17552
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19076 17338 19104 17546
rect 19536 17338 19564 17682
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19628 17202 19656 17614
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17776 16584 17828 16590
rect 17682 16552 17738 16561
rect 17776 16526 17828 16532
rect 17682 16487 17738 16496
rect 17696 15570 17724 16487
rect 17788 16114 17816 16526
rect 18248 16454 18276 17070
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17788 16017 17816 16050
rect 17774 16008 17830 16017
rect 17774 15943 17830 15952
rect 18248 15570 18276 16390
rect 18800 16250 18828 17002
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18892 16182 18920 16934
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20272 16794 20300 17138
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18892 15978 18920 16118
rect 19444 16046 19472 16662
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 17684 15564 17736 15570
rect 18236 15564 18288 15570
rect 17736 15524 17816 15552
rect 17684 15506 17736 15512
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17604 14482 17632 14826
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 14074 17632 14418
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16396 12038 16448 12044
rect 16486 12064 16542 12073
rect 16408 11626 16436 12038
rect 16486 11999 16542 12008
rect 16960 11830 16988 12174
rect 17328 11830 17356 12310
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16408 10810 16436 11562
rect 16960 11014 16988 11766
rect 17328 11218 17356 11766
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16026 10704 16082 10713
rect 16026 10639 16082 10648
rect 16040 10266 16068 10639
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16040 9586 16068 10202
rect 16408 10198 16436 10542
rect 16960 10198 16988 10950
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16316 9654 16344 9998
rect 16408 9722 16436 10134
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 8634 16160 9318
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 16132 8022 16160 8570
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 16120 8016 16172 8022
rect 16120 7958 16172 7964
rect 13542 7848 13598 7857
rect 13452 7812 13504 7818
rect 13504 7792 13542 7800
rect 13504 7783 13598 7792
rect 13504 7772 13584 7783
rect 13452 7754 13504 7760
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 16132 7546 16160 7958
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 16132 7342 16160 7482
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 16408 6254 16436 7822
rect 16592 7410 16620 8230
rect 16960 7993 16988 8366
rect 17144 8362 17172 8910
rect 17236 8430 17264 9046
rect 17328 8974 17356 9386
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 16946 7984 17002 7993
rect 16946 7919 17002 7928
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 17328 7206 17356 7822
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 16396 6248 16448 6254
rect 12622 6216 12678 6225
rect 17328 6225 17356 7142
rect 16396 6190 16448 6196
rect 17314 6216 17370 6225
rect 12622 6151 12678 6160
rect 17314 6151 17370 6160
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 17420 4154 17448 12854
rect 17512 12374 17540 13126
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17512 10606 17540 11154
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17512 9722 17540 10066
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17512 8090 17540 8298
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17604 7993 17632 8230
rect 17590 7984 17646 7993
rect 17590 7919 17646 7928
rect 17236 4126 17448 4154
rect 16118 4040 16174 4049
rect 16118 3975 16174 3984
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15474 2952 15530 2961
rect 15474 2887 15530 2896
rect 11794 2544 11850 2553
rect 11336 2508 11388 2514
rect 15488 2514 15516 2887
rect 11794 2479 11850 2488
rect 15476 2508 15528 2514
rect 11336 2450 11388 2456
rect 15476 2450 15528 2456
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 10874 1864 10930 1873
rect 10874 1799 10930 1808
rect 9034 54 9168 82
rect 9680 128 9732 134
rect 9680 70 9732 76
rect 10414 128 10470 480
rect 10414 76 10416 128
rect 10468 76 10470 128
rect 9034 0 9090 54
rect 10414 0 10470 76
rect 11794 82 11850 480
rect 11900 82 11928 2314
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 11794 54 11928 82
rect 13004 82 13032 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 13174 82 13230 480
rect 13004 54 13230 82
rect 11794 0 11850 54
rect 13174 0 13230 54
rect 14646 128 14702 480
rect 14646 76 14648 128
rect 14700 76 14702 128
rect 14646 0 14702 76
rect 16026 82 16082 480
rect 16132 82 16160 3975
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16408 2553 16436 2586
rect 16394 2544 16450 2553
rect 16394 2479 16450 2488
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 16026 54 16160 82
rect 17144 82 17172 2314
rect 17236 202 17264 4126
rect 17696 2514 17724 15302
rect 17788 14822 17816 15524
rect 18236 15506 18288 15512
rect 18248 14890 18276 15506
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 18524 14482 18552 15438
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18800 14618 18828 14826
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18800 13938 18828 14554
rect 18892 14550 18920 15914
rect 18984 15366 19012 15982
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19996 15706 20024 16526
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18984 15026 19012 15302
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18892 13734 18920 14486
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18432 13530 18460 13670
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17788 11778 17816 12650
rect 17880 12646 17908 13262
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17880 12442 17908 12582
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 18248 12374 18276 12718
rect 18432 12646 18460 13466
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 17788 11750 17908 11778
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17788 10198 17816 11562
rect 17880 10713 17908 11750
rect 18144 11620 18196 11626
rect 18064 11580 18144 11608
rect 18064 11014 18092 11580
rect 18144 11562 18196 11568
rect 18432 11286 18460 12582
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 17866 10704 17922 10713
rect 18064 10674 18092 10950
rect 17866 10639 17922 10648
rect 18052 10668 18104 10674
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9178 17816 9318
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17788 7954 17816 9114
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17880 2582 17908 10639
rect 18052 10610 18104 10616
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 17224 196 17276 202
rect 17224 138 17276 144
rect 17406 82 17462 480
rect 17972 134 18000 10542
rect 18156 9654 18184 10950
rect 18432 10538 18460 11222
rect 18524 11218 18552 12854
rect 19076 12646 19104 13126
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 19260 12306 19288 14894
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 20260 14544 20312 14550
rect 20260 14486 20312 14492
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19904 14006 19932 14418
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 19892 14000 19944 14006
rect 19892 13942 19944 13948
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20180 13530 20208 14282
rect 20272 14006 20300 14486
rect 20260 14000 20312 14006
rect 20260 13942 20312 13948
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19444 12850 19472 13398
rect 20180 12850 20208 13466
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18616 11937 18644 12106
rect 18602 11928 18658 11937
rect 18602 11863 18658 11872
rect 18800 11762 18828 12174
rect 19076 11898 19104 12242
rect 19260 11898 19288 12242
rect 20364 12186 20392 22374
rect 21468 22234 21496 22918
rect 21640 22432 21692 22438
rect 21640 22374 21692 22380
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20548 20058 20576 20402
rect 20640 20330 20668 21286
rect 20916 21078 20944 21966
rect 21468 21554 21496 22170
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21560 21434 21588 21490
rect 21468 21406 21588 21434
rect 20904 21072 20956 21078
rect 20904 21014 20956 21020
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20824 20466 20852 20810
rect 20916 20602 20944 21014
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20628 20324 20680 20330
rect 20628 20266 20680 20272
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20640 19514 20668 19790
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20548 18358 20576 19110
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20732 17882 20760 18702
rect 20824 18698 20852 20402
rect 21376 20262 21404 21014
rect 21468 20942 21496 21406
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21468 20516 21496 20878
rect 21548 20528 21600 20534
rect 21468 20488 21548 20516
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21376 19990 21404 20198
rect 21364 19984 21416 19990
rect 21364 19926 21416 19932
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20824 17678 20852 18634
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21192 18222 21220 18566
rect 21284 18426 21312 19178
rect 21468 18766 21496 20488
rect 21548 20470 21600 20476
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 21100 17814 21128 18022
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20456 16726 20484 17138
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16794 20760 16934
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20444 16720 20496 16726
rect 20824 16708 20852 17614
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20904 16720 20956 16726
rect 20824 16680 20904 16708
rect 20444 16662 20496 16668
rect 20904 16662 20956 16668
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20456 15026 20484 15302
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20536 14884 20588 14890
rect 20536 14826 20588 14832
rect 20548 14618 20576 14826
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 21008 14414 21036 17138
rect 21100 17066 21128 17750
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 21652 16998 21680 22374
rect 22376 22092 22428 22098
rect 22376 22034 22428 22040
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22204 21146 22232 21830
rect 22388 21690 22416 22034
rect 23768 21690 23796 27520
rect 25226 25664 25282 25673
rect 25226 25599 25282 25608
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 25148 22710 25176 23122
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 23940 22160 23992 22166
rect 23940 22102 23992 22108
rect 23952 21690 23980 22102
rect 25240 22098 25268 25599
rect 25424 22166 25452 27520
rect 27066 27532 27122 28000
rect 27066 27520 27068 27532
rect 26240 27474 26292 27480
rect 27120 27520 27122 27532
rect 27068 27474 27120 27480
rect 25502 23488 25558 23497
rect 25502 23423 25558 23432
rect 25516 22778 25544 23423
rect 25504 22772 25556 22778
rect 25504 22714 25556 22720
rect 25516 22574 25544 22714
rect 25504 22568 25556 22574
rect 25504 22510 25556 22516
rect 25502 22264 25558 22273
rect 25502 22199 25558 22208
rect 25412 22160 25464 22166
rect 25412 22102 25464 22108
rect 24676 22092 24728 22098
rect 24676 22034 24728 22040
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22008 20868 22060 20874
rect 22008 20810 22060 20816
rect 22020 19922 22048 20810
rect 22204 20466 22232 21082
rect 22848 21078 22876 21286
rect 22836 21072 22888 21078
rect 22836 21014 22888 21020
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22756 20602 22784 20878
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22848 20534 22876 21014
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22284 20324 22336 20330
rect 22284 20266 22336 20272
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22020 19378 22048 19858
rect 22112 19514 22140 19926
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22008 19236 22060 19242
rect 22008 19178 22060 19184
rect 22020 18698 22048 19178
rect 22296 18902 22324 20266
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22848 19174 22876 19858
rect 23124 19854 23152 20198
rect 23400 20058 23428 20538
rect 24044 20369 24072 21830
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21690 24716 22034
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 25134 21040 25190 21049
rect 25516 21010 25544 22199
rect 25134 20975 25190 20984
rect 25504 21004 25556 21010
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 25148 20602 25176 20975
rect 25504 20946 25556 20952
rect 25516 20602 25544 20946
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 25148 20398 25176 20538
rect 25136 20392 25188 20398
rect 24030 20360 24086 20369
rect 25136 20334 25188 20340
rect 24030 20295 24086 20304
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 24216 19916 24268 19922
rect 24216 19858 24268 19864
rect 23112 19848 23164 19854
rect 23018 19816 23074 19825
rect 23112 19790 23164 19796
rect 23018 19751 23074 19760
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22192 18896 22244 18902
rect 22192 18838 22244 18844
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 22020 17610 22048 18634
rect 22204 18086 22232 18838
rect 22296 18358 22324 18838
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22284 18352 22336 18358
rect 22284 18294 22336 18300
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22008 17604 22060 17610
rect 22008 17546 22060 17552
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21928 17066 21956 17478
rect 22204 17270 22232 18022
rect 22572 17882 22600 18158
rect 22664 18086 22692 18702
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22664 17882 22692 18022
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22848 17785 22876 19110
rect 22834 17776 22890 17785
rect 22468 17740 22520 17746
rect 22834 17711 22890 17720
rect 22928 17740 22980 17746
rect 22468 17682 22520 17688
rect 22928 17682 22980 17688
rect 22192 17264 22244 17270
rect 22480 17241 22508 17682
rect 22940 17338 22968 17682
rect 22928 17332 22980 17338
rect 22928 17274 22980 17280
rect 22192 17206 22244 17212
rect 22466 17232 22522 17241
rect 22466 17167 22522 17176
rect 22480 17134 22508 17167
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 21916 17060 21968 17066
rect 21916 17002 21968 17008
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21548 16516 21600 16522
rect 21548 16458 21600 16464
rect 21180 15972 21232 15978
rect 21180 15914 21232 15920
rect 21192 15638 21220 15914
rect 21180 15632 21232 15638
rect 21180 15574 21232 15580
rect 21192 15162 21220 15574
rect 21560 15502 21588 16458
rect 21652 16046 21680 16662
rect 21928 16250 21956 17002
rect 23032 16658 23060 19751
rect 24228 19446 24256 19858
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 24228 19174 24256 19382
rect 24216 19168 24268 19174
rect 24216 19110 24268 19116
rect 23112 18896 23164 18902
rect 23112 18838 23164 18844
rect 23124 18426 23152 18838
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23768 17678 23796 18022
rect 24044 17746 24072 18158
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22388 16250 22416 16390
rect 23032 16250 23060 16594
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21652 15910 21680 15982
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21928 15638 21956 16186
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 21824 15564 21876 15570
rect 21744 15524 21824 15552
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21272 14884 21324 14890
rect 21272 14826 21324 14832
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 20456 13938 20484 14350
rect 21100 14074 21128 14486
rect 21284 14414 21312 14826
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20456 13530 20484 13874
rect 20536 13796 20588 13802
rect 20536 13738 20588 13744
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20548 13462 20576 13738
rect 20536 13456 20588 13462
rect 20536 13398 20588 13404
rect 20720 13456 20772 13462
rect 20720 13398 20772 13404
rect 20732 12986 20760 13398
rect 21284 13258 21312 14350
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13462 21404 13670
rect 21364 13456 21416 13462
rect 21364 13398 21416 13404
rect 21456 13320 21508 13326
rect 21560 13308 21588 15438
rect 21744 15162 21772 15524
rect 21824 15506 21876 15512
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21744 15065 21772 15098
rect 21730 15056 21786 15065
rect 21730 14991 21786 15000
rect 21928 14872 21956 15574
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22204 15026 22232 15302
rect 22836 15088 22888 15094
rect 22836 15030 22888 15036
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22008 14884 22060 14890
rect 21928 14844 22008 14872
rect 21928 14618 21956 14844
rect 22008 14826 22060 14832
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22112 13734 22140 14350
rect 22756 14074 22784 14826
rect 22848 14414 22876 15030
rect 22940 14929 22968 15370
rect 22926 14920 22982 14929
rect 22926 14855 22982 14864
rect 22940 14822 22968 14855
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 23032 14550 23060 15846
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23112 15496 23164 15502
rect 23112 15438 23164 15444
rect 23020 14544 23072 14550
rect 23020 14486 23072 14492
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22756 13870 22784 14010
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22112 13530 22140 13670
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22204 13433 22232 13670
rect 22652 13456 22704 13462
rect 22190 13424 22246 13433
rect 22652 13398 22704 13404
rect 22190 13359 22246 13368
rect 21508 13280 21588 13308
rect 21456 13262 21508 13268
rect 21272 13252 21324 13258
rect 21272 13194 21324 13200
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21376 12714 21404 12922
rect 21560 12714 21588 13280
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21916 12708 21968 12714
rect 21916 12650 21968 12656
rect 22008 12708 22060 12714
rect 22008 12650 22060 12656
rect 20904 12232 20956 12238
rect 20364 12158 20484 12186
rect 20904 12174 20956 12180
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18800 11665 18828 11698
rect 20364 11694 20392 12038
rect 20352 11688 20404 11694
rect 18786 11656 18842 11665
rect 20352 11630 20404 11636
rect 18786 11591 18842 11600
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18432 10266 18460 10474
rect 19168 10266 19196 11086
rect 20180 10810 20208 11494
rect 20364 11286 20392 11630
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20456 11082 20484 12158
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20180 10470 20208 10746
rect 20916 10674 20944 12174
rect 21284 12170 21312 12650
rect 21928 12442 21956 12650
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 22020 11801 22048 12650
rect 22572 12442 22600 13262
rect 22664 12986 22692 13398
rect 22848 13326 22876 14350
rect 23032 14074 23060 14486
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 22836 13320 22888 13326
rect 23124 13297 23152 15438
rect 23308 14822 23336 15506
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23308 14385 23336 14758
rect 23294 14376 23350 14385
rect 23294 14311 23350 14320
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 22836 13262 22888 13268
rect 23110 13288 23166 13297
rect 23110 13223 23166 13232
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 23400 12918 23428 13806
rect 23388 12912 23440 12918
rect 23388 12854 23440 12860
rect 23754 12880 23810 12889
rect 23754 12815 23810 12824
rect 23204 12708 23256 12714
rect 23204 12650 23256 12656
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22848 12442 22876 12582
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22836 12436 22888 12442
rect 22836 12378 22888 12384
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 22006 11792 22062 11801
rect 22006 11727 22062 11736
rect 22296 11558 22324 12242
rect 23032 11558 23060 12242
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 21456 11280 21508 11286
rect 21456 11222 21508 11228
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21100 10742 21128 11018
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18984 9450 19012 9658
rect 18972 9444 19024 9450
rect 18972 9386 19024 9392
rect 18420 9104 18472 9110
rect 18420 9046 18472 9052
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8566 18092 8774
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 18432 8498 18460 9046
rect 18984 8974 19012 9386
rect 19444 9382 19472 10066
rect 19536 9450 19564 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 20548 10266 20576 10610
rect 21284 10538 21312 11086
rect 21468 10810 21496 11222
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19996 9586 20024 9862
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18432 8022 18460 8434
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18248 7546 18276 7890
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18892 4049 18920 8774
rect 19076 8294 19104 9046
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19076 8022 19104 8230
rect 19064 8016 19116 8022
rect 19064 7958 19116 7964
rect 19444 5681 19472 9318
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 9178 20024 9386
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19522 8936 19578 8945
rect 21008 8906 21036 9998
rect 21100 9586 21128 10134
rect 21284 10062 21312 10474
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 22006 10024 22062 10033
rect 21284 9654 21312 9998
rect 22006 9959 22062 9968
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 19522 8871 19578 8880
rect 20996 8900 21048 8906
rect 19430 5672 19486 5681
rect 19430 5607 19486 5616
rect 19444 5166 19472 5607
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 18878 4040 18934 4049
rect 18878 3975 18934 3984
rect 17144 54 17462 82
rect 17960 128 18012 134
rect 17960 70 18012 76
rect 18786 128 18842 480
rect 19536 134 19564 8871
rect 20996 8842 21048 8848
rect 21836 8566 21864 9522
rect 21824 8560 21876 8566
rect 21824 8502 21876 8508
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 18786 76 18788 128
rect 18840 76 18842 128
rect 16026 0 16082 54
rect 17406 0 17462 54
rect 18786 0 18842 76
rect 19524 128 19576 134
rect 19524 70 19576 76
rect 20166 128 20222 480
rect 20166 76 20168 128
rect 20220 76 20222 128
rect 20166 0 20222 76
rect 21376 82 21404 6326
rect 22020 1193 22048 9959
rect 22296 8838 22324 11494
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22848 10810 22876 11154
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22848 10713 22876 10746
rect 22834 10704 22890 10713
rect 22834 10639 22890 10648
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22480 10033 22508 10542
rect 22466 10024 22522 10033
rect 22466 9959 22522 9968
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 23216 7954 23244 12650
rect 23768 11937 23796 12815
rect 23754 11928 23810 11937
rect 23754 11863 23810 11872
rect 23572 11552 23624 11558
rect 23572 11494 23624 11500
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23308 9586 23336 9998
rect 23400 9722 23428 10066
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 22742 1864 22798 1873
rect 22742 1799 22798 1808
rect 22006 1184 22062 1193
rect 22006 1119 22062 1128
rect 21638 82 21694 480
rect 21376 54 21694 82
rect 22756 82 22784 1799
rect 23018 82 23074 480
rect 23584 134 23612 11494
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23768 8294 23796 8978
rect 23756 8288 23808 8294
rect 23756 8230 23808 8236
rect 23768 7857 23796 8230
rect 23754 7848 23810 7857
rect 23754 7783 23810 7792
rect 23860 4078 23888 17614
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 24044 17338 24072 17478
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23952 16250 23980 16594
rect 23940 16244 23992 16250
rect 23940 16186 23992 16192
rect 23952 16153 23980 16186
rect 23938 16144 23994 16153
rect 23938 16079 23994 16088
rect 24044 16017 24072 16934
rect 24228 16153 24256 19110
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 25228 17740 25280 17746
rect 25228 17682 25280 17688
rect 24950 17504 25006 17513
rect 24289 17436 24585 17456
rect 24950 17439 25006 17448
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24766 16416 24822 16425
rect 24289 16348 24585 16368
rect 24766 16351 24822 16360
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24214 16144 24270 16153
rect 24214 16079 24270 16088
rect 24030 16008 24086 16017
rect 24030 15943 24086 15952
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 23952 12306 23980 13194
rect 24044 12646 24072 15846
rect 24780 15706 24808 16351
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24136 14958 24164 15506
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24032 12640 24084 12646
rect 24032 12582 24084 12588
rect 23940 12300 23992 12306
rect 23940 12242 23992 12248
rect 23952 11898 23980 12242
rect 24136 12186 24164 14894
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24228 12986 24256 13330
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24964 12986 24992 17439
rect 25240 16998 25268 17682
rect 26252 17338 26280 27474
rect 27080 27443 27108 27474
rect 26790 26888 26846 26897
rect 26790 26823 26846 26832
rect 26804 21457 26832 26823
rect 27618 25120 27674 25129
rect 27618 25055 27674 25064
rect 27632 22710 27660 25055
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 26790 21448 26846 21457
rect 26790 21383 26846 21392
rect 27618 19272 27674 19281
rect 27618 19207 27674 19216
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 24228 12714 24256 12922
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 24216 12708 24268 12714
rect 24216 12650 24268 12656
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24044 12158 24164 12186
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 24044 10266 24072 12158
rect 24122 12064 24178 12073
rect 24122 11999 24178 12008
rect 24136 11694 24164 11999
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24124 11688 24176 11694
rect 24124 11630 24176 11636
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9722 24716 12582
rect 25148 12442 25176 12718
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 24766 11928 24822 11937
rect 24766 11863 24822 11872
rect 24780 11830 24808 11863
rect 24768 11824 24820 11830
rect 24768 11766 24820 11772
rect 24766 10568 24822 10577
rect 24766 10503 24822 10512
rect 24780 10266 24808 10503
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 25240 10198 25268 16934
rect 27632 15910 27660 19207
rect 27620 15904 27672 15910
rect 27620 15846 27672 15852
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27632 14657 27660 14758
rect 27618 14648 27674 14657
rect 27618 14583 27674 14592
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25516 11762 25544 12242
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25516 11665 25544 11698
rect 25502 11656 25558 11665
rect 25502 11591 25558 11600
rect 25228 10192 25280 10198
rect 25228 10134 25280 10140
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25148 9722 25176 10066
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 24674 9344 24730 9353
rect 24412 9178 24440 9318
rect 24674 9279 24730 9288
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 24688 9042 24716 9279
rect 24766 9208 24822 9217
rect 24766 9143 24822 9152
rect 24676 9036 24728 9042
rect 24676 8978 24728 8984
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24688 8634 24716 8978
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7546 24716 7890
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24780 6866 24808 9143
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 27632 7585 27660 7686
rect 27618 7576 27674 7585
rect 27618 7511 27674 7520
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24780 6458 24808 6802
rect 27620 6656 27672 6662
rect 27620 6598 27672 6604
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 27632 6361 27660 6598
rect 27618 6352 27674 6361
rect 27618 6287 27674 6296
rect 24858 6216 24914 6225
rect 24858 6151 24914 6160
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24596 5817 24624 5850
rect 24582 5808 24638 5817
rect 24582 5743 24638 5752
rect 24766 5536 24822 5545
rect 24289 5468 24585 5488
rect 24766 5471 24822 5480
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24780 5370 24808 5471
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24872 3194 24900 6151
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25240 5030 25268 5714
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 25240 3233 25268 4966
rect 27620 4208 27672 4214
rect 27620 4150 27672 4156
rect 27632 4049 27660 4150
rect 27618 4040 27674 4049
rect 27618 3975 27674 3984
rect 25226 3224 25282 3233
rect 24860 3188 24912 3194
rect 25226 3159 25282 3168
rect 24860 3130 24912 3136
rect 25136 2848 25188 2854
rect 25136 2790 25188 2796
rect 25148 2281 25176 2790
rect 25412 2576 25464 2582
rect 25412 2518 25464 2524
rect 25134 2272 25190 2281
rect 24289 2204 24585 2224
rect 25134 2207 25190 2216
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 22756 54 23074 82
rect 23572 128 23624 134
rect 23572 70 23624 76
rect 24398 128 24454 480
rect 24398 76 24400 128
rect 24452 76 24454 128
rect 21638 0 21694 54
rect 23018 0 23074 54
rect 24398 0 24454 76
rect 25424 82 25452 2518
rect 26884 2304 26936 2310
rect 26884 2246 26936 2252
rect 25778 82 25834 480
rect 25424 54 25834 82
rect 26896 82 26924 2246
rect 27158 82 27214 480
rect 26896 54 27214 82
rect 25778 0 25834 54
rect 27158 0 27214 54
<< via2 >>
rect 1030 22888 1086 22944
rect 18 15816 74 15872
rect 1490 26832 1546 26888
rect 1582 21664 1638 21720
rect 1582 20304 1638 20360
rect 110 14592 166 14648
rect 1122 13504 1178 13560
rect 110 12008 166 12064
rect 1674 19080 1730 19136
rect 1858 24384 1914 24440
rect 1858 19216 1914 19272
rect 1582 10104 1638 10160
rect 2778 17584 2834 17640
rect 5262 25472 5318 25528
rect 3698 15000 3754 15056
rect 1582 5072 1638 5128
rect 1674 4020 1676 4040
rect 1676 4020 1728 4040
rect 1728 4020 1730 4040
rect 1674 3984 1730 4020
rect 1490 1128 1546 1184
rect 2962 6160 3018 6216
rect 2962 4936 3018 4992
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 4526 10648 4582 10704
rect 3514 2352 3570 2408
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 7930 20304 7986 20360
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 6182 11736 6238 11792
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 6182 9152 6238 9208
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 4710 6296 4766 6352
rect 7838 13388 7894 13424
rect 7838 13368 7840 13388
rect 7840 13368 7892 13388
rect 7892 13368 7894 13388
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10138 19080 10194 19136
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 8942 17856 8998 17912
rect 8206 16496 8262 16552
rect 8942 16224 8998 16280
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 7286 7928 7342 7984
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 4710 5616 4766 5672
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5354 5752 5410 5808
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 8574 8472 8630 8528
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 12254 15000 12310 15056
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 13174 17176 13230 17232
rect 12990 14864 13046 14920
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11610 2896 11666 2952
rect 11886 9560 11942 9616
rect 13082 14320 13138 14376
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 13542 13368 13598 13424
rect 13450 9968 13506 10024
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 19154 21392 19210 21448
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 15842 16088 15898 16144
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15658 13368 15714 13424
rect 15382 13232 15438 13288
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 17590 17176 17646 17232
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 18694 17720 18750 17776
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 17682 16496 17738 16552
rect 17774 15952 17830 16008
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 16486 12008 16542 12064
rect 16026 10648 16082 10704
rect 13542 7792 13598 7848
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 16946 7928 17002 7984
rect 12622 6160 12678 6216
rect 17314 6160 17370 6216
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 17590 7928 17646 7984
rect 16118 3984 16174 4040
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15474 2896 15530 2952
rect 11794 2488 11850 2544
rect 10874 1808 10930 1864
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16394 2488 16450 2544
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 17866 10648 17922 10704
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 18602 11872 18658 11928
rect 25226 25608 25282 25664
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 25502 23432 25558 23488
rect 25502 22208 25558 22264
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 25134 20984 25190 21040
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24030 20304 24086 20360
rect 23018 19760 23074 19816
rect 22834 17720 22890 17776
rect 22466 17176 22522 17232
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 21730 15000 21786 15056
rect 22926 14864 22982 14920
rect 22190 13368 22246 13424
rect 18786 11600 18842 11656
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 23294 14320 23350 14376
rect 23110 13232 23166 13288
rect 23754 12824 23810 12880
rect 22006 11736 22062 11792
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19522 8880 19578 8936
rect 22006 9968 22062 10024
rect 19430 5616 19486 5672
rect 18878 3984 18934 4040
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 22834 10648 22890 10704
rect 22466 9968 22522 10024
rect 23754 11872 23810 11928
rect 22742 1808 22798 1864
rect 22006 1128 22062 1184
rect 23754 7792 23810 7848
rect 23938 16088 23994 16144
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24950 17448 25006 17504
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 16360 24822 16416
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24214 16088 24270 16144
rect 24030 15952 24086 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 26790 26832 26846 26888
rect 27618 25064 27674 25120
rect 26790 21392 26846 21448
rect 27618 19216 27674 19272
rect 24122 12008 24178 12064
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24766 11872 24822 11928
rect 24766 10512 24822 10568
rect 27618 14592 27674 14648
rect 25502 11600 25558 11656
rect 24674 9288 24730 9344
rect 24766 9152 24822 9208
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 27618 7520 27674 7576
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 27618 6296 27674 6352
rect 24858 6160 24914 6216
rect 24582 5752 24638 5808
rect 24766 5480 24822 5536
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 27618 3984 27674 4040
rect 25226 3168 25282 3224
rect 25134 2216 25190 2272
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
<< metal3 >>
rect 27520 27344 28000 27464
rect 0 27208 480 27328
rect 62 26890 122 27208
rect 1485 26890 1551 26893
rect 62 26888 1551 26890
rect 62 26832 1490 26888
rect 1546 26832 1551 26888
rect 62 26830 1551 26832
rect 1485 26827 1551 26830
rect 26785 26890 26851 26893
rect 27662 26890 27722 27344
rect 26785 26888 27722 26890
rect 26785 26832 26790 26888
rect 26846 26832 27722 26888
rect 26785 26830 27722 26832
rect 26785 26827 26851 26830
rect 27520 26120 28000 26240
rect 0 25984 480 26104
rect 62 25530 122 25984
rect 25221 25666 25287 25669
rect 27662 25666 27722 26120
rect 25221 25664 27722 25666
rect 25221 25608 25226 25664
rect 25282 25608 27722 25664
rect 25221 25606 27722 25608
rect 25221 25603 25287 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 5257 25530 5323 25533
rect 62 25528 5323 25530
rect 62 25472 5262 25528
rect 5318 25472 5323 25528
rect 62 25470 5323 25472
rect 5257 25467 5323 25470
rect 27520 25120 28000 25152
rect 27520 25064 27618 25120
rect 27674 25064 28000 25120
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 27520 25032 28000 25064
rect 24277 24991 24597 24992
rect 0 24624 480 24744
rect 62 24442 122 24624
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 1853 24442 1919 24445
rect 62 24440 1919 24442
rect 62 24384 1858 24440
rect 1914 24384 1919 24440
rect 62 24382 1919 24384
rect 1853 24379 1919 24382
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 27520 23808 28000 23928
rect 0 23400 480 23520
rect 25497 23490 25563 23493
rect 27662 23490 27722 23808
rect 25497 23488 27722 23490
rect 25497 23432 25502 23488
rect 25558 23432 27722 23488
rect 25497 23430 27722 23432
rect 25497 23427 25563 23430
rect 10277 23424 10597 23425
rect 62 22946 122 23400
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 1025 22946 1091 22949
rect 62 22944 1091 22946
rect 62 22888 1030 22944
rect 1086 22888 1091 22944
rect 62 22886 1091 22888
rect 1025 22883 1091 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 27520 22720 28000 22840
rect 10277 22336 10597 22337
rect 0 22176 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 25497 22266 25563 22269
rect 27662 22266 27722 22720
rect 25497 22264 27722 22266
rect 25497 22208 25502 22264
rect 25558 22208 27722 22264
rect 25497 22206 27722 22208
rect 25497 22203 25563 22206
rect 62 21722 122 22176
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1577 21722 1643 21725
rect 62 21720 1643 21722
rect 62 21664 1582 21720
rect 1638 21664 1643 21720
rect 62 21662 1643 21664
rect 1577 21659 1643 21662
rect 27520 21496 28000 21616
rect 19149 21450 19215 21453
rect 26785 21450 26851 21453
rect 19149 21448 26851 21450
rect 19149 21392 19154 21448
rect 19210 21392 26790 21448
rect 26846 21392 26851 21448
rect 19149 21390 26851 21392
rect 19149 21387 19215 21390
rect 26785 21387 26851 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 25129 21042 25195 21045
rect 27662 21042 27722 21496
rect 25129 21040 27722 21042
rect 25129 20984 25134 21040
rect 25190 20984 27722 21040
rect 25129 20982 27722 20984
rect 25129 20979 25195 20982
rect 0 20816 480 20936
rect 62 20362 122 20816
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 1577 20362 1643 20365
rect 62 20360 1643 20362
rect 62 20304 1582 20360
rect 1638 20304 1643 20360
rect 62 20302 1643 20304
rect 1577 20299 1643 20302
rect 7925 20362 7991 20365
rect 24025 20362 24091 20365
rect 7925 20360 24091 20362
rect 7925 20304 7930 20360
rect 7986 20304 24030 20360
rect 24086 20304 24091 20360
rect 7925 20302 24091 20304
rect 7925 20299 7991 20302
rect 24025 20299 24091 20302
rect 27520 20272 28000 20392
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 23013 19818 23079 19821
rect 27662 19818 27722 20272
rect 23013 19816 27722 19818
rect 23013 19760 23018 19816
rect 23074 19760 27722 19816
rect 23013 19758 27722 19760
rect 23013 19755 23079 19758
rect 0 19592 480 19712
rect 5610 19616 5930 19617
rect 62 19274 122 19592
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 1853 19274 1919 19277
rect 62 19272 1919 19274
rect 62 19216 1858 19272
rect 1914 19216 1919 19272
rect 62 19214 1919 19216
rect 1853 19211 1919 19214
rect 27520 19272 28000 19304
rect 27520 19216 27618 19272
rect 27674 19216 28000 19272
rect 27520 19184 28000 19216
rect 1669 19138 1735 19141
rect 10133 19138 10199 19141
rect 1669 19136 10199 19138
rect 1669 19080 1674 19136
rect 1730 19080 10138 19136
rect 10194 19080 10199 19136
rect 1669 19078 10199 19080
rect 1669 19075 1735 19078
rect 10133 19075 10199 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 5610 18528 5930 18529
rect 0 18368 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 62 17914 122 18368
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 18080
rect 19610 17919 19930 17920
rect 8937 17914 9003 17917
rect 62 17912 9003 17914
rect 62 17856 8942 17912
rect 8998 17856 9003 17912
rect 62 17854 9003 17856
rect 8937 17851 9003 17854
rect 18689 17778 18755 17781
rect 19374 17778 19380 17780
rect 18689 17776 19380 17778
rect 18689 17720 18694 17776
rect 18750 17720 19380 17776
rect 18689 17718 19380 17720
rect 18689 17715 18755 17718
rect 19374 17716 19380 17718
rect 19444 17778 19450 17780
rect 22829 17778 22895 17781
rect 19444 17776 22895 17778
rect 19444 17720 22834 17776
rect 22890 17720 22895 17776
rect 19444 17718 22895 17720
rect 19444 17716 19450 17718
rect 22829 17715 22895 17718
rect 2773 17642 2839 17645
rect 62 17640 2839 17642
rect 62 17584 2778 17640
rect 2834 17584 2839 17640
rect 62 17582 2839 17584
rect 62 17128 122 17582
rect 2773 17579 2839 17582
rect 24945 17506 25011 17509
rect 27662 17506 27722 17960
rect 24945 17504 27722 17506
rect 24945 17448 24950 17504
rect 25006 17448 27722 17504
rect 24945 17446 27722 17448
rect 24945 17443 25011 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 13169 17234 13235 17237
rect 17585 17234 17651 17237
rect 22461 17234 22527 17237
rect 13169 17232 22527 17234
rect 13169 17176 13174 17232
rect 13230 17176 17590 17232
rect 17646 17176 22466 17232
rect 22522 17176 22527 17232
rect 13169 17174 22527 17176
rect 13169 17171 13235 17174
rect 17585 17171 17651 17174
rect 22461 17171 22527 17174
rect 0 17008 480 17128
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 27520 16872 28000 16992
rect 19610 16831 19930 16832
rect 8201 16554 8267 16557
rect 17677 16554 17743 16557
rect 8201 16552 17743 16554
rect 8201 16496 8206 16552
rect 8262 16496 17682 16552
rect 17738 16496 17743 16552
rect 8201 16494 17743 16496
rect 8201 16491 8267 16494
rect 17677 16491 17743 16494
rect 24761 16418 24827 16421
rect 27662 16418 27722 16872
rect 24761 16416 27722 16418
rect 24761 16360 24766 16416
rect 24822 16360 27722 16416
rect 24761 16358 27722 16360
rect 24761 16355 24827 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 8937 16282 9003 16285
rect 8937 16280 13830 16282
rect 8937 16224 8942 16280
rect 8998 16224 13830 16280
rect 8937 16222 13830 16224
rect 8937 16219 9003 16222
rect 13770 16146 13830 16222
rect 15837 16146 15903 16149
rect 23933 16146 23999 16149
rect 13770 16144 23999 16146
rect 13770 16088 15842 16144
rect 15898 16088 23938 16144
rect 23994 16088 23999 16144
rect 13770 16086 23999 16088
rect 15837 16083 15903 16086
rect 23933 16083 23999 16086
rect 24209 16146 24275 16149
rect 24209 16144 27722 16146
rect 24209 16088 24214 16144
rect 24270 16088 27722 16144
rect 24209 16086 27722 16088
rect 24209 16083 24275 16086
rect 17769 16010 17835 16013
rect 24025 16010 24091 16013
rect 17769 16008 24091 16010
rect 17769 15952 17774 16008
rect 17830 15952 24030 16008
rect 24086 15952 24091 16008
rect 17769 15950 24091 15952
rect 17769 15947 17835 15950
rect 24025 15947 24091 15950
rect 0 15872 480 15904
rect 0 15816 18 15872
rect 74 15816 480 15872
rect 0 15784 480 15816
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 27662 15768 27722 16086
rect 19610 15743 19930 15744
rect 27520 15648 28000 15768
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 3693 15058 3759 15061
rect 12249 15058 12315 15061
rect 21725 15058 21791 15061
rect 3693 15056 21791 15058
rect 3693 15000 3698 15056
rect 3754 15000 12254 15056
rect 12310 15000 21730 15056
rect 21786 15000 21791 15056
rect 3693 14998 21791 15000
rect 3693 14995 3759 14998
rect 12249 14995 12315 14998
rect 21725 14995 21791 14998
rect 12985 14922 13051 14925
rect 22921 14922 22987 14925
rect 12985 14920 22987 14922
rect 12985 14864 12990 14920
rect 13046 14864 22926 14920
rect 22982 14864 22987 14920
rect 12985 14862 22987 14864
rect 12985 14859 13051 14862
rect 22921 14859 22987 14862
rect 10277 14720 10597 14721
rect 0 14648 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 0 14592 110 14648
rect 166 14592 480 14648
rect 0 14560 480 14592
rect 27520 14648 28000 14680
rect 27520 14592 27618 14648
rect 27674 14592 28000 14648
rect 27520 14560 28000 14592
rect 13077 14378 13143 14381
rect 23289 14378 23355 14381
rect 13077 14376 23355 14378
rect 13077 14320 13082 14376
rect 13138 14320 23294 14376
rect 23350 14320 23355 14376
rect 13077 14318 23355 14320
rect 13077 14315 13143 14318
rect 23289 14315 23355 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 1117 13562 1183 13565
rect 62 13560 1183 13562
rect 62 13504 1122 13560
rect 1178 13504 1183 13560
rect 62 13502 1183 13504
rect 62 13320 122 13502
rect 1117 13499 1183 13502
rect 7833 13426 7899 13429
rect 13537 13426 13603 13429
rect 7833 13424 13603 13426
rect 7833 13368 7838 13424
rect 7894 13368 13542 13424
rect 13598 13368 13603 13424
rect 7833 13366 13603 13368
rect 7833 13363 7899 13366
rect 13537 13363 13603 13366
rect 15653 13426 15719 13429
rect 22185 13426 22251 13429
rect 15653 13424 22251 13426
rect 15653 13368 15658 13424
rect 15714 13368 22190 13424
rect 22246 13368 22251 13424
rect 15653 13366 22251 13368
rect 15653 13363 15719 13366
rect 22185 13363 22251 13366
rect 27520 13336 28000 13456
rect 0 13200 480 13320
rect 15377 13290 15443 13293
rect 23105 13290 23171 13293
rect 15377 13288 23171 13290
rect 15377 13232 15382 13288
rect 15438 13232 23110 13288
rect 23166 13232 23171 13288
rect 15377 13230 23171 13232
rect 15377 13227 15443 13230
rect 23105 13227 23171 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 23749 12882 23815 12885
rect 27662 12882 27722 13336
rect 23749 12880 27722 12882
rect 23749 12824 23754 12880
rect 23810 12824 27722 12880
rect 23749 12822 27722 12824
rect 23749 12819 23815 12822
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 27520 12112 28000 12232
rect 0 12064 480 12096
rect 0 12008 110 12064
rect 166 12008 480 12064
rect 0 11976 480 12008
rect 16481 12066 16547 12069
rect 24117 12066 24183 12069
rect 16481 12064 24183 12066
rect 16481 12008 16486 12064
rect 16542 12008 24122 12064
rect 24178 12008 24183 12064
rect 16481 12006 24183 12008
rect 16481 12003 16547 12006
rect 24117 12003 24183 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 18597 11930 18663 11933
rect 23749 11930 23815 11933
rect 18597 11928 23815 11930
rect 18597 11872 18602 11928
rect 18658 11872 23754 11928
rect 23810 11872 23815 11928
rect 18597 11870 23815 11872
rect 18597 11867 18663 11870
rect 23749 11867 23815 11870
rect 24761 11930 24827 11933
rect 27662 11930 27722 12112
rect 24761 11928 27722 11930
rect 24761 11872 24766 11928
rect 24822 11872 27722 11928
rect 24761 11870 27722 11872
rect 24761 11867 24827 11870
rect 6177 11794 6243 11797
rect 22001 11794 22067 11797
rect 6177 11792 22067 11794
rect 6177 11736 6182 11792
rect 6238 11736 22006 11792
rect 22062 11736 22067 11792
rect 6177 11734 22067 11736
rect 6177 11731 6243 11734
rect 22001 11731 22067 11734
rect 18781 11658 18847 11661
rect 25497 11658 25563 11661
rect 18781 11656 25563 11658
rect 18781 11600 18786 11656
rect 18842 11600 25502 11656
rect 25558 11600 25563 11656
rect 18781 11598 25563 11600
rect 18781 11595 18847 11598
rect 25497 11595 25563 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 27520 11024 28000 11144
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10616 480 10736
rect 4521 10706 4587 10709
rect 16021 10706 16087 10709
rect 4521 10704 16087 10706
rect 4521 10648 4526 10704
rect 4582 10648 16026 10704
rect 16082 10648 16087 10704
rect 4521 10646 16087 10648
rect 4521 10643 4587 10646
rect 16021 10643 16087 10646
rect 17861 10706 17927 10709
rect 22829 10706 22895 10709
rect 17861 10704 22895 10706
rect 17861 10648 17866 10704
rect 17922 10648 22834 10704
rect 22890 10648 22895 10704
rect 17861 10646 22895 10648
rect 17861 10643 17927 10646
rect 22829 10643 22895 10646
rect 62 10162 122 10616
rect 24761 10570 24827 10573
rect 27662 10570 27722 11024
rect 24761 10568 27722 10570
rect 24761 10512 24766 10568
rect 24822 10512 27722 10568
rect 24761 10510 27722 10512
rect 24761 10507 24827 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 1577 10162 1643 10165
rect 62 10160 1643 10162
rect 62 10104 1582 10160
rect 1638 10104 1643 10160
rect 62 10102 1643 10104
rect 1577 10099 1643 10102
rect 13445 10026 13511 10029
rect 22001 10026 22067 10029
rect 22461 10026 22527 10029
rect 13445 10024 22527 10026
rect 13445 9968 13450 10024
rect 13506 9968 22006 10024
rect 22062 9968 22466 10024
rect 22522 9968 22527 10024
rect 13445 9966 22527 9968
rect 13445 9963 13511 9966
rect 22001 9963 22067 9966
rect 22461 9963 22527 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9920
rect 24277 9759 24597 9760
rect 11881 9618 11947 9621
rect 11881 9616 23490 9618
rect 11881 9560 11886 9616
rect 11942 9560 23490 9616
rect 11881 9558 23490 9560
rect 11881 9555 11947 9558
rect 0 9484 480 9512
rect 0 9420 60 9484
rect 124 9420 480 9484
rect 0 9392 480 9420
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 54 9148 60 9212
rect 124 9210 130 9212
rect 6177 9210 6243 9213
rect 124 9208 6243 9210
rect 124 9152 6182 9208
rect 6238 9152 6243 9208
rect 124 9150 6243 9152
rect 23430 9210 23490 9558
rect 24669 9346 24735 9349
rect 27662 9346 27722 9800
rect 24669 9344 27722 9346
rect 24669 9288 24674 9344
rect 24730 9288 27722 9344
rect 24669 9286 27722 9288
rect 24669 9283 24735 9286
rect 24761 9210 24827 9213
rect 23430 9208 27722 9210
rect 23430 9152 24766 9208
rect 24822 9152 27722 9208
rect 23430 9150 27722 9152
rect 124 9148 130 9150
rect 6177 9147 6243 9150
rect 24761 9147 24827 9150
rect 19374 8876 19380 8940
rect 19444 8938 19450 8940
rect 19517 8938 19583 8941
rect 19444 8936 19583 8938
rect 19444 8880 19522 8936
rect 19578 8880 19583 8936
rect 19444 8878 19583 8880
rect 19444 8876 19450 8878
rect 19517 8875 19583 8878
rect 27662 8832 27722 9150
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8832
rect 24277 8671 24597 8672
rect 8569 8530 8635 8533
rect 62 8528 8635 8530
rect 62 8472 8574 8528
rect 8630 8472 8635 8528
rect 62 8470 8635 8472
rect 62 8288 122 8470
rect 8569 8467 8635 8470
rect 0 8168 480 8288
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 7281 7986 7347 7989
rect 16941 7986 17007 7989
rect 17585 7986 17651 7989
rect 7281 7984 17651 7986
rect 7281 7928 7286 7984
rect 7342 7928 16946 7984
rect 17002 7928 17590 7984
rect 17646 7928 17651 7984
rect 7281 7926 17651 7928
rect 7281 7923 7347 7926
rect 16941 7923 17007 7926
rect 17585 7923 17651 7926
rect 13537 7850 13603 7853
rect 23749 7850 23815 7853
rect 13537 7848 23815 7850
rect 13537 7792 13542 7848
rect 13598 7792 23754 7848
rect 23810 7792 23815 7848
rect 13537 7790 23815 7792
rect 13537 7787 13603 7790
rect 23749 7787 23815 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 27520 7576 28000 7608
rect 27520 7520 27618 7576
rect 27674 7520 28000 7576
rect 27520 7488 28000 7520
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 0 6808 480 6928
rect 62 6354 122 6808
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 4705 6354 4771 6357
rect 62 6352 4771 6354
rect 62 6296 4710 6352
rect 4766 6296 4771 6352
rect 62 6294 4771 6296
rect 4705 6291 4771 6294
rect 27520 6352 28000 6384
rect 27520 6296 27618 6352
rect 27674 6296 28000 6352
rect 27520 6264 28000 6296
rect 2957 6218 3023 6221
rect 12617 6218 12683 6221
rect 2957 6216 12683 6218
rect 2957 6160 2962 6216
rect 3018 6160 12622 6216
rect 12678 6160 12683 6216
rect 2957 6158 12683 6160
rect 2957 6155 3023 6158
rect 12617 6155 12683 6158
rect 17309 6218 17375 6221
rect 24853 6218 24919 6221
rect 17309 6216 24919 6218
rect 17309 6160 17314 6216
rect 17370 6160 24858 6216
rect 24914 6160 24919 6216
rect 17309 6158 24919 6160
rect 17309 6155 17375 6158
rect 24853 6155 24919 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 5349 5810 5415 5813
rect 24577 5810 24643 5813
rect 5349 5808 24643 5810
rect 5349 5752 5354 5808
rect 5410 5752 24582 5808
rect 24638 5752 24643 5808
rect 5349 5750 24643 5752
rect 5349 5747 5415 5750
rect 24577 5747 24643 5750
rect 0 5584 480 5704
rect 4705 5674 4771 5677
rect 19425 5674 19491 5677
rect 4705 5672 19491 5674
rect 4705 5616 4710 5672
rect 4766 5616 19430 5672
rect 19486 5616 19491 5672
rect 4705 5614 19491 5616
rect 4705 5611 4771 5614
rect 19425 5611 19491 5614
rect 62 5130 122 5584
rect 24761 5538 24827 5541
rect 27654 5538 27660 5540
rect 24761 5536 27660 5538
rect 24761 5480 24766 5536
rect 24822 5480 27660 5536
rect 24761 5478 27660 5480
rect 24761 5475 24827 5478
rect 27654 5476 27660 5478
rect 27724 5476 27730 5540
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 27520 5268 28000 5296
rect 27520 5204 27660 5268
rect 27724 5204 28000 5268
rect 27520 5176 28000 5204
rect 1577 5130 1643 5133
rect 62 5128 1643 5130
rect 62 5072 1582 5128
rect 1638 5072 1643 5128
rect 62 5070 1643 5072
rect 1577 5067 1643 5070
rect 2957 4994 3023 4997
rect 62 4992 3023 4994
rect 62 4936 2962 4992
rect 3018 4936 3023 4992
rect 62 4934 3023 4936
rect 62 4480 122 4934
rect 2957 4931 3023 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 0 4360 480 4480
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 1669 4042 1735 4045
rect 16113 4042 16179 4045
rect 18873 4042 18939 4045
rect 1669 4040 18939 4042
rect 1669 3984 1674 4040
rect 1730 3984 16118 4040
rect 16174 3984 18878 4040
rect 18934 3984 18939 4040
rect 1669 3982 18939 3984
rect 1669 3979 1735 3982
rect 16113 3979 16179 3982
rect 18873 3979 18939 3982
rect 27520 4040 28000 4072
rect 27520 3984 27618 4040
rect 27674 3984 28000 4040
rect 27520 3952 28000 3984
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 25221 3226 25287 3229
rect 25221 3224 27722 3226
rect 25221 3168 25226 3224
rect 25282 3168 27722 3224
rect 25221 3166 27722 3168
rect 25221 3163 25287 3166
rect 0 3092 480 3120
rect 0 3028 60 3092
rect 124 3028 480 3092
rect 0 3000 480 3028
rect 27662 2984 27722 3166
rect 11605 2954 11671 2957
rect 15469 2954 15535 2957
rect 9630 2952 15535 2954
rect 9630 2896 11610 2952
rect 11666 2896 15474 2952
rect 15530 2896 15535 2952
rect 9630 2894 15535 2896
rect 54 2756 60 2820
rect 124 2818 130 2820
rect 9630 2818 9690 2894
rect 11605 2891 11671 2894
rect 15469 2891 15535 2894
rect 27520 2864 28000 2984
rect 124 2758 9690 2818
rect 124 2756 130 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 11789 2546 11855 2549
rect 16389 2546 16455 2549
rect 11789 2544 16455 2546
rect 11789 2488 11794 2544
rect 11850 2488 16394 2544
rect 16450 2488 16455 2544
rect 11789 2486 16455 2488
rect 11789 2483 11855 2486
rect 16389 2483 16455 2486
rect 3509 2410 3575 2413
rect 62 2408 3575 2410
rect 62 2352 3514 2408
rect 3570 2352 3575 2408
rect 62 2350 3575 2352
rect 62 1896 122 2350
rect 3509 2347 3575 2350
rect 25129 2274 25195 2277
rect 25129 2272 27722 2274
rect 25129 2216 25134 2272
rect 25190 2216 27722 2272
rect 25129 2214 27722 2216
rect 25129 2211 25195 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 0 1776 480 1896
rect 10869 1866 10935 1869
rect 22737 1866 22803 1869
rect 10869 1864 22803 1866
rect 10869 1808 10874 1864
rect 10930 1808 22742 1864
rect 22798 1808 22803 1864
rect 10869 1806 22803 1808
rect 10869 1803 10935 1806
rect 22737 1803 22803 1806
rect 27662 1760 27722 2214
rect 27520 1640 28000 1760
rect 1485 1186 1551 1189
rect 62 1184 1551 1186
rect 62 1128 1490 1184
rect 1546 1128 1551 1184
rect 62 1126 1551 1128
rect 62 672 122 1126
rect 1485 1123 1551 1126
rect 22001 1186 22067 1189
rect 22001 1184 27722 1186
rect 22001 1128 22006 1184
rect 22062 1128 27722 1184
rect 22001 1126 27722 1128
rect 22001 1123 22067 1126
rect 27662 672 27722 1126
rect 0 552 480 672
rect 27520 552 28000 672
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 19380 17716 19444 17780
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 60 9420 124 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 60 9148 124 9212
rect 19380 8876 19444 8940
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 27660 5476 27724 5540
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 27660 5204 27724 5268
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 60 3028 124 3092
rect 60 2756 124 2820
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 59 9484 125 9485
rect 59 9420 60 9484
rect 124 9420 125 9484
rect 59 9419 125 9420
rect 62 9213 122 9419
rect 59 9212 125 9213
rect 59 9148 60 9212
rect 124 9148 125 9212
rect 59 9147 125 9148
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 59 3092 125 3093
rect 59 3028 60 3092
rect 124 3028 125 3092
rect 59 3027 125 3028
rect 62 2821 122 3027
rect 59 2820 125 2821
rect 59 2756 60 2820
rect 124 2756 125 2820
rect 59 2755 125 2756
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19379 17780 19445 17781
rect 19379 17716 19380 17780
rect 19444 17716 19445 17780
rect 19379 17715 19445 17716
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 19382 8941 19442 17715
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19379 8940 19445 8941
rect 19379 8876 19380 8940
rect 19444 8876 19445 8940
rect 19379 8875 19445 8876
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 27659 5540 27725 5541
rect 27659 5476 27660 5540
rect 27724 5476 27725 5540
rect 27659 5475 27725 5476
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 27662 5269 27722 5475
rect 27659 5268 27725 5269
rect 27659 5204 27660 5268
rect 27724 5204 27725 5268
rect 27659 5203 27725 5204
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_40 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_44 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_48
timestamp 1586364061
transform 1 0 5520 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_60
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_75 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_81
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_103
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _171_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_111
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _170_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_153
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_164
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_184
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_236
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_4  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_262
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_274
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _176_
timestamp 1586364061
transform 1 0 23828 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_251
timestamp 1586364061
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_255
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_267
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_275
timestamp 1586364061
transform 1 0 26404 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _173_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_42
timestamp 1586364061
transform 1 0 4968 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_47
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_35
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_49
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use scs8hd_buf_2  _175_
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_259
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_263
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_275
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_22
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_conb_1  _158_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_8  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_37
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_54
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_78
timestamp 1586364061
transform 1 0 8280 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_89
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_90
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_102
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_109
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_121
timestamp 1586364061
transform 1 0 12236 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 590 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_206
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_222
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_242
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_253
timestamp 1586364061
transform 1 0 24380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_270
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_6  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_8  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_6  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_103
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_111
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _174_
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 774 592
use scs8hd_decap_6  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 590 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 406 592
use scs8hd_conb_1  _155_
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_58
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_67
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_84
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_169
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_173
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_177
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_200
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_212
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_224
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_13
timestamp 1586364061
transform 1 0 2300 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__C
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_8  _077_
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_55
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_96
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_100
timestamp 1586364061
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_116
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 1142 592
use scs8hd_conb_1  _153_
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_159
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_176
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_180
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _169_
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_259
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_or3_4  _084_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__138__D
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_20
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_24
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_30
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_45
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_49
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 590 592
use scs8hd_decap_4  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_100
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_111
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_nor4_4  _136_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__136__D
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_145
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_164
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_201
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_249
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_inv_8  _060_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _138_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__D
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__148__C
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_77
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 130 592
use scs8hd_nor4_4  _152_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__C
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_114
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _135_
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_219
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_231
timestamp 1586364061
transform 1 0 22356 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_243
timestamp 1586364061
transform 1 0 23460 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_270
timestamp 1586364061
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_8  _062_
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _064_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_12
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_24
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_20
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_24
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_nor4_4  _137_
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 1602 592
use scs8hd_nor4_4  _148_
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__148__D
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_45
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_50
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_38
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _147_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__D
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_54
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_58
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_82
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__D
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__C
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 866 592
use scs8hd_nor4_4  _151_
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_115
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__C
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_124
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use scs8hd_conb_1  _157_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_130
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_126
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__D
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__D
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_134
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _144_
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 1602 592
use scs8hd_inv_8  _071_
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_160
timestamp 1586364061
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_165
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_173
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_194
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _074_
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_203
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_199
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_213
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_230
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_242
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_249
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_236
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _183_
timestamp 1586364061
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_263
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_275
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_or3_4  _097_
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_10
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _061_
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_45
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_nor4_4  _150_
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _161_
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_162
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_201
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_207
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_223
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_230
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_234
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_238
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_or3_4  _134_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_8
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_12
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _063_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _078_
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_54
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_75
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_4  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__C
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _149_
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_169
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_173
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_176
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_235
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_259
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_or3_4  _105_
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_9
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _181_
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__105__C
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_38
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _070_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__142__D
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_87
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _142_
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__C
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_nor4_4  _143_
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _160_
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _079_
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_17_211
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 590 592
use scs8hd_inv_8  _073_
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_228
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_239
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_243
timestamp 1586364061
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_buf_2  _180_
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_250
timestamp 1586364061
transform 1 0 24104 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_263
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_267
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _069_
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_8
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_25
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_nor4_4  _140_
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_73
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_77
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _179_
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__141__C
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_115
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _133_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_183
timestamp 1586364061
transform 1 0 17940 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_188
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_200
timestamp 1586364061
transform 1 0 19504 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_204
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_212
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _156_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_218
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_222
timestamp 1586364061
transform 1 0 21528 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_229
timestamp 1586364061
transform 1 0 22172 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23920 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_240
timestamp 1586364061
transform 1 0 23184 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_262
timestamp 1586364061
transform 1 0 25208 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_274
timestamp 1586364061
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__C
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 1050 592
use scs8hd_nor4_4  _139_
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 1602 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__D
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_45
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 314 592
use scs8hd_or3_4  _095_
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_58
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_70
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_82
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _072_
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_109
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__D
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use scs8hd_nor4_4  _141_
timestamp 1586364061
transform 1 0 12512 0 1 12512
box -38 -48 1602 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_141
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_126
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_143
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_145
timestamp 1586364061
transform 1 0 14444 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_169
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_163
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_176
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_6  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 590 592
use scs8hd_decap_3  FILLER_19_170
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_184
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_buf_2  _168_
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_196
timestamp 1586364061
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_194
timestamp 1586364061
transform 1 0 18952 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_190
timestamp 1586364061
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18124 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_200
timestamp 1586364061
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_212
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_208
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_211
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_227
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_231
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_6  FILLER_19_238
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_241
timestamp 1586364061
transform 1 0 23276 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_251
timestamp 1586364061
transform 1 0 24196 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_252
timestamp 1586364061
transform 1 0 24288 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_264
timestamp 1586364061
transform 1 0 25392 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_272
timestamp 1586364061
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _178_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_12
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 314 592
use scs8hd_nor4_4  _145_
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 1602 592
use scs8hd_or3_4  _098_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_or3_4  _120_
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_155
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_176
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_188
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_202
timestamp 1586364061
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_206
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_221
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_225
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_248
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_252
timestamp 1586364061
transform 1 0 24288 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_264
timestamp 1586364061
transform 1 0 25392 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use scs8hd_or3_4  _089_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_conb_1  _159_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__C
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_or3_4  _093_
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__C
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_42
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__C
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_60
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_74
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_143
timestamp 1586364061
transform 1 0 14260 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 17388 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_170
timestamp 1586364061
transform 1 0 16744 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_176
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_205
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_228
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_241
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_253
timestamp 1586364061
transform 1 0 24380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_265
timestamp 1586364061
transform 1 0 25484 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_273
timestamp 1586364061
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_nor4_4  _146_
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 1602 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__C
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_8
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_33
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 406 592
use scs8hd_inv_8  _057_
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _059_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_90
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_94
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_129
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_139
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_205
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_218
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_222
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 23276 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_235
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_239
timestamp 1586364061
transform 1 0 23092 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_243
timestamp 1586364061
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_248
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_252
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_or3_4  _087_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_8  _058_
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_50
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_54
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_73
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__C
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_123
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_or3_4  _106_
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_136
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_140
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_170
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 17756 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_196
timestamp 1586364061
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _165_
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_201
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_205
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_226
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_230
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 406 592
use scs8hd_or3_4  _085_
timestamp 1586364061
transform 1 0 22632 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_243
timestamp 1586364061
transform 1 0 23460 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_10
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_40
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_67
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_84
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _164_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_130
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_144
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_148
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_157
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_161
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_174
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18952 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_190
timestamp 1586364061
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_205
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_209
timestamp 1586364061
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_224
timestamp 1586364061
transform 1 0 21712 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_228
timestamp 1586364061
transform 1 0 22080 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _163_
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23920 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_235
timestamp 1586364061
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_239
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_250
timestamp 1586364061
transform 1 0 24104 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_262
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_274
timestamp 1586364061
transform 1 0 26312 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_6
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_10
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _076_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_46
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_38
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_58
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_87
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_112
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_120
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_116
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_or3_4  _113_
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_138
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_142
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_157
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_165
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_169
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_161
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_182
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_194
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_212
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_219
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_229
timestamp 1586364061
transform 1 0 22172 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_27_238
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_234
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_240
timestamp 1586364061
transform 1 0 23184 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24012 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_251
timestamp 1586364061
transform 1 0 24196 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_262
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_266
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_274
timestamp 1586364061
transform 1 0 26312 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_10
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_50
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_65
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_113
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_123
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_172
timestamp 1586364061
transform 1 0 16928 0 -1 17952
box -38 -48 590 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_187
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_191
timestamp 1586364061
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_204
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_208
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_228
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_241
timestamp 1586364061
transform 1 0 23276 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_247
timestamp 1586364061
transform 1 0 23828 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_252
timestamp 1586364061
transform 1 0 24288 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_conb_1  _154_
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_9
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_13
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_17
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_30
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_42
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_72
timestamp 1586364061
transform 1 0 7728 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_102
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_144
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_158
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_162
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_187
timestamp 1586364061
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_191
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_212
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20976 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_227
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_231
timestamp 1586364061
transform 1 0 22356 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_235
timestamp 1586364061
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_239
timestamp 1586364061
transform 1 0 23092 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_254
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_274
timestamp 1586364061
transform 1 0 26312 0 1 17952
box -38 -48 314 592
use scs8hd_inv_8  _075_
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_13
timestamp 1586364061
transform 1 0 2300 0 -1 19040
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_29
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_6  FILLER_30_49
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_72
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_86
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 590 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_99
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_111
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_30_138
timestamp 1586364061
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_158
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_168
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 17664 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_189
timestamp 1586364061
transform 1 0 18492 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_195
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_219
timestamp 1586364061
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_229
timestamp 1586364061
transform 1 0 22172 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22908 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_12  FILLER_30_246
timestamp 1586364061
transform 1 0 23736 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_258
timestamp 1586364061
transform 1 0 24840 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_270
timestamp 1586364061
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _177_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_18
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_42
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 7084 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_76
timestamp 1586364061
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_102
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_134
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_138
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_151
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_169
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_188
timestamp 1586364061
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_192
timestamp 1586364061
transform 1 0 18768 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_204
timestamp 1586364061
transform 1 0 19872 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_213
timestamp 1586364061
transform 1 0 20700 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_226
timestamp 1586364061
transform 1 0 21896 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_230
timestamp 1586364061
transform 1 0 22264 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_238
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_249
timestamp 1586364061
transform 1 0 24012 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_261
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_31_273
timestamp 1586364061
transform 1 0 26220 0 1 19040
box -38 -48 406 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_29
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_43
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_47
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_62
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_66
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_79
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_87
timestamp 1586364061
transform 1 0 9108 0 -1 20128
box -38 -48 406 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_99
timestamp 1586364061
transform 1 0 10212 0 -1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_109
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_113
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_128
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_132
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_165
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_169
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_32_182
timestamp 1586364061
transform 1 0 17848 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_201
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_205
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_209
timestamp 1586364061
transform 1 0 20332 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_212
timestamp 1586364061
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_228
timestamp 1586364061
transform 1 0 22080 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_250
timestamp 1586364061
transform 1 0 24104 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_262
timestamp 1586364061
transform 1 0 25208 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_conb_1  _167_
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_49
timestamp 1586364061
transform 1 0 5612 0 -1 21216
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_6  FILLER_34_75
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_72
timestamp 1586364061
transform 1 0 7728 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_96
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_90
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_101
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_104
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_111
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_134
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_128
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_132
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_149
timestamp 1586364061
transform 1 0 14812 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_145
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_157
timestamp 1586364061
transform 1 0 15548 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15732 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_34_165
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_161
timestamp 1586364061
transform 1 0 15916 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_164
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_177
timestamp 1586364061
transform 1 0 17388 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_170
timestamp 1586364061
transform 1 0 16744 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_183
timestamp 1586364061
transform 1 0 17940 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_193
timestamp 1586364061
transform 1 0 18860 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_189
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_188
timestamp 1586364061
transform 1 0 18400 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19044 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18676 0 1 20128
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_206
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_206
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_219
timestamp 1586364061
transform 1 0 21252 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_230
timestamp 1586364061
transform 1 0 22264 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_226
timestamp 1586364061
transform 1 0 21896 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_223
timestamp 1586364061
transform 1 0 21620 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_236
timestamp 1586364061
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_243
timestamp 1586364061
transform 1 0 23460 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_258
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_262
timestamp 1586364061
transform 1 0 25208 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_266
timestamp 1586364061
transform 1 0 25576 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_258
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_274
timestamp 1586364061
transform 1 0 26312 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_270
timestamp 1586364061
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_19
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_31
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_43
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_49
timestamp 1586364061
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_72
timestamp 1586364061
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_76
timestamp 1586364061
transform 1 0 8096 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_89
timestamp 1586364061
transform 1 0 9292 0 1 21216
box -38 -48 406 592
use scs8hd_buf_2  _172_
timestamp 1586364061
transform 1 0 10028 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_101
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_105
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_117
timestamp 1586364061
transform 1 0 11868 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_142
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 14444 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_154
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_193
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_197
timestamp 1586364061
transform 1 0 19228 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_204
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_216
timestamp 1586364061
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_229
timestamp 1586364061
transform 1 0 22172 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_233
timestamp 1586364061
transform 1 0 22540 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_35_241
timestamp 1586364061
transform 1 0 23276 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_249
timestamp 1586364061
transform 1 0 24012 0 1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_6
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_18
timestamp 1586364061
transform 1 0 2760 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_30
timestamp 1586364061
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_65
timestamp 1586364061
transform 1 0 7084 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_82
timestamp 1586364061
transform 1 0 8648 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_86
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_96
timestamp 1586364061
transform 1 0 9936 0 -1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_36_120
timestamp 1586364061
transform 1 0 12144 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 866 592
use scs8hd_fill_2  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_136
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 774 592
use scs8hd_conb_1  _166_
timestamp 1586364061
transform 1 0 15548 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_144
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_147
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_3  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_160
timestamp 1586364061
transform 1 0 15824 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 22304
box -38 -48 866 592
use scs8hd_fill_1  FILLER_36_168
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_189
timestamp 1586364061
transform 1 0 18492 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_201
timestamp 1586364061
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_213
timestamp 1586364061
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use scs8hd_conb_1  _162_
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_218
timestamp 1586364061
transform 1 0 21160 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_222
timestamp 1586364061
transform 1 0 21528 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_229
timestamp 1586364061
transform 1 0 22172 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_241
timestamp 1586364061
transform 1 0 23276 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_246
timestamp 1586364061
transform 1 0 23736 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_254
timestamp 1586364061
transform 1 0 24472 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_258
timestamp 1586364061
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_270
timestamp 1586364061
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_6
timestamp 1586364061
transform 1 0 1656 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_10
timestamp 1586364061
transform 1 0 2024 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_22
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_34
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_46
timestamp 1586364061
transform 1 0 5336 0 1 22304
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_58
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_79
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_85
timestamp 1586364061
transform 1 0 8924 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_89
timestamp 1586364061
transform 1 0 9292 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_101
timestamp 1586364061
transform 1 0 10396 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 774 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_131
timestamp 1586364061
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_144
timestamp 1586364061
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_148
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_166
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_178
timestamp 1586364061
transform 1 0 17480 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_182
timestamp 1586364061
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19964 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_204
timestamp 1586364061
transform 1 0 19872 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_212
timestamp 1586364061
transform 1 0 20608 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_224
timestamp 1586364061
transform 1 0 21712 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 774 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_262
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_266
timestamp 1586364061
transform 1 0 25576 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_274
timestamp 1586364061
transform 1 0 26312 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_76
timestamp 1586364061
transform 1 0 8096 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_88
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_137
timestamp 1586364061
transform 1 0 13708 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16192 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_162
timestamp 1586364061
transform 1 0 16008 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_167
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_179
timestamp 1586364061
transform 1 0 17572 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_191
timestamp 1586364061
transform 1 0 18676 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_203
timestamp 1586364061
transform 1 0 19780 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_211
timestamp 1586364061
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_258
timestamp 1586364061
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_270
timestamp 1586364061
transform 1 0 25944 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_45
timestamp 1586364061
transform 1 0 5244 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_49
timestamp 1586364061
transform 1 0 5612 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_49
timestamp 1586364061
transform 1 0 5612 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_61
timestamp 1586364061
transform 1 0 6716 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_73
timestamp 1586364061
transform 1 0 7820 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_85
timestamp 1586364061
transform 1 0 8924 0 -1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_91
timestamp 1586364061
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _182_
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 13340 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_131
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_138
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_137
timestamp 1586364061
transform 1 0 13708 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_154
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_149
timestamp 1586364061
transform 1 0 14812 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_178
timestamp 1586364061
transform 1 0 17480 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_182
timestamp 1586364061
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 21252 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_216
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 3422 0 3478 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 4802 0 4858 480 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 552 480 672 6 address[2]
port 2 nsew default input
rlabel metal2 s 754 27520 810 28000 6 address[3]
port 3 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 1776 480 1896 6 address[5]
port 5 nsew default input
rlabel metal2 s 3974 27520 4030 28000 6 address[6]
port 6 nsew default input
rlabel metal2 s 6182 0 6238 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal2 s 7286 27520 7342 28000 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 27520 552 28000 672 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 27520 1640 28000 1760 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 27520 2864 28000 2984 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 27520 3952 28000 4072 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 27520 5176 28000 5296 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 27520 6264 28000 6384 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal2 s 8942 27520 8998 28000 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal2 s 13174 0 13230 480 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 27520 7488 28000 7608 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal2 s 14646 0 14702 480 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal2 s 16026 0 16082 480 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal2 s 10598 27520 10654 28000 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal2 s 15474 27520 15530 28000 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 27520 12112 28000 12232 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 13200 480 13320 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal3 s 27520 14560 28000 14680 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal2 s 17130 27520 17186 28000 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal2 s 18786 27520 18842 28000 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal2 s 20166 0 20222 480 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal3 s 0 18368 480 18488 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal3 s 27520 15648 28000 15768 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal3 s 27520 16872 28000 16992 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal2 s 20442 27520 20498 28000 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal2 s 21638 0 21694 480 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal3 s 27520 19184 28000 19304 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal2 s 2042 0 2098 480 6 data_in
port 63 nsew default input
rlabel metal2 s 662 0 718 480 6 enable
port 64 nsew default input
rlabel metal3 s 27520 20272 28000 20392 6 left_bottom_grid_pin_12_
port 65 nsew default input
rlabel metal2 s 24398 0 24454 480 6 left_top_grid_pin_11_
port 66 nsew default input
rlabel metal3 s 27520 25032 28000 25152 6 left_top_grid_pin_13_
port 67 nsew default input
rlabel metal2 s 25778 0 25834 480 6 left_top_grid_pin_15_
port 68 nsew default input
rlabel metal3 s 27520 21496 28000 21616 6 left_top_grid_pin_1_
port 69 nsew default input
rlabel metal3 s 27520 22720 28000 22840 6 left_top_grid_pin_3_
port 70 nsew default input
rlabel metal3 s 27520 23808 28000 23928 6 left_top_grid_pin_5_
port 71 nsew default input
rlabel metal2 s 23754 27520 23810 28000 6 left_top_grid_pin_7_
port 72 nsew default input
rlabel metal2 s 23018 0 23074 480 6 left_top_grid_pin_9_
port 73 nsew default input
rlabel metal2 s 25410 27520 25466 28000 6 right_bottom_grid_pin_12_
port 74 nsew default input
rlabel metal3 s 27520 27344 28000 27464 6 right_top_grid_pin_11_
port 75 nsew default input
rlabel metal2 s 27158 0 27214 480 6 right_top_grid_pin_13_
port 76 nsew default input
rlabel metal3 s 0 27208 480 27328 6 right_top_grid_pin_15_
port 77 nsew default input
rlabel metal3 s 0 23400 480 23520 6 right_top_grid_pin_1_
port 78 nsew default input
rlabel metal3 s 27520 26120 28000 26240 6 right_top_grid_pin_3_
port 79 nsew default input
rlabel metal3 s 0 24624 480 24744 6 right_top_grid_pin_5_
port 80 nsew default input
rlabel metal2 s 27066 27520 27122 28000 6 right_top_grid_pin_7_
port 81 nsew default input
rlabel metal3 s 0 25984 480 26104 6 right_top_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
