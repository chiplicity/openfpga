magic
tech sky130A
magscale 1 2
timestamp 1605013381
<< locali >>
rect 10609 22015 10643 22321
rect 11621 2975 11655 3145
<< viali >>
rect 10609 22321 10643 22355
rect 10609 21981 10643 22015
rect 19257 20961 19291 20995
rect 21557 20961 21591 20995
rect 21741 20825 21775 20859
rect 19441 20757 19475 20791
rect 8677 20553 8711 20587
rect 10149 20553 10183 20587
rect 19349 20553 19383 20587
rect 21557 20553 21591 20587
rect 20637 20485 20671 20519
rect 23857 20485 23891 20519
rect 8493 20349 8527 20383
rect 9045 20349 9079 20383
rect 12541 20349 12575 20383
rect 13093 20349 13127 20383
rect 16313 20349 16347 20383
rect 16957 20349 16991 20383
rect 18061 20349 18095 20383
rect 19165 20349 19199 20383
rect 19717 20349 19751 20383
rect 20453 20349 20487 20383
rect 21097 20349 21131 20383
rect 21741 20349 21775 20383
rect 22293 20349 22327 20383
rect 23673 20349 23707 20383
rect 24225 20349 24259 20383
rect 20177 20281 20211 20315
rect 12725 20213 12759 20247
rect 16497 20213 16531 20247
rect 18245 20213 18279 20247
rect 18705 20213 18739 20247
rect 21925 20213 21959 20247
rect 18613 20009 18647 20043
rect 21097 20009 21131 20043
rect 17325 19873 17359 19907
rect 18429 19873 18463 19907
rect 19533 19873 19567 19907
rect 20913 19873 20947 19907
rect 17509 19737 17543 19771
rect 19717 19737 19751 19771
rect 17325 19465 17359 19499
rect 18521 19125 18555 19159
rect 19533 19125 19567 19159
rect 20913 19125 20947 19159
rect 11805 14501 11839 14535
rect 11897 14433 11931 14467
rect 12081 14365 12115 14399
rect 11437 14229 11471 14263
rect 11529 14025 11563 14059
rect 12173 14025 12207 14059
rect 13553 13889 13587 13923
rect 2513 13821 2547 13855
rect 13645 13821 13679 13855
rect 13912 13821 13946 13855
rect 11805 13753 11839 13787
rect 1685 13685 1719 13719
rect 3065 13685 3099 13719
rect 10241 13685 10275 13719
rect 15025 13685 15059 13719
rect 2421 13481 2455 13515
rect 12173 13481 12207 13515
rect 12633 13413 12667 13447
rect 2789 13345 2823 13379
rect 4629 13345 4663 13379
rect 5264 13345 5298 13379
rect 9956 13345 9990 13379
rect 12541 13345 12575 13379
rect 2329 13277 2363 13311
rect 2881 13277 2915 13311
rect 3065 13277 3099 13311
rect 4997 13277 5031 13311
rect 7757 13277 7791 13311
rect 9505 13277 9539 13311
rect 9689 13277 9723 13311
rect 12725 13277 12759 13311
rect 1685 13141 1719 13175
rect 6377 13141 6411 13175
rect 11069 13141 11103 13175
rect 13737 13141 13771 13175
rect 2973 12937 3007 12971
rect 4537 12937 4571 12971
rect 11805 12937 11839 12971
rect 12265 12937 12299 12971
rect 1409 12869 1443 12903
rect 9045 12869 9079 12903
rect 9781 12869 9815 12903
rect 11529 12869 11563 12903
rect 1869 12801 1903 12835
rect 2053 12801 2087 12835
rect 3433 12801 3467 12835
rect 3617 12801 3651 12835
rect 5181 12801 5215 12835
rect 7665 12801 7699 12835
rect 10609 12801 10643 12835
rect 10793 12801 10827 12835
rect 13001 12801 13035 12835
rect 14749 12801 14783 12835
rect 1777 12733 1811 12767
rect 2881 12733 2915 12767
rect 3341 12733 3375 12767
rect 4905 12733 4939 12767
rect 4997 12733 5031 12767
rect 12817 12733 12851 12767
rect 14933 12733 14967 12767
rect 15189 12733 15223 12767
rect 2513 12665 2547 12699
rect 4445 12665 4479 12699
rect 7910 12665 7944 12699
rect 4077 12597 4111 12631
rect 5641 12597 5675 12631
rect 7481 12597 7515 12631
rect 10149 12597 10183 12631
rect 10517 12597 10551 12631
rect 12449 12597 12483 12631
rect 12909 12597 12943 12631
rect 13461 12597 13495 12631
rect 16313 12597 16347 12631
rect 2421 12393 2455 12427
rect 3525 12393 3559 12427
rect 4537 12393 4571 12427
rect 4997 12393 5031 12427
rect 7205 12393 7239 12427
rect 9505 12393 9539 12427
rect 9689 12393 9723 12427
rect 10793 12393 10827 12427
rect 12173 12393 12207 12427
rect 12817 12393 12851 12427
rect 13093 12393 13127 12427
rect 13645 12393 13679 12427
rect 1685 12325 1719 12359
rect 6092 12325 6126 12359
rect 2329 12257 2363 12291
rect 2789 12257 2823 12291
rect 5825 12257 5859 12291
rect 10057 12257 10091 12291
rect 12081 12257 12115 12291
rect 13737 12257 13771 12291
rect 15025 12257 15059 12291
rect 16497 12257 16531 12291
rect 16753 12257 16787 12291
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 12357 12189 12391 12223
rect 13829 12189 13863 12223
rect 11713 12053 11747 12087
rect 13277 12053 13311 12087
rect 17877 12053 17911 12087
rect 18521 12053 18555 12087
rect 2605 11849 2639 11883
rect 2789 11849 2823 11883
rect 3801 11849 3835 11883
rect 4261 11849 4295 11883
rect 5917 11849 5951 11883
rect 9413 11849 9447 11883
rect 9597 11849 9631 11883
rect 11437 11849 11471 11883
rect 12449 11849 12483 11883
rect 16589 11849 16623 11883
rect 18245 11849 18279 11883
rect 6193 11781 6227 11815
rect 11805 11781 11839 11815
rect 2053 11713 2087 11747
rect 3433 11713 3467 11747
rect 8769 11713 8803 11747
rect 10149 11713 10183 11747
rect 12265 11713 12299 11747
rect 13001 11713 13035 11747
rect 1409 11645 1443 11679
rect 10057 11645 10091 11679
rect 12817 11645 12851 11679
rect 14197 11645 14231 11679
rect 16957 11645 16991 11679
rect 18429 11645 18463 11679
rect 18696 11645 18730 11679
rect 26433 11645 26467 11679
rect 26985 11645 27019 11679
rect 3157 11577 3191 11611
rect 9045 11577 9079 11611
rect 13553 11577 13587 11611
rect 1593 11509 1627 11543
rect 3249 11509 3283 11543
rect 9965 11509 9999 11543
rect 10701 11509 10735 11543
rect 12909 11509 12943 11543
rect 13829 11509 13863 11543
rect 19809 11509 19843 11543
rect 26617 11509 26651 11543
rect 2329 11305 2363 11339
rect 2421 11305 2455 11339
rect 3433 11305 3467 11339
rect 4077 11305 4111 11339
rect 8125 11305 8159 11339
rect 10241 11305 10275 11339
rect 11805 11305 11839 11339
rect 12541 11305 12575 11339
rect 12909 11305 12943 11339
rect 13369 11305 13403 11339
rect 7012 11237 7046 11271
rect 12173 11237 12207 11271
rect 2789 11169 2823 11203
rect 4445 11169 4479 11203
rect 6745 11169 6779 11203
rect 13277 11169 13311 11203
rect 17693 11169 17727 11203
rect 26525 11169 26559 11203
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 13461 11101 13495 11135
rect 17785 11101 17819 11135
rect 17969 11101 18003 11135
rect 9965 11033 9999 11067
rect 16497 11033 16531 11067
rect 26709 11033 26743 11067
rect 17325 10965 17359 10999
rect 18429 10965 18463 10999
rect 1593 10761 1627 10795
rect 2053 10761 2087 10795
rect 2421 10761 2455 10795
rect 3249 10761 3283 10795
rect 7389 10761 7423 10795
rect 13001 10761 13035 10795
rect 13553 10761 13587 10795
rect 26525 10761 26559 10795
rect 18061 10693 18095 10727
rect 2789 10625 2823 10659
rect 3893 10625 3927 10659
rect 9965 10625 9999 10659
rect 10609 10625 10643 10659
rect 13093 10625 13127 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 17785 10625 17819 10659
rect 18613 10625 18647 10659
rect 19073 10625 19107 10659
rect 1409 10557 1443 10591
rect 9229 10557 9263 10591
rect 15945 10557 15979 10591
rect 16773 10557 16807 10591
rect 18521 10557 18555 10591
rect 3157 10489 3191 10523
rect 9597 10489 9631 10523
rect 10517 10489 10551 10523
rect 16313 10489 16347 10523
rect 3617 10421 3651 10455
rect 3709 10421 3743 10455
rect 4353 10421 4387 10455
rect 4629 10421 4663 10455
rect 5089 10421 5123 10455
rect 7113 10421 7147 10455
rect 10057 10421 10091 10455
rect 10425 10421 10459 10455
rect 16405 10421 16439 10455
rect 17417 10421 17451 10455
rect 18429 10421 18463 10455
rect 1593 10217 1627 10251
rect 2789 10217 2823 10251
rect 3341 10217 3375 10251
rect 4445 10217 4479 10251
rect 6929 10217 6963 10251
rect 7941 10217 7975 10251
rect 11069 10217 11103 10251
rect 13001 10217 13035 10251
rect 14749 10217 14783 10251
rect 16589 10217 16623 10251
rect 17693 10217 17727 10251
rect 18705 10217 18739 10251
rect 26709 10217 26743 10251
rect 9934 10149 9968 10183
rect 1409 10081 1443 10115
rect 4537 10081 4571 10115
rect 8125 10081 8159 10115
rect 14933 10081 14967 10115
rect 16497 10081 16531 10115
rect 18061 10081 18095 10115
rect 26525 10081 26559 10115
rect 4721 10013 4755 10047
rect 9689 10013 9723 10047
rect 12173 10013 12207 10047
rect 16773 10013 16807 10047
rect 17325 10013 17359 10047
rect 18153 10013 18187 10047
rect 18337 10013 18371 10047
rect 2513 9945 2547 9979
rect 4077 9945 4111 9979
rect 16129 9877 16163 9911
rect 2421 9673 2455 9707
rect 4537 9673 4571 9707
rect 4905 9673 4939 9707
rect 8217 9673 8251 9707
rect 10793 9673 10827 9707
rect 1593 9605 1627 9639
rect 2053 9605 2087 9639
rect 4169 9605 4203 9639
rect 9321 9605 9355 9639
rect 10609 9605 10643 9639
rect 17049 9605 17083 9639
rect 19441 9605 19475 9639
rect 6837 9537 6871 9571
rect 11253 9537 11287 9571
rect 11437 9537 11471 9571
rect 14013 9537 14047 9571
rect 18521 9537 18555 9571
rect 18705 9537 18739 9571
rect 19073 9537 19107 9571
rect 1409 9469 1443 9503
rect 11161 9469 11195 9503
rect 13921 9469 13955 9503
rect 14280 9469 14314 9503
rect 16589 9469 16623 9503
rect 17693 9469 17727 9503
rect 18429 9469 18463 9503
rect 19809 9469 19843 9503
rect 26525 9469 26559 9503
rect 6653 9401 6687 9435
rect 7104 9401 7138 9435
rect 9781 9401 9815 9435
rect 10333 9401 10367 9435
rect 8769 9333 8803 9367
rect 15393 9333 15427 9367
rect 16221 9333 16255 9367
rect 17325 9333 17359 9367
rect 18061 9333 18095 9367
rect 1593 9129 1627 9163
rect 3157 9129 3191 9163
rect 10885 9129 10919 9163
rect 11161 9129 11195 9163
rect 11529 9129 11563 9163
rect 14013 9129 14047 9163
rect 15669 9129 15703 9163
rect 16129 9129 16163 9163
rect 17325 9129 17359 9163
rect 17785 9129 17819 9163
rect 18889 9129 18923 9163
rect 19257 9129 19291 9163
rect 26709 9129 26743 9163
rect 16221 9061 16255 9095
rect 16865 9061 16899 9095
rect 19349 9061 19383 9095
rect 1409 8993 1443 9027
rect 2513 8993 2547 9027
rect 5733 8993 5767 9027
rect 5989 8993 6023 9027
rect 11621 8993 11655 9027
rect 17693 8993 17727 9027
rect 18613 8993 18647 9027
rect 26525 8993 26559 9027
rect 11805 8925 11839 8959
rect 16313 8925 16347 8959
rect 17969 8925 18003 8959
rect 19441 8925 19475 8959
rect 15761 8857 15795 8891
rect 2697 8789 2731 8823
rect 7113 8789 7147 8823
rect 8953 8789 8987 8823
rect 14749 8789 14783 8823
rect 1593 8585 1627 8619
rect 2513 8585 2547 8619
rect 5825 8585 5859 8619
rect 7205 8585 7239 8619
rect 11621 8585 11655 8619
rect 17417 8585 17451 8619
rect 17785 8585 17819 8619
rect 18521 8585 18555 8619
rect 19533 8585 19567 8619
rect 26617 8585 26651 8619
rect 6193 8517 6227 8551
rect 8861 8517 8895 8551
rect 11253 8517 11287 8551
rect 13829 8517 13863 8551
rect 17049 8517 17083 8551
rect 27353 8517 27387 8551
rect 27721 8517 27755 8551
rect 2053 8449 2087 8483
rect 3249 8449 3283 8483
rect 3433 8449 3467 8483
rect 7941 8449 7975 8483
rect 9505 8449 9539 8483
rect 14749 8449 14783 8483
rect 18337 8449 18371 8483
rect 18981 8449 19015 8483
rect 19165 8449 19199 8483
rect 1409 8381 1443 8415
rect 7665 8381 7699 8415
rect 8769 8381 8803 8415
rect 9229 8381 9263 8415
rect 14013 8381 14047 8415
rect 14841 8381 14875 8415
rect 15108 8381 15142 8415
rect 26433 8381 26467 8415
rect 26985 8381 27019 8415
rect 27537 8381 27571 8415
rect 28089 8381 28123 8415
rect 3157 8313 3191 8347
rect 3893 8313 3927 8347
rect 4353 8313 4387 8347
rect 6653 8313 6687 8347
rect 7757 8313 7791 8347
rect 8401 8313 8435 8347
rect 9321 8313 9355 8347
rect 14289 8313 14323 8347
rect 19901 8313 19935 8347
rect 2789 8245 2823 8279
rect 7297 8245 7331 8279
rect 11989 8245 12023 8279
rect 16221 8245 16255 8279
rect 18889 8245 18923 8279
rect 2329 8041 2363 8075
rect 2881 8041 2915 8075
rect 7021 8041 7055 8075
rect 7665 8041 7699 8075
rect 14105 8041 14139 8075
rect 14841 8041 14875 8075
rect 16221 8041 16255 8075
rect 18613 8041 18647 8075
rect 18981 8041 19015 8075
rect 19441 8041 19475 8075
rect 26709 8041 26743 8075
rect 6929 7973 6963 8007
rect 2789 7905 2823 7939
rect 9045 7905 9079 7939
rect 11345 7905 11379 7939
rect 14013 7905 14047 7939
rect 15853 7905 15887 7939
rect 16753 7905 16787 7939
rect 26525 7905 26559 7939
rect 1685 7837 1719 7871
rect 3065 7837 3099 7871
rect 7113 7837 7147 7871
rect 14197 7837 14231 7871
rect 16497 7837 16531 7871
rect 12633 7769 12667 7803
rect 2421 7701 2455 7735
rect 3525 7701 3559 7735
rect 4353 7701 4387 7735
rect 6561 7701 6595 7735
rect 8861 7701 8895 7735
rect 10793 7701 10827 7735
rect 13461 7701 13495 7735
rect 13645 7701 13679 7735
rect 17877 7701 17911 7735
rect 2329 7497 2363 7531
rect 5641 7497 5675 7531
rect 6653 7497 6687 7531
rect 7113 7497 7147 7531
rect 7481 7497 7515 7531
rect 8309 7497 8343 7531
rect 10517 7497 10551 7531
rect 14289 7497 14323 7531
rect 16589 7497 16623 7531
rect 27353 7497 27387 7531
rect 9137 7429 9171 7463
rect 16865 7429 16899 7463
rect 1961 7361 1995 7395
rect 3065 7361 3099 7395
rect 9045 7361 9079 7395
rect 9689 7361 9723 7395
rect 11161 7361 11195 7395
rect 11345 7361 11379 7395
rect 12817 7361 12851 7395
rect 13737 7361 13771 7395
rect 13921 7361 13955 7395
rect 2789 7293 2823 7327
rect 4261 7293 4295 7327
rect 26433 7293 26467 7327
rect 26985 7293 27019 7327
rect 2881 7225 2915 7259
rect 3525 7225 3559 7259
rect 4169 7225 4203 7259
rect 4528 7225 4562 7259
rect 8677 7225 8711 7259
rect 9505 7225 9539 7259
rect 11713 7225 11747 7259
rect 13093 7225 13127 7259
rect 13645 7225 13679 7259
rect 14841 7225 14875 7259
rect 2421 7157 2455 7191
rect 9597 7157 9631 7191
rect 10701 7157 10735 7191
rect 11069 7157 11103 7191
rect 13277 7157 13311 7191
rect 14749 7157 14783 7191
rect 26617 7157 26651 7191
rect 2053 6953 2087 6987
rect 13277 6953 13311 6987
rect 14013 6953 14047 6987
rect 2329 6885 2363 6919
rect 5978 6885 6012 6919
rect 1409 6817 1443 6851
rect 2513 6817 2547 6851
rect 4077 6817 4111 6851
rect 8401 6817 8435 6851
rect 10057 6817 10091 6851
rect 11417 6817 11451 6851
rect 13369 6817 13403 6851
rect 18144 6817 18178 6851
rect 26525 6817 26559 6851
rect 5733 6749 5767 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 10701 6749 10735 6783
rect 11161 6749 11195 6783
rect 13461 6749 13495 6783
rect 17877 6749 17911 6783
rect 2697 6681 2731 6715
rect 4261 6681 4295 6715
rect 9689 6681 9723 6715
rect 12541 6681 12575 6715
rect 26709 6681 26743 6715
rect 1593 6613 1627 6647
rect 3065 6613 3099 6647
rect 7113 6613 7147 6647
rect 8217 6613 8251 6647
rect 9229 6613 9263 6647
rect 12909 6613 12943 6647
rect 16037 6613 16071 6647
rect 19257 6613 19291 6647
rect 1685 6409 1719 6443
rect 3065 6409 3099 6443
rect 4169 6409 4203 6443
rect 5733 6409 5767 6443
rect 9873 6409 9907 6443
rect 12265 6409 12299 6443
rect 15761 6409 15795 6443
rect 18613 6409 18647 6443
rect 3801 6341 3835 6375
rect 4629 6341 4663 6375
rect 8769 6341 8803 6375
rect 2605 6273 2639 6307
rect 9781 6273 9815 6307
rect 10425 6273 10459 6307
rect 10885 6273 10919 6307
rect 11253 6273 11287 6307
rect 13369 6273 13403 6307
rect 16497 6273 16531 6307
rect 2421 6205 2455 6239
rect 2513 6205 2547 6239
rect 3617 6205 3651 6239
rect 7205 6205 7239 6239
rect 7389 6205 7423 6239
rect 10333 6205 10367 6239
rect 13461 6205 13495 6239
rect 13728 6205 13762 6239
rect 16313 6205 16347 6239
rect 26525 6205 26559 6239
rect 3433 6137 3467 6171
rect 7634 6137 7668 6171
rect 13001 6137 13035 6171
rect 15485 6137 15519 6171
rect 16405 6137 16439 6171
rect 2053 6069 2087 6103
rect 6193 6069 6227 6103
rect 9321 6069 9355 6103
rect 10241 6069 10275 6103
rect 11621 6069 11655 6103
rect 14841 6069 14875 6103
rect 15945 6069 15979 6103
rect 18245 6069 18279 6103
rect 2145 5865 2179 5899
rect 2421 5865 2455 5899
rect 2789 5865 2823 5899
rect 4077 5865 4111 5899
rect 8309 5865 8343 5899
rect 10609 5865 10643 5899
rect 13001 5865 13035 5899
rect 13553 5865 13587 5899
rect 14289 5865 14323 5899
rect 15669 5865 15703 5899
rect 16221 5865 16255 5899
rect 17325 5865 17359 5899
rect 17693 5865 17727 5899
rect 26709 5865 26743 5899
rect 9965 5797 9999 5831
rect 4445 5729 4479 5763
rect 14473 5729 14507 5763
rect 16129 5729 16163 5763
rect 26525 5729 26559 5763
rect 2881 5661 2915 5695
rect 3065 5661 3099 5695
rect 3893 5661 3927 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 16313 5661 16347 5695
rect 17785 5661 17819 5695
rect 17877 5661 17911 5695
rect 18337 5661 18371 5695
rect 7389 5525 7423 5559
rect 10241 5525 10275 5559
rect 15761 5525 15795 5559
rect 2053 5321 2087 5355
rect 3893 5321 3927 5355
rect 4997 5321 5031 5355
rect 13277 5321 13311 5355
rect 15577 5321 15611 5355
rect 16405 5321 16439 5355
rect 18061 5321 18095 5355
rect 26249 5321 26283 5355
rect 26617 5321 26651 5355
rect 26985 5253 27019 5287
rect 4537 5185 4571 5219
rect 15945 5185 15979 5219
rect 16957 5185 16991 5219
rect 18613 5185 18647 5219
rect 1409 5117 1443 5151
rect 2421 5117 2455 5151
rect 2513 5117 2547 5151
rect 3433 5117 3467 5151
rect 4261 5117 4295 5151
rect 13369 5117 13403 5151
rect 13625 5117 13659 5151
rect 16773 5117 16807 5151
rect 18429 5117 18463 5151
rect 26433 5117 26467 5151
rect 5365 5049 5399 5083
rect 18521 5049 18555 5083
rect 1593 4981 1627 5015
rect 2697 4981 2731 5015
rect 3801 4981 3835 5015
rect 4353 4981 4387 5015
rect 5733 4981 5767 5015
rect 14749 4981 14783 5015
rect 16313 4981 16347 5015
rect 16865 4981 16899 5015
rect 17509 4981 17543 5015
rect 17785 4981 17819 5015
rect 2053 4777 2087 4811
rect 4077 4777 4111 4811
rect 7297 4777 7331 4811
rect 12725 4777 12759 4811
rect 13369 4777 13403 4811
rect 14381 4777 14415 4811
rect 15761 4777 15795 4811
rect 16497 4777 16531 4811
rect 17693 4777 17727 4811
rect 18153 4777 18187 4811
rect 26709 4777 26743 4811
rect 2421 4709 2455 4743
rect 3065 4709 3099 4743
rect 15669 4709 15703 4743
rect 17417 4709 17451 4743
rect 1409 4641 1443 4675
rect 2513 4641 2547 4675
rect 3893 4641 3927 4675
rect 4445 4641 4479 4675
rect 6173 4641 6207 4675
rect 12817 4641 12851 4675
rect 26525 4641 26559 4675
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 5917 4573 5951 4607
rect 12909 4573 12943 4607
rect 15853 4573 15887 4607
rect 1593 4437 1627 4471
rect 2697 4437 2731 4471
rect 12357 4437 12391 4471
rect 15301 4437 15335 4471
rect 3985 4233 4019 4267
rect 5457 4233 5491 4267
rect 12265 4233 12299 4267
rect 13093 4233 13127 4267
rect 15393 4233 15427 4267
rect 16129 4233 16163 4267
rect 27353 4233 27387 4267
rect 1961 4097 1995 4131
rect 3433 4097 3467 4131
rect 4629 4097 4663 4131
rect 4997 4097 5031 4131
rect 5917 4097 5951 4131
rect 15025 4097 15059 4131
rect 1409 4029 1443 4063
rect 2421 4029 2455 4063
rect 2513 4029 2547 4063
rect 4353 4029 4387 4063
rect 7665 4029 7699 4063
rect 8493 4029 8527 4063
rect 15853 4029 15887 4063
rect 26433 4029 26467 4063
rect 26985 4029 27019 4063
rect 3157 3961 3191 3995
rect 7941 3961 7975 3995
rect 1593 3893 1627 3927
rect 2697 3893 2731 3927
rect 3893 3893 3927 3927
rect 4445 3893 4479 3927
rect 6285 3893 6319 3927
rect 12725 3893 12759 3927
rect 26617 3893 26651 3927
rect 1961 3689 1995 3723
rect 3157 3689 3191 3723
rect 3893 3689 3927 3723
rect 4077 3689 4111 3723
rect 4445 3689 4479 3723
rect 14933 3689 14967 3723
rect 26709 3689 26743 3723
rect 8677 3621 8711 3655
rect 1409 3553 1443 3587
rect 2513 3553 2547 3587
rect 4537 3553 4571 3587
rect 9781 3553 9815 3587
rect 11069 3553 11103 3587
rect 11325 3553 11359 3587
rect 15301 3553 15335 3587
rect 25329 3553 25363 3587
rect 26525 3553 26559 3587
rect 4629 3485 4663 3519
rect 1593 3349 1627 3383
rect 2697 3349 2731 3383
rect 5089 3349 5123 3383
rect 9965 3349 9999 3383
rect 12449 3349 12483 3383
rect 15485 3349 15519 3383
rect 25513 3349 25547 3383
rect 2237 3145 2271 3179
rect 2605 3145 2639 3179
rect 3617 3145 3651 3179
rect 4813 3145 4847 3179
rect 5273 3145 5307 3179
rect 6193 3145 6227 3179
rect 9965 3145 9999 3179
rect 10517 3145 10551 3179
rect 11621 3145 11655 3179
rect 11897 3145 11931 3179
rect 14473 3145 14507 3179
rect 25145 3145 25179 3179
rect 25881 3145 25915 3179
rect 26617 3145 26651 3179
rect 27353 3145 27387 3179
rect 3985 3077 4019 3111
rect 8585 3009 8619 3043
rect 12173 3009 12207 3043
rect 1409 2941 1443 2975
rect 2789 2941 2823 2975
rect 3065 2941 3099 2975
rect 4077 2941 4111 2975
rect 5365 2941 5399 2975
rect 11253 2941 11287 2975
rect 11621 2941 11655 2975
rect 12449 2941 12483 2975
rect 12716 2941 12750 2975
rect 14749 2941 14783 2975
rect 14933 2941 14967 2975
rect 18153 2941 18187 2975
rect 18705 2941 18739 2975
rect 25329 2941 25363 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 27537 2941 27571 2975
rect 28089 2941 28123 2975
rect 1685 2873 1719 2907
rect 4353 2873 4387 2907
rect 5641 2873 5675 2907
rect 8830 2873 8864 2907
rect 11069 2873 11103 2907
rect 15178 2873 15212 2907
rect 8401 2805 8435 2839
rect 11437 2805 11471 2839
rect 13829 2805 13863 2839
rect 16313 2805 16347 2839
rect 18337 2805 18371 2839
rect 25513 2805 25547 2839
rect 27721 2805 27755 2839
rect 2237 2601 2271 2635
rect 2605 2601 2639 2635
rect 3341 2601 3375 2635
rect 5733 2601 5767 2635
rect 11621 2601 11655 2635
rect 12081 2601 12115 2635
rect 12817 2601 12851 2635
rect 14105 2601 14139 2635
rect 14473 2601 14507 2635
rect 15209 2601 15243 2635
rect 16865 2601 16899 2635
rect 19625 2601 19659 2635
rect 23029 2601 23063 2635
rect 27077 2601 27111 2635
rect 6285 2533 6319 2567
rect 6745 2533 6779 2567
rect 7450 2533 7484 2567
rect 11161 2533 11195 2567
rect 15730 2533 15764 2567
rect 1501 2465 1535 2499
rect 2789 2465 2823 2499
rect 3893 2465 3927 2499
rect 4620 2465 4654 2499
rect 7205 2465 7239 2499
rect 11437 2465 11471 2499
rect 13185 2465 13219 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 19441 2465 19475 2499
rect 19993 2465 20027 2499
rect 22845 2465 22879 2499
rect 23397 2465 23431 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 25697 2465 25731 2499
rect 26249 2465 26283 2499
rect 26893 2465 26927 2499
rect 27445 2465 27479 2499
rect 1777 2397 1811 2431
rect 4353 2397 4387 2431
rect 13829 2397 13863 2431
rect 13369 2329 13403 2363
rect 2973 2261 3007 2295
rect 8585 2261 8619 2295
rect 9965 2261 9999 2295
rect 18521 2261 18555 2295
rect 24777 2261 24811 2295
rect 25881 2261 25915 2295
<< metal1 >>
rect 4062 22312 4068 22364
rect 4120 22352 4126 22364
rect 10597 22355 10655 22361
rect 10597 22352 10609 22355
rect 4120 22324 10609 22352
rect 4120 22312 4126 22324
rect 10597 22321 10609 22324
rect 10643 22321 10655 22355
rect 10597 22315 10655 22321
rect 2958 22176 2964 22228
rect 3016 22216 3022 22228
rect 13170 22216 13176 22228
rect 3016 22188 13176 22216
rect 3016 22176 3022 22188
rect 13170 22176 13176 22188
rect 13228 22176 13234 22228
rect 12526 22108 12532 22160
rect 12584 22148 12590 22160
rect 24854 22148 24860 22160
rect 12584 22120 24860 22148
rect 12584 22108 12590 22120
rect 24854 22108 24860 22120
rect 24912 22108 24918 22160
rect 10594 22012 10600 22024
rect 10555 21984 10600 22012
rect 10594 21972 10600 21984
rect 10652 21972 10658 22024
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 25314 21632 25320 21684
rect 25372 21672 25378 21684
rect 25682 21672 25688 21684
rect 25372 21644 25688 21672
rect 25372 21632 25378 21644
rect 25682 21632 25688 21644
rect 25740 21632 25746 21684
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 14182 21020 14188 21072
rect 14240 21060 14246 21072
rect 25774 21060 25780 21072
rect 14240 21032 25780 21060
rect 14240 21020 14246 21032
rect 25774 21020 25780 21032
rect 25832 21020 25838 21072
rect 3878 20952 3884 21004
rect 3936 20992 3942 21004
rect 13170 20992 13176 21004
rect 3936 20964 13176 20992
rect 3936 20952 3942 20964
rect 13170 20952 13176 20964
rect 13228 20952 13234 21004
rect 19245 20995 19303 21001
rect 19245 20961 19257 20995
rect 19291 20992 19303 20995
rect 20162 20992 20168 21004
rect 19291 20964 20168 20992
rect 19291 20961 19303 20964
rect 19245 20955 19303 20961
rect 20162 20952 20168 20964
rect 20220 20952 20226 21004
rect 21542 20992 21548 21004
rect 21503 20964 21548 20992
rect 21542 20952 21548 20964
rect 21600 20952 21606 21004
rect 3142 20884 3148 20936
rect 3200 20924 3206 20936
rect 25682 20924 25688 20936
rect 3200 20896 25688 20924
rect 3200 20884 3206 20896
rect 25682 20884 25688 20896
rect 25740 20884 25746 20936
rect 8202 20816 8208 20868
rect 8260 20856 8266 20868
rect 21729 20859 21787 20865
rect 21729 20856 21741 20859
rect 8260 20828 21741 20856
rect 8260 20816 8266 20828
rect 21729 20825 21741 20828
rect 21775 20825 21787 20859
rect 21729 20819 21787 20825
rect 5166 20748 5172 20800
rect 5224 20788 5230 20800
rect 19429 20791 19487 20797
rect 19429 20788 19441 20791
rect 5224 20760 19441 20788
rect 5224 20748 5230 20760
rect 19429 20757 19441 20760
rect 19475 20757 19487 20791
rect 19429 20751 19487 20757
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 8665 20587 8723 20593
rect 8665 20553 8677 20587
rect 8711 20584 8723 20587
rect 9582 20584 9588 20596
rect 8711 20556 9588 20584
rect 8711 20553 8723 20556
rect 8665 20547 8723 20553
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 10137 20587 10195 20593
rect 10137 20553 10149 20587
rect 10183 20584 10195 20587
rect 11330 20584 11336 20596
rect 10183 20556 11336 20584
rect 10183 20553 10195 20556
rect 10137 20547 10195 20553
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 19337 20587 19395 20593
rect 19337 20553 19349 20587
rect 19383 20584 19395 20587
rect 19426 20584 19432 20596
rect 19383 20556 19432 20584
rect 19383 20553 19395 20556
rect 19337 20547 19395 20553
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 21542 20584 21548 20596
rect 21503 20556 21548 20584
rect 21542 20544 21548 20556
rect 21600 20584 21606 20596
rect 22002 20584 22008 20596
rect 21600 20556 22008 20584
rect 21600 20544 21606 20556
rect 22002 20544 22008 20556
rect 22060 20544 22066 20596
rect 20622 20516 20628 20528
rect 20583 20488 20628 20516
rect 20622 20476 20628 20488
rect 20680 20476 20686 20528
rect 23842 20516 23848 20528
rect 23803 20488 23848 20516
rect 23842 20476 23848 20488
rect 23900 20476 23906 20528
rect 8481 20383 8539 20389
rect 8481 20349 8493 20383
rect 8527 20380 8539 20383
rect 8570 20380 8576 20392
rect 8527 20352 8576 20380
rect 8527 20349 8539 20352
rect 8481 20343 8539 20349
rect 8570 20340 8576 20352
rect 8628 20380 8634 20392
rect 9033 20383 9091 20389
rect 9033 20380 9045 20383
rect 8628 20352 9045 20380
rect 8628 20340 8634 20352
rect 9033 20349 9045 20352
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 12529 20383 12587 20389
rect 12529 20349 12541 20383
rect 12575 20380 12587 20383
rect 12710 20380 12716 20392
rect 12575 20352 12716 20380
rect 12575 20349 12587 20352
rect 12529 20343 12587 20349
rect 12710 20340 12716 20352
rect 12768 20380 12774 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 12768 20352 13093 20380
rect 12768 20340 12774 20352
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 16301 20383 16359 20389
rect 16301 20349 16313 20383
rect 16347 20380 16359 20383
rect 16945 20383 17003 20389
rect 16945 20380 16957 20383
rect 16347 20352 16957 20380
rect 16347 20349 16359 20352
rect 16301 20343 16359 20349
rect 16945 20349 16957 20352
rect 16991 20380 17003 20383
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 16991 20352 18061 20380
rect 16991 20349 17003 20352
rect 16945 20343 17003 20349
rect 18049 20349 18061 20352
rect 18095 20380 18107 20383
rect 18095 20352 18736 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 12710 20244 12716 20256
rect 12671 20216 12716 20244
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 16482 20244 16488 20256
rect 16443 20216 16488 20244
rect 16482 20204 16488 20216
rect 16540 20204 16546 20256
rect 18230 20244 18236 20256
rect 18191 20216 18236 20244
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 18708 20253 18736 20352
rect 18966 20340 18972 20392
rect 19024 20380 19030 20392
rect 19153 20383 19211 20389
rect 19153 20380 19165 20383
rect 19024 20352 19165 20380
rect 19024 20340 19030 20352
rect 19153 20349 19165 20352
rect 19199 20380 19211 20383
rect 19705 20383 19763 20389
rect 19705 20380 19717 20383
rect 19199 20352 19717 20380
rect 19199 20349 19211 20352
rect 19153 20343 19211 20349
rect 19705 20349 19717 20352
rect 19751 20349 19763 20383
rect 19705 20343 19763 20349
rect 20441 20383 20499 20389
rect 20441 20349 20453 20383
rect 20487 20380 20499 20383
rect 21085 20383 21143 20389
rect 21085 20380 21097 20383
rect 20487 20352 21097 20380
rect 20487 20349 20499 20352
rect 20441 20343 20499 20349
rect 21085 20349 21097 20352
rect 21131 20380 21143 20383
rect 21729 20383 21787 20389
rect 21729 20380 21741 20383
rect 21131 20352 21741 20380
rect 21131 20349 21143 20352
rect 21085 20343 21143 20349
rect 21729 20349 21741 20352
rect 21775 20380 21787 20383
rect 22278 20380 22284 20392
rect 21775 20352 22284 20380
rect 21775 20349 21787 20352
rect 21729 20343 21787 20349
rect 22278 20340 22284 20352
rect 22336 20340 22342 20392
rect 23658 20380 23664 20392
rect 23619 20352 23664 20380
rect 23658 20340 23664 20352
rect 23716 20380 23722 20392
rect 24213 20383 24271 20389
rect 24213 20380 24225 20383
rect 23716 20352 24225 20380
rect 23716 20340 23722 20352
rect 24213 20349 24225 20352
rect 24259 20349 24271 20383
rect 24213 20343 24271 20349
rect 20162 20312 20168 20324
rect 20075 20284 20168 20312
rect 20162 20272 20168 20284
rect 20220 20312 20226 20324
rect 20714 20312 20720 20324
rect 20220 20284 20720 20312
rect 20220 20272 20226 20284
rect 20714 20272 20720 20284
rect 20772 20272 20778 20324
rect 18693 20247 18751 20253
rect 18693 20213 18705 20247
rect 18739 20244 18751 20247
rect 18874 20244 18880 20256
rect 18739 20216 18880 20244
rect 18739 20213 18751 20216
rect 18693 20207 18751 20213
rect 18874 20204 18880 20216
rect 18932 20204 18938 20256
rect 21910 20244 21916 20256
rect 21871 20216 21916 20244
rect 21910 20204 21916 20216
rect 21968 20204 21974 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 18598 20040 18604 20052
rect 18559 20012 18604 20040
rect 18598 20000 18604 20012
rect 18656 20000 18662 20052
rect 21085 20043 21143 20049
rect 21085 20009 21097 20043
rect 21131 20040 21143 20043
rect 21542 20040 21548 20052
rect 21131 20012 21548 20040
rect 21131 20009 21143 20012
rect 21085 20003 21143 20009
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 17310 19904 17316 19916
rect 17271 19876 17316 19904
rect 17310 19864 17316 19876
rect 17368 19864 17374 19916
rect 18417 19907 18475 19913
rect 18417 19873 18429 19907
rect 18463 19904 18475 19907
rect 19426 19904 19432 19916
rect 18463 19876 19432 19904
rect 18463 19873 18475 19876
rect 18417 19867 18475 19873
rect 19426 19864 19432 19876
rect 19484 19904 19490 19916
rect 19521 19907 19579 19913
rect 19521 19904 19533 19907
rect 19484 19876 19533 19904
rect 19484 19864 19490 19876
rect 19521 19873 19533 19876
rect 19567 19873 19579 19907
rect 19521 19867 19579 19873
rect 20714 19864 20720 19916
rect 20772 19904 20778 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20772 19876 20913 19904
rect 20772 19864 20778 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 17494 19768 17500 19780
rect 17455 19740 17500 19768
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 19702 19768 19708 19780
rect 19663 19740 19708 19768
rect 19702 19728 19708 19740
rect 19760 19728 19766 19780
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 17310 19496 17316 19508
rect 17271 19468 17316 19496
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 16482 19360 16488 19372
rect 15804 19332 16488 19360
rect 15804 19320 15810 19332
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 17328 19360 17356 19456
rect 17402 19388 17408 19440
rect 17460 19428 17466 19440
rect 17770 19428 17776 19440
rect 17460 19400 17776 19428
rect 17460 19388 17466 19400
rect 17770 19388 17776 19400
rect 17828 19388 17834 19440
rect 19058 19360 19064 19372
rect 17328 19332 19064 19360
rect 19058 19320 19064 19332
rect 19116 19320 19122 19372
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14550 19292 14556 19304
rect 14332 19264 14556 19292
rect 14332 19252 14338 19264
rect 14550 19252 14556 19264
rect 14608 19252 14614 19304
rect 19426 19184 19432 19236
rect 19484 19184 19490 19236
rect 18509 19159 18567 19165
rect 18509 19125 18521 19159
rect 18555 19156 18567 19159
rect 19444 19156 19472 19184
rect 19521 19159 19579 19165
rect 19521 19156 19533 19159
rect 18555 19128 19533 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 19521 19125 19533 19128
rect 19567 19156 19579 19159
rect 19794 19156 19800 19168
rect 19567 19128 19800 19156
rect 19567 19125 19579 19128
rect 19521 19119 19579 19125
rect 19794 19116 19800 19128
rect 19852 19116 19858 19168
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 20901 19159 20959 19165
rect 20901 19156 20913 19159
rect 20772 19128 20913 19156
rect 20772 19116 20778 19128
rect 20901 19125 20913 19128
rect 20947 19125 20959 19159
rect 20901 19119 20959 19125
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 21358 16028 21364 16040
rect 19392 16000 21364 16028
rect 19392 15988 19398 16000
rect 21358 15988 21364 16000
rect 21416 15988 21422 16040
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 11790 14532 11796 14544
rect 11751 14504 11796 14532
rect 11790 14492 11796 14504
rect 11848 14492 11854 14544
rect 11882 14464 11888 14476
rect 11843 14436 11888 14464
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 12158 14396 12164 14408
rect 12115 14368 12164 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 11425 14263 11483 14269
rect 11425 14229 11437 14263
rect 11471 14260 11483 14263
rect 12434 14260 12440 14272
rect 11471 14232 12440 14260
rect 11471 14229 11483 14232
rect 11425 14223 11483 14229
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11790 14056 11796 14068
rect 11563 14028 11796 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11940 14028 12173 14056
rect 11940 14016 11946 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 12158 13920 12164 13932
rect 11808 13892 12164 13920
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 2682 13852 2688 13864
rect 2547 13824 2688 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 2682 13812 2688 13824
rect 2740 13812 2746 13864
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 11808 13793 11836 13892
rect 12158 13880 12164 13892
rect 12216 13920 12222 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 12216 13892 13553 13920
rect 12216 13880 12222 13892
rect 13541 13889 13553 13892
rect 13587 13920 13599 13923
rect 13587 13892 13768 13920
rect 13587 13889 13599 13892
rect 13541 13883 13599 13889
rect 13630 13852 13636 13864
rect 13591 13824 13636 13852
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 13740 13852 13768 13892
rect 13906 13861 13912 13864
rect 13900 13852 13912 13861
rect 13740 13824 13912 13852
rect 13900 13815 13912 13824
rect 13906 13812 13912 13815
rect 13964 13812 13970 13864
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 10836 13756 11805 13784
rect 10836 13744 10842 13756
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 11793 13747 11851 13753
rect 1670 13716 1676 13728
rect 1631 13688 1676 13716
rect 1670 13676 1676 13688
rect 1728 13676 1734 13728
rect 3053 13719 3111 13725
rect 3053 13685 3065 13719
rect 3099 13716 3111 13719
rect 4890 13716 4896 13728
rect 3099 13688 4896 13716
rect 3099 13685 3111 13688
rect 3053 13679 3111 13685
rect 4890 13676 4896 13688
rect 4948 13676 4954 13728
rect 10226 13716 10232 13728
rect 10187 13688 10232 13716
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 15010 13716 15016 13728
rect 14971 13688 15016 13716
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 1728 13484 2421 13512
rect 1728 13472 1734 13484
rect 2409 13481 2421 13484
rect 2455 13481 2467 13515
rect 2409 13475 2467 13481
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 2774 13512 2780 13524
rect 2556 13484 2780 13512
rect 2556 13472 2562 13484
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12161 13515 12219 13521
rect 12161 13512 12173 13515
rect 11940 13484 12173 13512
rect 11940 13472 11946 13484
rect 12161 13481 12173 13484
rect 12207 13481 12219 13515
rect 12161 13475 12219 13481
rect 9490 13404 9496 13456
rect 9548 13444 9554 13456
rect 12250 13444 12256 13456
rect 9548 13416 12256 13444
rect 9548 13404 9554 13416
rect 12250 13404 12256 13416
rect 12308 13444 12314 13456
rect 12621 13447 12679 13453
rect 12621 13444 12633 13447
rect 12308 13416 12633 13444
rect 12308 13404 12314 13416
rect 12621 13413 12633 13416
rect 12667 13413 12679 13447
rect 12621 13407 12679 13413
rect 2682 13336 2688 13388
rect 2740 13376 2746 13388
rect 2777 13379 2835 13385
rect 2777 13376 2789 13379
rect 2740 13348 2789 13376
rect 2740 13336 2746 13348
rect 2777 13345 2789 13348
rect 2823 13376 2835 13379
rect 4522 13376 4528 13388
rect 2823 13348 4528 13376
rect 2823 13345 2835 13348
rect 2777 13339 2835 13345
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 5258 13385 5264 13388
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 5252 13376 5264 13385
rect 4663 13348 5264 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 5252 13339 5264 13348
rect 5258 13336 5264 13339
rect 5316 13336 5322 13388
rect 9950 13385 9956 13388
rect 9944 13376 9956 13385
rect 9911 13348 9956 13376
rect 9944 13339 9956 13348
rect 9950 13336 9956 13339
rect 10008 13336 10014 13388
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 12529 13379 12587 13385
rect 12529 13376 12541 13379
rect 11848 13348 12541 13376
rect 11848 13336 11854 13348
rect 12529 13345 12541 13348
rect 12575 13376 12587 13379
rect 12894 13376 12900 13388
rect 12575 13348 12900 13376
rect 12575 13345 12587 13348
rect 12529 13339 12587 13345
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13308 2375 13311
rect 2866 13308 2872 13320
rect 2363 13280 2872 13308
rect 2363 13277 2375 13280
rect 2317 13271 2375 13277
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 3050 13308 3056 13320
rect 3011 13280 3056 13308
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 4982 13308 4988 13320
rect 4943 13280 4988 13308
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 7650 13268 7656 13320
rect 7708 13308 7714 13320
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 7708 13280 7757 13308
rect 7708 13268 7714 13280
rect 7745 13277 7757 13280
rect 7791 13308 7803 13311
rect 9493 13311 9551 13317
rect 9493 13308 9505 13311
rect 7791 13280 9505 13308
rect 7791 13277 7803 13280
rect 7745 13271 7803 13277
rect 9493 13277 9505 13280
rect 9539 13308 9551 13311
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9539 13280 9689 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 12710 13308 12716 13320
rect 12671 13280 12716 13308
rect 9677 13271 9735 13277
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 1854 13172 1860 13184
rect 1719 13144 1860 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 6362 13172 6368 13184
rect 6323 13144 6368 13172
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10836 13144 11069 13172
rect 10836 13132 10842 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 13725 13175 13783 13181
rect 13725 13172 13737 13175
rect 13688 13144 13737 13172
rect 13688 13132 13694 13144
rect 13725 13141 13737 13144
rect 13771 13172 13783 13175
rect 14918 13172 14924 13184
rect 13771 13144 14924 13172
rect 13771 13141 13783 13144
rect 13725 13135 13783 13141
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 2866 12928 2872 12980
rect 2924 12968 2930 12980
rect 2961 12971 3019 12977
rect 2961 12968 2973 12971
rect 2924 12940 2973 12968
rect 2924 12928 2930 12940
rect 2961 12937 2973 12940
rect 3007 12937 3019 12971
rect 3510 12968 3516 12980
rect 2961 12931 3019 12937
rect 3436 12940 3516 12968
rect 1397 12903 1455 12909
rect 1397 12869 1409 12903
rect 1443 12900 1455 12903
rect 2590 12900 2596 12912
rect 1443 12872 2596 12900
rect 1443 12869 1455 12872
rect 1397 12863 1455 12869
rect 2590 12860 2596 12872
rect 2648 12860 2654 12912
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 2038 12832 2044 12844
rect 1999 12804 2044 12832
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 3436 12841 3464 12940
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 4522 12968 4528 12980
rect 4483 12940 4528 12968
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 12250 12968 12256 12980
rect 12211 12940 12256 12968
rect 12250 12928 12256 12940
rect 12308 12968 12314 12980
rect 17954 12968 17960 12980
rect 12308 12940 17960 12968
rect 12308 12928 12314 12940
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 9033 12903 9091 12909
rect 9033 12869 9045 12903
rect 9079 12900 9091 12903
rect 9769 12903 9827 12909
rect 9769 12900 9781 12903
rect 9079 12872 9781 12900
rect 9079 12869 9091 12872
rect 9033 12863 9091 12869
rect 9769 12869 9781 12872
rect 9815 12900 9827 12903
rect 9950 12900 9956 12912
rect 9815 12872 9956 12900
rect 9815 12869 9827 12872
rect 9769 12863 9827 12869
rect 9950 12860 9956 12872
rect 10008 12900 10014 12912
rect 10134 12900 10140 12912
rect 10008 12872 10140 12900
rect 10008 12860 10014 12872
rect 10134 12860 10140 12872
rect 10192 12900 10198 12912
rect 11517 12903 11575 12909
rect 11517 12900 11529 12903
rect 10192 12872 11529 12900
rect 10192 12860 10198 12872
rect 11517 12869 11529 12872
rect 11563 12900 11575 12903
rect 12710 12900 12716 12912
rect 11563 12872 12716 12900
rect 11563 12869 11575 12872
rect 11517 12863 11575 12869
rect 12710 12860 12716 12872
rect 12768 12860 12774 12912
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12801 3479 12835
rect 3602 12832 3608 12844
rect 3515 12804 3608 12832
rect 3421 12795 3479 12801
rect 1670 12724 1676 12776
rect 1728 12764 1734 12776
rect 1765 12767 1823 12773
rect 1765 12764 1777 12767
rect 1728 12736 1777 12764
rect 1728 12724 1734 12736
rect 1765 12733 1777 12736
rect 1811 12733 1823 12767
rect 1765 12727 1823 12733
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 2869 12767 2927 12773
rect 2869 12764 2881 12767
rect 2832 12736 2881 12764
rect 2832 12724 2838 12736
rect 2869 12733 2881 12736
rect 2915 12764 2927 12767
rect 3326 12764 3332 12776
rect 2915 12736 3332 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 3326 12724 3332 12736
rect 3384 12724 3390 12776
rect 2501 12699 2559 12705
rect 2501 12665 2513 12699
rect 2547 12696 2559 12699
rect 3436 12696 3464 12795
rect 3602 12792 3608 12804
rect 3660 12832 3666 12844
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 3660 12804 5181 12832
rect 3660 12792 3666 12804
rect 5169 12801 5181 12804
rect 5215 12832 5227 12835
rect 5258 12832 5264 12844
rect 5215 12804 5264 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5258 12792 5264 12804
rect 5316 12832 5322 12844
rect 7650 12832 7656 12844
rect 5316 12804 5672 12832
rect 7611 12804 7656 12832
rect 5316 12792 5322 12804
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 4890 12764 4896 12776
rect 4580 12736 4896 12764
rect 4580 12724 4586 12736
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12764 5043 12767
rect 5074 12764 5080 12776
rect 5031 12736 5080 12764
rect 5031 12733 5043 12736
rect 4985 12727 5043 12733
rect 4430 12696 4436 12708
rect 2547 12668 3464 12696
rect 4343 12668 4436 12696
rect 2547 12665 2559 12668
rect 2501 12659 2559 12665
rect 3344 12640 3372 12668
rect 4430 12656 4436 12668
rect 4488 12696 4494 12708
rect 5000 12696 5028 12727
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 4488 12668 5028 12696
rect 4488 12656 4494 12668
rect 3326 12588 3332 12640
rect 3384 12588 3390 12640
rect 4062 12628 4068 12640
rect 4023 12600 4068 12628
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 5644 12637 5672 12804
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 10226 12832 10232 12844
rect 9732 12804 10232 12832
rect 9732 12792 9738 12804
rect 10226 12792 10232 12804
rect 10284 12832 10290 12844
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 10284 12804 10609 12832
rect 10284 12792 10290 12804
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10778 12832 10784 12844
rect 10739 12804 10784 12832
rect 10597 12795 10655 12801
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12952 12804 13001 12832
rect 12952 12792 12958 12804
rect 12989 12801 13001 12804
rect 13035 12832 13047 12835
rect 14737 12835 14795 12841
rect 14737 12832 14749 12835
rect 13035 12804 14749 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 14737 12801 14749 12804
rect 14783 12832 14795 12835
rect 14783 12804 15056 12832
rect 14783 12801 14795 12804
rect 14737 12795 14795 12801
rect 15028 12776 15056 12804
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12492 12736 12817 12764
rect 12492 12724 12498 12736
rect 12805 12733 12817 12736
rect 12851 12764 12863 12767
rect 13078 12764 13084 12776
rect 12851 12736 13084 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 14918 12764 14924 12776
rect 14879 12736 14924 12764
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 15010 12724 15016 12776
rect 15068 12764 15074 12776
rect 15177 12767 15235 12773
rect 15177 12764 15189 12767
rect 15068 12736 15189 12764
rect 15068 12724 15074 12736
rect 15177 12733 15189 12736
rect 15223 12733 15235 12767
rect 15177 12727 15235 12733
rect 7898 12699 7956 12705
rect 7898 12696 7910 12699
rect 7484 12668 7910 12696
rect 5629 12631 5687 12637
rect 5629 12597 5641 12631
rect 5675 12628 5687 12631
rect 6822 12628 6828 12640
rect 5675 12600 6828 12628
rect 5675 12597 5687 12600
rect 5629 12591 5687 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7190 12588 7196 12640
rect 7248 12628 7254 12640
rect 7484 12637 7512 12668
rect 7898 12665 7910 12668
rect 7944 12665 7956 12699
rect 7898 12659 7956 12665
rect 10152 12668 12940 12696
rect 10152 12637 10180 12668
rect 7469 12631 7527 12637
rect 7469 12628 7481 12631
rect 7248 12600 7481 12628
rect 7248 12588 7254 12600
rect 7469 12597 7481 12600
rect 7515 12597 7527 12631
rect 7469 12591 7527 12597
rect 10137 12631 10195 12637
rect 10137 12597 10149 12631
rect 10183 12597 10195 12631
rect 10502 12628 10508 12640
rect 10463 12600 10508 12628
rect 10137 12591 10195 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 12434 12628 12440 12640
rect 12395 12600 12440 12628
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 12912 12637 12940 12668
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13449 12631 13507 12637
rect 13449 12628 13461 12631
rect 12943 12600 13461 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13449 12597 13461 12600
rect 13495 12597 13507 12631
rect 13449 12591 13507 12597
rect 16301 12631 16359 12637
rect 16301 12597 16313 12631
rect 16347 12628 16359 12631
rect 16390 12628 16396 12640
rect 16347 12600 16396 12628
rect 16347 12597 16359 12600
rect 16301 12591 16359 12597
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 1912 12396 2421 12424
rect 1912 12384 1918 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 2409 12387 2467 12393
rect 3513 12427 3571 12433
rect 3513 12393 3525 12427
rect 3559 12424 3571 12427
rect 3602 12424 3608 12436
rect 3559 12396 3608 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 4522 12424 4528 12436
rect 4483 12396 4528 12424
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 4982 12424 4988 12436
rect 4943 12396 4988 12424
rect 4982 12384 4988 12396
rect 5040 12384 5046 12436
rect 7190 12424 7196 12436
rect 7151 12396 7196 12424
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 9493 12427 9551 12433
rect 9493 12393 9505 12427
rect 9539 12424 9551 12427
rect 9677 12427 9735 12433
rect 9677 12424 9689 12427
rect 9539 12396 9689 12424
rect 9539 12393 9551 12396
rect 9493 12387 9551 12393
rect 9677 12393 9689 12396
rect 9723 12424 9735 12427
rect 10502 12424 10508 12436
rect 9723 12396 10508 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 10502 12384 10508 12396
rect 10560 12384 10566 12436
rect 10778 12424 10784 12436
rect 10739 12396 10784 12424
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 12161 12427 12219 12433
rect 12161 12424 12173 12427
rect 11480 12396 12173 12424
rect 11480 12384 11486 12396
rect 12161 12393 12173 12396
rect 12207 12424 12219 12427
rect 12434 12424 12440 12436
rect 12207 12396 12440 12424
rect 12207 12393 12219 12396
rect 12161 12387 12219 12393
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 12894 12424 12900 12436
rect 12851 12396 12900 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13078 12424 13084 12436
rect 13039 12396 13084 12424
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13633 12427 13691 12433
rect 13633 12393 13645 12427
rect 13679 12424 13691 12427
rect 13722 12424 13728 12436
rect 13679 12396 13728 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 1673 12359 1731 12365
rect 1673 12325 1685 12359
rect 1719 12356 1731 12359
rect 2038 12356 2044 12368
rect 1719 12328 2044 12356
rect 1719 12325 1731 12328
rect 1673 12319 1731 12325
rect 2038 12316 2044 12328
rect 2096 12316 2102 12368
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2774 12288 2780 12300
rect 2363 12260 2780 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2774 12248 2780 12260
rect 2832 12288 2838 12300
rect 5000 12288 5028 12384
rect 6080 12359 6138 12365
rect 6080 12325 6092 12359
rect 6126 12356 6138 12359
rect 6362 12356 6368 12368
rect 6126 12328 6368 12356
rect 6126 12325 6138 12328
rect 6080 12319 6138 12325
rect 6362 12316 6368 12328
rect 6420 12316 6426 12368
rect 16942 12356 16948 12368
rect 16500 12328 16948 12356
rect 5810 12288 5816 12300
rect 2832 12260 2877 12288
rect 5000 12260 5816 12288
rect 2832 12248 2838 12260
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10686 12288 10692 12300
rect 10091 12260 10692 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 12069 12291 12127 12297
rect 12069 12257 12081 12291
rect 12115 12288 12127 12291
rect 12434 12288 12440 12300
rect 12115 12260 12440 12288
rect 12115 12257 12127 12260
rect 12069 12251 12127 12257
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 13538 12248 13544 12300
rect 13596 12288 13602 12300
rect 13725 12291 13783 12297
rect 13725 12288 13737 12291
rect 13596 12260 13737 12288
rect 13596 12248 13602 12260
rect 13725 12257 13737 12260
rect 13771 12257 13783 12291
rect 13725 12251 13783 12257
rect 14918 12248 14924 12300
rect 14976 12288 14982 12300
rect 16500 12297 16528 12328
rect 16942 12316 16948 12328
rect 17000 12316 17006 12368
rect 15013 12291 15071 12297
rect 15013 12288 15025 12291
rect 14976 12260 15025 12288
rect 14976 12248 14982 12260
rect 15013 12257 15025 12260
rect 15059 12288 15071 12291
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 15059 12260 16497 12288
rect 15059 12257 15071 12260
rect 15013 12251 15071 12257
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 16741 12291 16799 12297
rect 16741 12288 16753 12291
rect 16632 12260 16753 12288
rect 16632 12248 16638 12260
rect 16741 12257 16753 12260
rect 16787 12257 16799 12291
rect 16741 12251 16799 12257
rect 2866 12220 2872 12232
rect 2827 12192 2872 12220
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 3050 12220 3056 12232
rect 2963 12192 3056 12220
rect 3050 12180 3056 12192
rect 3108 12220 3114 12232
rect 4062 12220 4068 12232
rect 3108 12192 4068 12220
rect 3108 12180 3114 12192
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 10134 12220 10140 12232
rect 9088 12192 10140 12220
rect 9088 12180 9094 12192
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 12342 12220 12348 12232
rect 10284 12192 10329 12220
rect 12303 12192 12348 12220
rect 10284 12180 10290 12192
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 13814 12220 13820 12232
rect 13775 12192 13820 12220
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 26234 12112 26240 12164
rect 26292 12152 26298 12164
rect 26510 12152 26516 12164
rect 26292 12124 26516 12152
rect 26292 12112 26298 12124
rect 26510 12112 26516 12124
rect 26568 12112 26574 12164
rect 11698 12084 11704 12096
rect 11659 12056 11704 12084
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 12802 12044 12808 12096
rect 12860 12084 12866 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 12860 12056 13277 12084
rect 12860 12044 12866 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 13265 12047 13323 12053
rect 15470 12044 15476 12096
rect 15528 12084 15534 12096
rect 16482 12084 16488 12096
rect 15528 12056 16488 12084
rect 15528 12044 15534 12056
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 17865 12087 17923 12093
rect 17865 12053 17877 12087
rect 17911 12084 17923 12087
rect 18230 12084 18236 12096
rect 17911 12056 18236 12084
rect 17911 12053 17923 12056
rect 17865 12047 17923 12053
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 18506 12084 18512 12096
rect 18467 12056 18512 12084
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 2593 11883 2651 11889
rect 2593 11880 2605 11883
rect 2556 11852 2605 11880
rect 2556 11840 2562 11852
rect 2593 11849 2605 11852
rect 2639 11849 2651 11883
rect 2593 11843 2651 11849
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 2832 11852 2877 11880
rect 2832 11840 2838 11852
rect 3602 11840 3608 11892
rect 3660 11880 3666 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3660 11852 3801 11880
rect 3660 11840 3666 11852
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4249 11883 4307 11889
rect 4249 11880 4261 11883
rect 4120 11852 4261 11880
rect 4120 11840 4126 11852
rect 4249 11849 4261 11852
rect 4295 11880 4307 11883
rect 5905 11883 5963 11889
rect 5905 11880 5917 11883
rect 4295 11852 5917 11880
rect 4295 11849 4307 11852
rect 4249 11843 4307 11849
rect 5905 11849 5917 11852
rect 5951 11880 5963 11883
rect 6362 11880 6368 11892
rect 5951 11852 6368 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 9398 11880 9404 11892
rect 9359 11852 9404 11880
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9582 11880 9588 11892
rect 9543 11852 9588 11880
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 11422 11880 11428 11892
rect 11383 11852 11428 11880
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 16574 11880 16580 11892
rect 12492 11852 12537 11880
rect 16535 11852 16580 11880
rect 12492 11840 12498 11852
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 18230 11880 18236 11892
rect 18191 11852 18236 11880
rect 18230 11840 18236 11852
rect 18288 11880 18294 11892
rect 18690 11880 18696 11892
rect 18288 11852 18696 11880
rect 18288 11840 18294 11852
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 2041 11747 2099 11753
rect 2041 11744 2053 11747
rect 1412 11716 2053 11744
rect 1412 11685 1440 11716
rect 2041 11713 2053 11716
rect 2087 11744 2099 11747
rect 2682 11744 2688 11756
rect 2087 11716 2688 11744
rect 2087 11713 2099 11716
rect 2041 11707 2099 11713
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11744 3479 11747
rect 3620 11744 3648 11840
rect 5810 11772 5816 11824
rect 5868 11812 5874 11824
rect 6181 11815 6239 11821
rect 6181 11812 6193 11815
rect 5868 11784 6193 11812
rect 5868 11772 5874 11784
rect 6181 11781 6193 11784
rect 6227 11812 6239 11815
rect 6730 11812 6736 11824
rect 6227 11784 6736 11812
rect 6227 11781 6239 11784
rect 6181 11775 6239 11781
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 11793 11815 11851 11821
rect 11793 11781 11805 11815
rect 11839 11812 11851 11815
rect 12342 11812 12348 11824
rect 11839 11784 12348 11812
rect 11839 11781 11851 11784
rect 11793 11775 11851 11781
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 3467 11716 3648 11744
rect 8757 11747 8815 11753
rect 3467 11713 3479 11716
rect 3421 11707 3479 11713
rect 8757 11713 8769 11747
rect 8803 11744 8815 11747
rect 10137 11747 10195 11753
rect 10137 11744 10149 11747
rect 8803 11716 10149 11744
rect 8803 11713 8815 11716
rect 8757 11707 8815 11713
rect 10137 11713 10149 11716
rect 10183 11744 10195 11747
rect 10226 11744 10232 11756
rect 10183 11716 10232 11744
rect 10183 11713 10195 11716
rect 10137 11707 10195 11713
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12894 11744 12900 11756
rect 12299 11716 12900 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12894 11704 12900 11716
rect 12952 11744 12958 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12952 11716 13001 11744
rect 12952 11704 12958 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11645 1455 11679
rect 1397 11639 1455 11645
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 9766 11676 9772 11688
rect 9456 11648 9772 11676
rect 9456 11636 9462 11648
rect 9766 11636 9772 11648
rect 9824 11676 9830 11688
rect 10045 11679 10103 11685
rect 10045 11676 10057 11679
rect 9824 11648 10057 11676
rect 9824 11636 9830 11648
rect 10045 11645 10057 11648
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 12158 11636 12164 11688
rect 12216 11676 12222 11688
rect 12802 11676 12808 11688
rect 12216 11648 12808 11676
rect 12216 11636 12222 11648
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13814 11676 13820 11688
rect 13504 11648 13820 11676
rect 13504 11636 13510 11648
rect 13814 11636 13820 11648
rect 13872 11676 13878 11688
rect 14185 11679 14243 11685
rect 14185 11676 14197 11679
rect 13872 11648 14197 11676
rect 13872 11636 13878 11648
rect 14185 11645 14197 11648
rect 14231 11645 14243 11679
rect 16942 11676 16948 11688
rect 16855 11648 16948 11676
rect 14185 11639 14243 11645
rect 16942 11636 16948 11648
rect 17000 11676 17006 11688
rect 18417 11679 18475 11685
rect 18417 11676 18429 11679
rect 17000 11648 18429 11676
rect 17000 11636 17006 11648
rect 18417 11645 18429 11648
rect 18463 11676 18475 11679
rect 18506 11676 18512 11688
rect 18463 11648 18512 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 18690 11685 18696 11688
rect 18684 11676 18696 11685
rect 18651 11648 18696 11676
rect 18684 11639 18696 11648
rect 18690 11636 18696 11639
rect 18748 11636 18754 11688
rect 26418 11676 26424 11688
rect 26379 11648 26424 11676
rect 26418 11636 26424 11648
rect 26476 11676 26482 11688
rect 26973 11679 27031 11685
rect 26973 11676 26985 11679
rect 26476 11648 26985 11676
rect 26476 11636 26482 11648
rect 26973 11645 26985 11648
rect 27019 11645 27031 11679
rect 26973 11639 27031 11645
rect 3145 11611 3203 11617
rect 3145 11577 3157 11611
rect 3191 11608 3203 11611
rect 3326 11608 3332 11620
rect 3191 11580 3332 11608
rect 3191 11577 3203 11580
rect 3145 11571 3203 11577
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 2498 11500 2504 11552
rect 2556 11540 2562 11552
rect 3160 11540 3188 11571
rect 3326 11568 3332 11580
rect 3384 11568 3390 11620
rect 9030 11608 9036 11620
rect 8991 11580 9036 11608
rect 9030 11568 9036 11580
rect 9088 11568 9094 11620
rect 13538 11608 13544 11620
rect 13499 11580 13544 11608
rect 13538 11568 13544 11580
rect 13596 11568 13602 11620
rect 2556 11512 3188 11540
rect 3237 11543 3295 11549
rect 2556 11500 2562 11512
rect 3237 11509 3249 11543
rect 3283 11540 3295 11543
rect 3418 11540 3424 11552
rect 3283 11512 3424 11540
rect 3283 11509 3295 11512
rect 3237 11503 3295 11509
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 9950 11540 9956 11552
rect 9911 11512 9956 11540
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10686 11540 10692 11552
rect 10647 11512 10692 11540
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13078 11500 13084 11552
rect 13136 11540 13142 11552
rect 13722 11540 13728 11552
rect 13136 11512 13728 11540
rect 13136 11500 13142 11512
rect 13722 11500 13728 11512
rect 13780 11540 13786 11552
rect 13817 11543 13875 11549
rect 13817 11540 13829 11543
rect 13780 11512 13829 11540
rect 13780 11500 13786 11512
rect 13817 11509 13829 11512
rect 13863 11509 13875 11543
rect 13817 11503 13875 11509
rect 19426 11500 19432 11552
rect 19484 11540 19490 11552
rect 19797 11543 19855 11549
rect 19797 11540 19809 11543
rect 19484 11512 19809 11540
rect 19484 11500 19490 11512
rect 19797 11509 19809 11512
rect 19843 11509 19855 11543
rect 26602 11540 26608 11552
rect 26563 11512 26608 11540
rect 19797 11503 19855 11509
rect 26602 11500 26608 11512
rect 26660 11500 26666 11552
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 2363 11308 2421 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2409 11305 2421 11308
rect 2455 11336 2467 11339
rect 2866 11336 2872 11348
rect 2455 11308 2872 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3418 11336 3424 11348
rect 3379 11308 3424 11336
rect 3418 11296 3424 11308
rect 3476 11336 3482 11348
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 3476 11308 4077 11336
rect 3476 11296 3482 11308
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4065 11299 4123 11305
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 6972 11308 8125 11336
rect 6972 11296 6978 11308
rect 8113 11305 8125 11308
rect 8159 11305 8171 11339
rect 10226 11336 10232 11348
rect 10187 11308 10232 11336
rect 8113 11299 8171 11305
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 11793 11339 11851 11345
rect 11793 11305 11805 11339
rect 11839 11336 11851 11339
rect 12434 11336 12440 11348
rect 11839 11308 12440 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 12529 11339 12587 11345
rect 12529 11305 12541 11339
rect 12575 11336 12587 11339
rect 12894 11336 12900 11348
rect 12575 11308 12900 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 13357 11339 13415 11345
rect 13357 11305 13369 11339
rect 13403 11336 13415 11339
rect 13538 11336 13544 11348
rect 13403 11308 13544 11336
rect 13403 11305 13415 11308
rect 13357 11299 13415 11305
rect 13538 11296 13544 11308
rect 13596 11336 13602 11348
rect 13998 11336 14004 11348
rect 13596 11308 14004 11336
rect 13596 11296 13602 11308
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 7000 11271 7058 11277
rect 7000 11237 7012 11271
rect 7046 11268 7058 11271
rect 7098 11268 7104 11280
rect 7046 11240 7104 11268
rect 7046 11237 7058 11240
rect 7000 11231 7058 11237
rect 7098 11228 7104 11240
rect 7156 11228 7162 11280
rect 12158 11268 12164 11280
rect 12119 11240 12164 11268
rect 12158 11228 12164 11240
rect 12216 11228 12222 11280
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 4433 11203 4491 11209
rect 2832 11172 2877 11200
rect 2832 11160 2838 11172
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4614 11200 4620 11212
rect 4479 11172 4620 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 6730 11200 6736 11212
rect 6691 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 13262 11200 13268 11212
rect 13223 11172 13268 11200
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 17678 11200 17684 11212
rect 17368 11172 17684 11200
rect 17368 11160 17374 11172
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 26510 11200 26516 11212
rect 26471 11172 26516 11200
rect 26510 11160 26516 11172
rect 26568 11160 26574 11212
rect 2866 11132 2872 11144
rect 2827 11104 2872 11132
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3602 11132 3608 11144
rect 3099 11104 3608 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 2406 11024 2412 11076
rect 2464 11064 2470 11076
rect 3068 11064 3096 11095
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 4522 11132 4528 11144
rect 4396 11104 4528 11132
rect 4396 11092 4402 11104
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 4890 11132 4896 11144
rect 4755 11104 4896 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 13446 11132 13452 11144
rect 13407 11104 13452 11132
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 17402 11092 17408 11144
rect 17460 11132 17466 11144
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 17460 11104 17785 11132
rect 17460 11092 17466 11104
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11132 18015 11135
rect 18230 11132 18236 11144
rect 18003 11104 18236 11132
rect 18003 11101 18015 11104
rect 17957 11095 18015 11101
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 9950 11064 9956 11076
rect 2464 11036 3096 11064
rect 9863 11036 9956 11064
rect 2464 11024 2470 11036
rect 9950 11024 9956 11036
rect 10008 11064 10014 11076
rect 10410 11064 10416 11076
rect 10008 11036 10416 11064
rect 10008 11024 10014 11036
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 16482 11064 16488 11076
rect 16443 11036 16488 11064
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 26694 11064 26700 11076
rect 26655 11036 26700 11064
rect 26694 11024 26700 11036
rect 26752 11024 26758 11076
rect 16758 10956 16764 11008
rect 16816 10996 16822 11008
rect 17313 10999 17371 11005
rect 17313 10996 17325 10999
rect 16816 10968 17325 10996
rect 16816 10956 16822 10968
rect 17313 10965 17325 10968
rect 17359 10965 17371 10999
rect 18414 10996 18420 11008
rect 18375 10968 18420 10996
rect 17313 10959 17371 10965
rect 18414 10956 18420 10968
rect 18472 10956 18478 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 2038 10792 2044 10804
rect 1999 10764 2044 10792
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2406 10792 2412 10804
rect 2367 10764 2412 10792
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 2832 10764 3249 10792
rect 2832 10752 2838 10764
rect 3237 10761 3249 10764
rect 3283 10761 3295 10795
rect 3237 10755 3295 10761
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 6972 10764 7389 10792
rect 6972 10752 6978 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 7377 10755 7435 10761
rect 12989 10795 13047 10801
rect 12989 10761 13001 10795
rect 13035 10792 13047 10795
rect 13262 10792 13268 10804
rect 13035 10764 13268 10792
rect 13035 10761 13047 10764
rect 12989 10755 13047 10761
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 13538 10792 13544 10804
rect 13499 10764 13544 10792
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 26510 10792 26516 10804
rect 26471 10764 26516 10792
rect 26510 10752 26516 10764
rect 26568 10752 26574 10804
rect 18049 10727 18107 10733
rect 18049 10724 18061 10727
rect 16868 10696 18061 10724
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 3881 10659 3939 10665
rect 3881 10656 3893 10659
rect 2823 10628 3893 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 3881 10625 3893 10628
rect 3927 10656 3939 10659
rect 4890 10656 4896 10668
rect 3927 10628 4896 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 9950 10656 9956 10668
rect 9863 10628 9956 10656
rect 9950 10616 9956 10628
rect 10008 10656 10014 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10008 10628 10609 10656
rect 10008 10616 10014 10628
rect 10597 10625 10609 10628
rect 10643 10656 10655 10659
rect 10870 10656 10876 10668
rect 10643 10628 10876 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 13078 10656 13084 10668
rect 13039 10628 13084 10656
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 16868 10665 16896 10696
rect 18049 10693 18061 10696
rect 18095 10693 18107 10727
rect 18049 10687 18107 10693
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16632 10628 16865 10656
rect 16632 10616 16638 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 17034 10656 17040 10668
rect 16995 10628 17040 10656
rect 16853 10619 16911 10625
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 17770 10656 17776 10668
rect 17731 10628 17776 10656
rect 17770 10616 17776 10628
rect 17828 10616 17834 10668
rect 18230 10616 18236 10668
rect 18288 10656 18294 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18288 10628 18613 10656
rect 18288 10616 18294 10628
rect 18601 10625 18613 10628
rect 18647 10656 18659 10659
rect 18690 10656 18696 10668
rect 18647 10628 18696 10656
rect 18647 10625 18659 10628
rect 18601 10619 18659 10625
rect 18690 10616 18696 10628
rect 18748 10656 18754 10668
rect 19061 10659 19119 10665
rect 19061 10656 19073 10659
rect 18748 10628 19073 10656
rect 18748 10616 18754 10628
rect 19061 10625 19073 10628
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 2038 10588 2044 10600
rect 1443 10560 2044 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 2038 10548 2044 10560
rect 2096 10548 2102 10600
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10588 9275 10591
rect 15933 10591 15991 10597
rect 9263 10560 10916 10588
rect 9263 10557 9275 10560
rect 9217 10551 9275 10557
rect 3145 10523 3203 10529
rect 3145 10489 3157 10523
rect 3191 10520 3203 10523
rect 9585 10523 9643 10529
rect 3191 10492 3740 10520
rect 3191 10489 3203 10492
rect 3145 10483 3203 10489
rect 3712 10464 3740 10492
rect 9585 10489 9597 10523
rect 9631 10520 9643 10523
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 9631 10492 10517 10520
rect 9631 10489 9643 10492
rect 9585 10483 9643 10489
rect 10505 10489 10517 10492
rect 10551 10520 10563 10523
rect 10778 10520 10784 10532
rect 10551 10492 10784 10520
rect 10551 10489 10563 10492
rect 10505 10483 10563 10489
rect 10778 10480 10784 10492
rect 10836 10480 10842 10532
rect 3418 10412 3424 10464
rect 3476 10452 3482 10464
rect 3605 10455 3663 10461
rect 3605 10452 3617 10455
rect 3476 10424 3617 10452
rect 3476 10412 3482 10424
rect 3605 10421 3617 10424
rect 3651 10421 3663 10455
rect 3605 10415 3663 10421
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 4341 10455 4399 10461
rect 3752 10424 3797 10452
rect 3752 10412 3758 10424
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 4430 10452 4436 10464
rect 4387 10424 4436 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 4614 10452 4620 10464
rect 4575 10424 4620 10452
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 5077 10455 5135 10461
rect 5077 10452 5089 10455
rect 4948 10424 5089 10452
rect 4948 10412 4954 10424
rect 5077 10421 5089 10424
rect 5123 10452 5135 10455
rect 7098 10452 7104 10464
rect 5123 10424 7104 10452
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10413 10455 10471 10461
rect 10413 10421 10425 10455
rect 10459 10452 10471 10455
rect 10888 10452 10916 10560
rect 15933 10557 15945 10591
rect 15979 10588 15991 10591
rect 16758 10588 16764 10600
rect 15979 10560 16764 10588
rect 15979 10557 15991 10560
rect 15933 10551 15991 10557
rect 16758 10548 16764 10560
rect 16816 10548 16822 10600
rect 17788 10588 17816 10616
rect 18322 10588 18328 10600
rect 17788 10560 18328 10588
rect 18322 10548 18328 10560
rect 18380 10588 18386 10600
rect 18509 10591 18567 10597
rect 18509 10588 18521 10591
rect 18380 10560 18521 10588
rect 18380 10548 18386 10560
rect 18509 10557 18521 10560
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 16301 10523 16359 10529
rect 16301 10489 16313 10523
rect 16347 10520 16359 10523
rect 17034 10520 17040 10532
rect 16347 10492 17040 10520
rect 16347 10489 16359 10492
rect 16301 10483 16359 10489
rect 17034 10480 17040 10492
rect 17092 10480 17098 10532
rect 11330 10452 11336 10464
rect 10459 10424 11336 10452
rect 10459 10421 10471 10424
rect 10413 10415 10471 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 16390 10452 16396 10464
rect 16351 10424 16396 10452
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 17402 10452 17408 10464
rect 17000 10424 17408 10452
rect 17000 10412 17006 10424
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 18414 10452 18420 10464
rect 18375 10424 18420 10452
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 3329 10251 3387 10257
rect 2832 10220 2877 10248
rect 2832 10208 2838 10220
rect 3329 10217 3341 10251
rect 3375 10248 3387 10251
rect 3418 10248 3424 10260
rect 3375 10220 3424 10248
rect 3375 10217 3387 10220
rect 3329 10211 3387 10217
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 4433 10251 4491 10257
rect 4433 10217 4445 10251
rect 4479 10248 4491 10251
rect 4522 10248 4528 10260
rect 4479 10220 4528 10248
rect 4479 10217 4491 10220
rect 4433 10211 4491 10217
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 6914 10248 6920 10260
rect 6875 10220 6920 10248
rect 6914 10208 6920 10220
rect 6972 10248 6978 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 6972 10220 7941 10248
rect 6972 10208 6978 10220
rect 7929 10217 7941 10220
rect 7975 10248 7987 10251
rect 8110 10248 8116 10260
rect 7975 10220 8116 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 10870 10208 10876 10260
rect 10928 10248 10934 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 10928 10220 11069 10248
rect 10928 10208 10934 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 11057 10211 11115 10217
rect 12989 10251 13047 10257
rect 12989 10217 13001 10251
rect 13035 10248 13047 10251
rect 13446 10248 13452 10260
rect 13035 10220 13452 10248
rect 13035 10217 13047 10220
rect 12989 10211 13047 10217
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14056 10220 14749 10248
rect 14056 10208 14062 10220
rect 14737 10217 14749 10220
rect 14783 10248 14795 10251
rect 14918 10248 14924 10260
rect 14783 10220 14924 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 16577 10251 16635 10257
rect 16577 10217 16589 10251
rect 16623 10248 16635 10251
rect 16850 10248 16856 10260
rect 16623 10220 16856 10248
rect 16623 10217 16635 10220
rect 16577 10211 16635 10217
rect 16850 10208 16856 10220
rect 16908 10248 16914 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 16908 10220 17693 10248
rect 16908 10208 16914 10220
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 18138 10248 18144 10260
rect 17681 10211 17739 10217
rect 17880 10220 18144 10248
rect 9858 10140 9864 10192
rect 9916 10189 9922 10192
rect 9916 10183 9980 10189
rect 9916 10149 9934 10183
rect 9968 10149 9980 10183
rect 9916 10143 9980 10149
rect 9916 10140 9922 10143
rect 17218 10140 17224 10192
rect 17276 10180 17282 10192
rect 17880 10180 17908 10220
rect 18138 10208 18144 10220
rect 18196 10248 18202 10260
rect 18690 10248 18696 10260
rect 18196 10220 18552 10248
rect 18651 10220 18696 10248
rect 18196 10208 18202 10220
rect 17276 10152 17908 10180
rect 18524 10180 18552 10220
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 26694 10248 26700 10260
rect 26655 10220 26700 10248
rect 26694 10208 26700 10220
rect 26752 10208 26758 10260
rect 21358 10180 21364 10192
rect 18524 10152 21364 10180
rect 17276 10140 17282 10152
rect 21358 10140 21364 10152
rect 21416 10140 21422 10192
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10112 4583 10115
rect 4798 10112 4804 10124
rect 4571 10084 4804 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10112 8171 10115
rect 8202 10112 8208 10124
rect 8159 10084 8208 10112
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 14918 10112 14924 10124
rect 14879 10084 14924 10112
rect 14918 10072 14924 10084
rect 14976 10072 14982 10124
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 15838 10112 15844 10124
rect 15712 10084 15844 10112
rect 15712 10072 15718 10084
rect 15838 10072 15844 10084
rect 15896 10112 15902 10124
rect 16485 10115 16543 10121
rect 16485 10112 16497 10115
rect 15896 10084 16497 10112
rect 15896 10072 15902 10084
rect 16485 10081 16497 10084
rect 16531 10081 16543 10115
rect 18046 10112 18052 10124
rect 18007 10084 18052 10112
rect 16485 10075 16543 10081
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 26510 10112 26516 10124
rect 26471 10084 26516 10112
rect 26510 10072 26516 10084
rect 26568 10072 26574 10124
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10044 4767 10047
rect 4890 10044 4896 10056
rect 4755 10016 4896 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 12158 10044 12164 10056
rect 12119 10016 12164 10044
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10044 16819 10047
rect 17034 10044 17040 10056
rect 16807 10016 17040 10044
rect 16807 10013 16819 10016
rect 16761 10007 16819 10013
rect 17034 10004 17040 10016
rect 17092 10004 17098 10056
rect 17310 10044 17316 10056
rect 17271 10016 17316 10044
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 17402 10004 17408 10056
rect 17460 10044 17466 10056
rect 18141 10047 18199 10053
rect 18141 10044 18153 10047
rect 17460 10016 18153 10044
rect 17460 10004 17466 10016
rect 18141 10013 18153 10016
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10044 18383 10047
rect 18690 10044 18696 10056
rect 18371 10016 18696 10044
rect 18371 10013 18383 10016
rect 18325 10007 18383 10013
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 2501 9979 2559 9985
rect 2501 9945 2513 9979
rect 2547 9976 2559 9979
rect 2866 9976 2872 9988
rect 2547 9948 2872 9976
rect 2547 9945 2559 9948
rect 2501 9939 2559 9945
rect 2866 9936 2872 9948
rect 2924 9976 2930 9988
rect 4065 9979 4123 9985
rect 4065 9976 4077 9979
rect 2924 9948 4077 9976
rect 2924 9936 2930 9948
rect 4065 9945 4077 9948
rect 4111 9945 4123 9979
rect 4065 9939 4123 9945
rect 2314 9868 2320 9920
rect 2372 9908 2378 9920
rect 2958 9908 2964 9920
rect 2372 9880 2964 9908
rect 2372 9868 2378 9880
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 16117 9911 16175 9917
rect 16117 9877 16129 9911
rect 16163 9908 16175 9911
rect 16482 9908 16488 9920
rect 16163 9880 16488 9908
rect 16163 9877 16175 9880
rect 16117 9871 16175 9877
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2409 9707 2467 9713
rect 2409 9704 2421 9707
rect 1452 9676 2421 9704
rect 1452 9664 1458 9676
rect 2409 9673 2421 9676
rect 2455 9704 2467 9707
rect 4246 9704 4252 9716
rect 2455 9676 4252 9704
rect 2455 9673 2467 9676
rect 2409 9667 2467 9673
rect 4246 9664 4252 9676
rect 4304 9664 4310 9716
rect 4522 9704 4528 9716
rect 4483 9676 4528 9704
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 4890 9704 4896 9716
rect 4851 9676 4896 9704
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 7156 9676 8217 9704
rect 7156 9664 7162 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 9674 9704 9680 9716
rect 8205 9667 8263 9673
rect 9600 9676 9680 9704
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 2041 9639 2099 9645
rect 2041 9605 2053 9639
rect 2087 9636 2099 9639
rect 3142 9636 3148 9648
rect 2087 9608 3148 9636
rect 2087 9605 2099 9608
rect 2041 9599 2099 9605
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 2056 9500 2084 9599
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 4157 9639 4215 9645
rect 4157 9605 4169 9639
rect 4203 9636 4215 9639
rect 4798 9636 4804 9648
rect 4203 9608 4804 9636
rect 4203 9605 4215 9608
rect 4157 9599 4215 9605
rect 4798 9596 4804 9608
rect 4856 9596 4862 9648
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 9309 9639 9367 9645
rect 9309 9636 9321 9639
rect 8168 9608 9321 9636
rect 8168 9596 8174 9608
rect 9309 9605 9321 9608
rect 9355 9636 9367 9639
rect 9600 9636 9628 9676
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 10778 9704 10784 9716
rect 10739 9676 10784 9704
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 11974 9704 11980 9716
rect 11572 9676 11980 9704
rect 11572 9664 11578 9676
rect 11974 9664 11980 9676
rect 12032 9664 12038 9716
rect 18690 9704 18696 9716
rect 15120 9676 16620 9704
rect 10594 9636 10600 9648
rect 9355 9608 9628 9636
rect 10555 9608 10600 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 12066 9636 12072 9648
rect 11256 9608 12072 9636
rect 6822 9568 6828 9580
rect 6783 9540 6828 9568
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 1443 9472 2084 9500
rect 10612 9500 10640 9596
rect 10870 9528 10876 9580
rect 10928 9568 10934 9580
rect 11256 9577 11284 9608
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 10928 9540 11253 9568
rect 10928 9528 10934 9540
rect 11241 9537 11253 9540
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 11425 9571 11483 9577
rect 11425 9537 11437 9571
rect 11471 9568 11483 9571
rect 11790 9568 11796 9580
rect 11471 9540 11796 9568
rect 11471 9537 11483 9540
rect 11425 9531 11483 9537
rect 11146 9500 11152 9512
rect 10612 9472 11152 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 7098 9441 7104 9444
rect 6641 9435 6699 9441
rect 6641 9401 6653 9435
rect 6687 9432 6699 9435
rect 7092 9432 7104 9441
rect 6687 9404 7104 9432
rect 6687 9401 6699 9404
rect 6641 9395 6699 9401
rect 7092 9395 7104 9404
rect 7098 9392 7104 9395
rect 7156 9392 7162 9444
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 9769 9435 9827 9441
rect 9769 9432 9781 9435
rect 9548 9404 9781 9432
rect 9548 9392 9554 9404
rect 9769 9401 9781 9404
rect 9815 9432 9827 9435
rect 9858 9432 9864 9444
rect 9815 9404 9864 9432
rect 9815 9401 9827 9404
rect 9769 9395 9827 9401
rect 9858 9392 9864 9404
rect 9916 9432 9922 9444
rect 10321 9435 10379 9441
rect 10321 9432 10333 9435
rect 9916 9404 10333 9432
rect 9916 9392 9922 9404
rect 10321 9401 10333 9404
rect 10367 9432 10379 9435
rect 11440 9432 11468 9531
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 13998 9568 14004 9580
rect 13959 9540 14004 9568
rect 13998 9528 14004 9540
rect 14056 9528 14062 9580
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9500 13967 9503
rect 14268 9503 14326 9509
rect 14268 9500 14280 9503
rect 13955 9472 14280 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 14268 9469 14280 9472
rect 14314 9500 14326 9503
rect 15120 9500 15148 9676
rect 16592 9509 16620 9676
rect 17880 9676 18696 9704
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 17880 9636 17908 9676
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 19794 9704 19800 9716
rect 19576 9676 19800 9704
rect 19576 9664 19582 9676
rect 19794 9664 19800 9676
rect 19852 9664 19858 9716
rect 17083 9608 17908 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 17954 9596 17960 9648
rect 18012 9596 18018 9648
rect 19429 9639 19487 9645
rect 19429 9636 19441 9639
rect 18524 9608 19441 9636
rect 14314 9472 15148 9500
rect 16577 9503 16635 9509
rect 14314 9469 14326 9472
rect 14268 9463 14326 9469
rect 16577 9469 16589 9503
rect 16623 9500 16635 9503
rect 17034 9500 17040 9512
rect 16623 9472 17040 9500
rect 16623 9469 16635 9472
rect 16577 9463 16635 9469
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 17310 9460 17316 9512
rect 17368 9500 17374 9512
rect 17681 9503 17739 9509
rect 17681 9500 17693 9503
rect 17368 9472 17693 9500
rect 17368 9460 17374 9472
rect 17681 9469 17693 9472
rect 17727 9469 17739 9503
rect 17681 9463 17739 9469
rect 17402 9432 17408 9444
rect 10367 9404 11468 9432
rect 15396 9404 17408 9432
rect 10367 9401 10379 9404
rect 10321 9395 10379 9401
rect 15396 9376 15424 9404
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 17972 9432 18000 9596
rect 18524 9580 18552 9608
rect 19429 9605 19441 9608
rect 19475 9605 19487 9639
rect 19429 9599 19487 9605
rect 18506 9568 18512 9580
rect 18467 9540 18512 9568
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 18690 9568 18696 9580
rect 18603 9540 18696 9568
rect 18690 9528 18696 9540
rect 18748 9568 18754 9580
rect 19061 9571 19119 9577
rect 19061 9568 19073 9571
rect 18748 9540 19073 9568
rect 18748 9528 18754 9540
rect 19061 9537 19073 9540
rect 19107 9537 19119 9571
rect 19061 9531 19119 9537
rect 18414 9500 18420 9512
rect 18375 9472 18420 9500
rect 18414 9460 18420 9472
rect 18472 9500 18478 9512
rect 19797 9503 19855 9509
rect 19797 9500 19809 9503
rect 18472 9472 19809 9500
rect 18472 9460 18478 9472
rect 19797 9469 19809 9472
rect 19843 9469 19855 9503
rect 26510 9500 26516 9512
rect 26471 9472 26516 9500
rect 19797 9463 19855 9469
rect 26510 9460 26516 9472
rect 26568 9460 26574 9512
rect 19150 9432 19156 9444
rect 17972 9404 19156 9432
rect 19150 9392 19156 9404
rect 19208 9392 19214 9444
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8754 9364 8760 9376
rect 8352 9336 8760 9364
rect 8352 9324 8358 9336
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 15378 9364 15384 9376
rect 15291 9336 15384 9364
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15838 9324 15844 9376
rect 15896 9364 15902 9376
rect 16209 9367 16267 9373
rect 16209 9364 16221 9367
rect 15896 9336 16221 9364
rect 15896 9324 15902 9336
rect 16209 9333 16221 9336
rect 16255 9364 16267 9367
rect 16482 9364 16488 9376
rect 16255 9336 16488 9364
rect 16255 9333 16267 9336
rect 16209 9327 16267 9333
rect 16482 9324 16488 9336
rect 16540 9324 16546 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 17218 9364 17224 9376
rect 16724 9336 17224 9364
rect 16724 9324 16730 9336
rect 17218 9324 17224 9336
rect 17276 9364 17282 9376
rect 17313 9367 17371 9373
rect 17313 9364 17325 9367
rect 17276 9336 17325 9364
rect 17276 9324 17282 9336
rect 17313 9333 17325 9336
rect 17359 9333 17371 9367
rect 18046 9364 18052 9376
rect 18007 9336 18052 9364
rect 17313 9327 17371 9333
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 3142 9160 3148 9172
rect 3103 9132 3148 9160
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 10870 9160 10876 9172
rect 10831 9132 10876 9160
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 11149 9163 11207 9169
rect 11149 9129 11161 9163
rect 11195 9160 11207 9163
rect 11330 9160 11336 9172
rect 11195 9132 11336 9160
rect 11195 9129 11207 9132
rect 11149 9123 11207 9129
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 11517 9163 11575 9169
rect 11517 9129 11529 9163
rect 11563 9160 11575 9163
rect 11606 9160 11612 9172
rect 11563 9132 11612 9160
rect 11563 9129 11575 9132
rect 11517 9123 11575 9129
rect 11606 9120 11612 9132
rect 11664 9160 11670 9172
rect 12158 9160 12164 9172
rect 11664 9132 12164 9160
rect 11664 9120 11670 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 13998 9160 14004 9172
rect 13959 9132 14004 9160
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 15657 9163 15715 9169
rect 15657 9129 15669 9163
rect 15703 9160 15715 9163
rect 16117 9163 16175 9169
rect 16117 9160 16129 9163
rect 15703 9132 16129 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 16117 9129 16129 9132
rect 16163 9160 16175 9163
rect 17313 9163 17371 9169
rect 17313 9160 17325 9163
rect 16163 9132 17325 9160
rect 16163 9129 16175 9132
rect 16117 9123 16175 9129
rect 17313 9129 17325 9132
rect 17359 9129 17371 9163
rect 17770 9160 17776 9172
rect 17683 9132 17776 9160
rect 17313 9123 17371 9129
rect 17770 9120 17776 9132
rect 17828 9160 17834 9172
rect 18877 9163 18935 9169
rect 18877 9160 18889 9163
rect 17828 9132 18889 9160
rect 17828 9120 17834 9132
rect 18877 9129 18889 9132
rect 18923 9129 18935 9163
rect 18877 9123 18935 9129
rect 18966 9120 18972 9172
rect 19024 9160 19030 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 19024 9132 19257 9160
rect 19024 9120 19030 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 26694 9160 26700 9172
rect 26655 9132 26700 9160
rect 19245 9123 19303 9129
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 6270 9092 6276 9104
rect 5736 9064 6276 9092
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 2498 9024 2504 9036
rect 2459 8996 2504 9024
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 5736 9033 5764 9064
rect 6270 9052 6276 9064
rect 6328 9092 6334 9104
rect 6822 9092 6828 9104
rect 6328 9064 6828 9092
rect 6328 9052 6334 9064
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 16206 9092 16212 9104
rect 16167 9064 16212 9092
rect 16206 9052 16212 9064
rect 16264 9052 16270 9104
rect 16850 9092 16856 9104
rect 16811 9064 16856 9092
rect 16850 9052 16856 9064
rect 16908 9052 16914 9104
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 19337 9095 19395 9101
rect 17092 9064 18644 9092
rect 17092 9052 17098 9064
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 5810 8984 5816 9036
rect 5868 9024 5874 9036
rect 5977 9027 6035 9033
rect 5977 9024 5989 9027
rect 5868 8996 5989 9024
rect 5868 8984 5874 8996
rect 5977 8993 5989 8996
rect 6023 8993 6035 9027
rect 5977 8987 6035 8993
rect 11514 8984 11520 9036
rect 11572 9024 11578 9036
rect 11609 9027 11667 9033
rect 11609 9024 11621 9027
rect 11572 8996 11621 9024
rect 11572 8984 11578 8996
rect 11609 8993 11621 8996
rect 11655 8993 11667 9027
rect 11609 8987 11667 8993
rect 17681 9027 17739 9033
rect 17681 8993 17693 9027
rect 17727 9024 17739 9027
rect 18506 9024 18512 9036
rect 17727 8996 18512 9024
rect 17727 8993 17739 8996
rect 17681 8987 17739 8993
rect 18506 8984 18512 8996
rect 18564 8984 18570 9036
rect 18616 9033 18644 9064
rect 19337 9061 19349 9095
rect 19383 9092 19395 9095
rect 19610 9092 19616 9104
rect 19383 9064 19616 9092
rect 19383 9061 19395 9064
rect 19337 9055 19395 9061
rect 19610 9052 19616 9064
rect 19668 9052 19674 9104
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 9024 18659 9027
rect 26510 9024 26516 9036
rect 18647 8996 19472 9024
rect 26471 8996 26516 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 19444 8968 19472 8996
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 11790 8956 11796 8968
rect 11751 8928 11796 8956
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 16356 8928 16401 8956
rect 16356 8916 16362 8928
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17460 8928 17969 8956
rect 17460 8916 17466 8928
rect 17957 8925 17969 8928
rect 18003 8956 18015 8959
rect 18690 8956 18696 8968
rect 18003 8928 18696 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 19484 8928 19529 8956
rect 19484 8916 19490 8928
rect 12250 8848 12256 8900
rect 12308 8888 12314 8900
rect 15749 8891 15807 8897
rect 15749 8888 15761 8891
rect 12308 8860 15761 8888
rect 12308 8848 12314 8860
rect 15749 8857 15761 8860
rect 15795 8857 15807 8891
rect 15749 8851 15807 8857
rect 2682 8820 2688 8832
rect 2643 8792 2688 8820
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 7098 8820 7104 8832
rect 7059 8792 7104 8820
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 8941 8823 8999 8829
rect 8941 8789 8953 8823
rect 8987 8820 8999 8823
rect 9490 8820 9496 8832
rect 8987 8792 9496 8820
rect 8987 8789 8999 8792
rect 8941 8783 8999 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 14737 8823 14795 8829
rect 14737 8820 14749 8823
rect 14424 8792 14749 8820
rect 14424 8780 14430 8792
rect 14737 8789 14749 8792
rect 14783 8820 14795 8823
rect 14918 8820 14924 8832
rect 14783 8792 14924 8820
rect 14783 8789 14795 8792
rect 14737 8783 14795 8789
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 18322 8820 18328 8832
rect 18012 8792 18328 8820
rect 18012 8780 18018 8792
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2498 8616 2504 8628
rect 2459 8588 2504 8616
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 5810 8616 5816 8628
rect 5723 8588 5816 8616
rect 5810 8576 5816 8588
rect 5868 8616 5874 8628
rect 7193 8619 7251 8625
rect 7193 8616 7205 8619
rect 5868 8588 7205 8616
rect 5868 8576 5874 8588
rect 7193 8585 7205 8588
rect 7239 8616 7251 8619
rect 7926 8616 7932 8628
rect 7239 8588 7932 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 11606 8616 11612 8628
rect 11567 8588 11612 8616
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 16482 8576 16488 8628
rect 16540 8616 16546 8628
rect 17126 8616 17132 8628
rect 16540 8588 17132 8616
rect 16540 8576 16546 8588
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 17402 8616 17408 8628
rect 17363 8588 17408 8616
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17770 8616 17776 8628
rect 17731 8588 17776 8616
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 18506 8616 18512 8628
rect 18467 8588 18512 8616
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 18966 8576 18972 8628
rect 19024 8616 19030 8628
rect 19521 8619 19579 8625
rect 19521 8616 19533 8619
rect 19024 8588 19533 8616
rect 19024 8576 19030 8588
rect 19521 8585 19533 8588
rect 19567 8616 19579 8619
rect 19886 8616 19892 8628
rect 19567 8588 19892 8616
rect 19567 8585 19579 8588
rect 19521 8579 19579 8585
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 26602 8616 26608 8628
rect 26563 8588 26608 8616
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 6181 8551 6239 8557
rect 6181 8517 6193 8551
rect 6227 8548 6239 8551
rect 6270 8548 6276 8560
rect 6227 8520 6276 8548
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 8849 8551 8907 8557
rect 8849 8548 8861 8551
rect 7668 8520 8861 8548
rect 2038 8480 2044 8492
rect 1412 8452 2044 8480
rect 1412 8421 1440 8452
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 3237 8483 3295 8489
rect 3237 8480 3249 8483
rect 3200 8452 3249 8480
rect 3200 8440 3206 8452
rect 3237 8449 3249 8452
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 3510 8480 3516 8492
rect 3467 8452 3516 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 7668 8424 7696 8520
rect 8849 8517 8861 8520
rect 8895 8517 8907 8551
rect 8849 8511 8907 8517
rect 11241 8551 11299 8557
rect 11241 8517 11253 8551
rect 11287 8548 11299 8551
rect 11514 8548 11520 8560
rect 11287 8520 11520 8548
rect 11287 8517 11299 8520
rect 11241 8511 11299 8517
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 13817 8551 13875 8557
rect 13817 8517 13829 8551
rect 13863 8548 13875 8551
rect 14366 8548 14372 8560
rect 13863 8520 14372 8548
rect 13863 8517 13875 8520
rect 13817 8511 13875 8517
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 17037 8551 17095 8557
rect 17037 8517 17049 8551
rect 17083 8548 17095 8551
rect 18524 8548 18552 8576
rect 19242 8548 19248 8560
rect 17083 8520 18552 8548
rect 18984 8520 19248 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 7926 8480 7932 8492
rect 7887 8452 7932 8480
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 9490 8480 9496 8492
rect 9451 8452 9496 8480
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8480 14795 8483
rect 18322 8480 18328 8492
rect 14783 8452 14964 8480
rect 18283 8452 18328 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 7650 8412 7656 8424
rect 7563 8384 7656 8412
rect 1397 8375 1455 8381
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8412 8815 8415
rect 9214 8412 9220 8424
rect 8803 8384 9220 8412
rect 8803 8381 8815 8384
rect 8757 8375 8815 8381
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8344 3203 8347
rect 3881 8347 3939 8353
rect 3881 8344 3893 8347
rect 3191 8316 3893 8344
rect 3191 8313 3203 8316
rect 3145 8307 3203 8313
rect 3881 8313 3893 8316
rect 3927 8344 3939 8347
rect 4341 8347 4399 8353
rect 4341 8344 4353 8347
rect 3927 8316 4353 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4341 8313 4353 8316
rect 4387 8313 4399 8347
rect 4341 8307 4399 8313
rect 6641 8347 6699 8353
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 7745 8347 7803 8353
rect 7745 8344 7757 8347
rect 6687 8316 7757 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 7745 8313 7757 8316
rect 7791 8344 7803 8347
rect 8389 8347 8447 8353
rect 7791 8316 8340 8344
rect 7791 8313 7803 8316
rect 7745 8307 7803 8313
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 7282 8276 7288 8288
rect 2832 8248 2877 8276
rect 7243 8248 7288 8276
rect 2832 8236 2838 8248
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 8312 8276 8340 8316
rect 8389 8313 8401 8347
rect 8435 8344 8447 8347
rect 9309 8347 9367 8353
rect 9309 8344 9321 8347
rect 8435 8316 9321 8344
rect 8435 8313 8447 8316
rect 8389 8307 8447 8313
rect 9309 8313 9321 8316
rect 9355 8344 9367 8347
rect 9582 8344 9588 8356
rect 9355 8316 9588 8344
rect 9355 8313 9367 8316
rect 9309 8307 9367 8313
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 14016 8344 14044 8375
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 14826 8412 14832 8424
rect 14148 8384 14832 8412
rect 14148 8372 14154 8384
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 14936 8412 14964 8452
rect 18322 8440 18328 8452
rect 18380 8480 18386 8492
rect 18984 8489 19012 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 26510 8508 26516 8560
rect 26568 8548 26574 8560
rect 27341 8551 27399 8557
rect 27341 8548 27353 8551
rect 26568 8520 27353 8548
rect 26568 8508 26574 8520
rect 27341 8517 27353 8520
rect 27387 8517 27399 8551
rect 27706 8548 27712 8560
rect 27667 8520 27712 8548
rect 27341 8511 27399 8517
rect 27706 8508 27712 8520
rect 27764 8508 27770 8560
rect 18969 8483 19027 8489
rect 18969 8480 18981 8483
rect 18380 8452 18981 8480
rect 18380 8440 18386 8452
rect 18969 8449 18981 8452
rect 19015 8449 19027 8483
rect 18969 8443 19027 8449
rect 19153 8483 19211 8489
rect 19153 8449 19165 8483
rect 19199 8480 19211 8483
rect 19426 8480 19432 8492
rect 19199 8452 19432 8480
rect 19199 8449 19211 8452
rect 19153 8443 19211 8449
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 15096 8415 15154 8421
rect 15096 8412 15108 8415
rect 14936 8384 15108 8412
rect 15096 8381 15108 8384
rect 15142 8412 15154 8415
rect 15378 8412 15384 8424
rect 15142 8384 15384 8412
rect 15142 8381 15154 8384
rect 15096 8375 15154 8381
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 26418 8412 26424 8424
rect 26379 8384 26424 8412
rect 26418 8372 26424 8384
rect 26476 8412 26482 8424
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26476 8384 26985 8412
rect 26476 8372 26482 8384
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 27522 8412 27528 8424
rect 27483 8384 27528 8412
rect 26973 8375 27031 8381
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27580 8384 28089 8412
rect 27580 8372 27586 8384
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 14277 8347 14335 8353
rect 14277 8344 14289 8347
rect 13740 8316 14289 8344
rect 8478 8276 8484 8288
rect 8312 8248 8484 8276
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 11977 8279 12035 8285
rect 11977 8276 11989 8279
rect 11848 8248 11989 8276
rect 11848 8236 11854 8248
rect 11977 8245 11989 8248
rect 12023 8276 12035 8279
rect 12526 8276 12532 8288
rect 12023 8248 12532 8276
rect 12023 8245 12035 8248
rect 11977 8239 12035 8245
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 13740 8276 13768 8316
rect 14277 8313 14289 8316
rect 14323 8313 14335 8347
rect 14277 8307 14335 8313
rect 17402 8304 17408 8356
rect 17460 8344 17466 8356
rect 19610 8344 19616 8356
rect 17460 8316 19616 8344
rect 17460 8304 17466 8316
rect 19610 8304 19616 8316
rect 19668 8344 19674 8356
rect 19889 8347 19947 8353
rect 19889 8344 19901 8347
rect 19668 8316 19901 8344
rect 19668 8304 19674 8316
rect 19889 8313 19901 8316
rect 19935 8313 19947 8347
rect 19889 8307 19947 8313
rect 12676 8248 13768 8276
rect 16209 8279 16267 8285
rect 12676 8236 12682 8248
rect 16209 8245 16221 8279
rect 16255 8276 16267 8279
rect 16298 8276 16304 8288
rect 16255 8248 16304 8276
rect 16255 8245 16267 8248
rect 16209 8239 16267 8245
rect 16298 8236 16304 8248
rect 16356 8276 16362 8288
rect 16574 8276 16580 8288
rect 16356 8248 16580 8276
rect 16356 8236 16362 8248
rect 16574 8236 16580 8248
rect 16632 8236 16638 8288
rect 18874 8276 18880 8288
rect 18835 8248 18880 8276
rect 18874 8236 18880 8248
rect 18932 8236 18938 8288
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 2317 8075 2375 8081
rect 2317 8041 2329 8075
rect 2363 8072 2375 8075
rect 2774 8072 2780 8084
rect 2363 8044 2780 8072
rect 2363 8041 2375 8044
rect 2317 8035 2375 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 3970 8072 3976 8084
rect 2924 8044 3976 8072
rect 2924 8032 2930 8044
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 7009 8075 7067 8081
rect 7009 8041 7021 8075
rect 7055 8072 7067 8075
rect 7282 8072 7288 8084
rect 7055 8044 7288 8072
rect 7055 8041 7067 8044
rect 7009 8035 7067 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7650 8072 7656 8084
rect 7611 8044 7656 8072
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 14093 8075 14151 8081
rect 14093 8041 14105 8075
rect 14139 8072 14151 8075
rect 14182 8072 14188 8084
rect 14139 8044 14188 8072
rect 14139 8041 14151 8044
rect 14093 8035 14151 8041
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 14826 8072 14832 8084
rect 14787 8044 14832 8072
rect 14826 8032 14832 8044
rect 14884 8032 14890 8084
rect 16209 8075 16267 8081
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 16390 8072 16396 8084
rect 16255 8044 16396 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 18601 8075 18659 8081
rect 18601 8041 18613 8075
rect 18647 8072 18659 8075
rect 18874 8072 18880 8084
rect 18647 8044 18880 8072
rect 18647 8041 18659 8044
rect 18601 8035 18659 8041
rect 18874 8032 18880 8044
rect 18932 8072 18938 8084
rect 18969 8075 19027 8081
rect 18969 8072 18981 8075
rect 18932 8044 18981 8072
rect 18932 8032 18938 8044
rect 18969 8041 18981 8044
rect 19015 8041 19027 8075
rect 19426 8072 19432 8084
rect 19387 8044 19432 8072
rect 18969 8035 19027 8041
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 26694 8072 26700 8084
rect 26655 8044 26700 8072
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 6917 8007 6975 8013
rect 6917 7973 6929 8007
rect 6963 8004 6975 8007
rect 7466 8004 7472 8016
rect 6963 7976 7472 8004
rect 6963 7973 6975 7976
rect 6917 7967 6975 7973
rect 7466 7964 7472 7976
rect 7524 7964 7530 8016
rect 2314 7896 2320 7948
rect 2372 7936 2378 7948
rect 2777 7939 2835 7945
rect 2777 7936 2789 7939
rect 2372 7908 2789 7936
rect 2372 7896 2378 7908
rect 2777 7905 2789 7908
rect 2823 7936 2835 7939
rect 3878 7936 3884 7948
rect 2823 7908 3884 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 9030 7936 9036 7948
rect 8991 7908 9036 7936
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 11698 7936 11704 7948
rect 11379 7908 11704 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 13998 7936 14004 7948
rect 13959 7908 14004 7936
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7936 15899 7939
rect 16574 7936 16580 7948
rect 15887 7908 16580 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 16574 7896 16580 7908
rect 16632 7936 16638 7948
rect 16741 7939 16799 7945
rect 16741 7936 16753 7939
rect 16632 7908 16753 7936
rect 16632 7896 16638 7908
rect 16741 7905 16753 7908
rect 16787 7905 16799 7939
rect 26510 7936 26516 7948
rect 26471 7908 26516 7936
rect 16741 7899 16799 7905
rect 26510 7896 26516 7908
rect 26568 7896 26574 7948
rect 1394 7828 1400 7880
rect 1452 7868 1458 7880
rect 1673 7871 1731 7877
rect 1673 7868 1685 7871
rect 1452 7840 1685 7868
rect 1452 7828 1458 7840
rect 1673 7837 1685 7840
rect 1719 7868 1731 7871
rect 2682 7868 2688 7880
rect 1719 7840 2688 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3099 7840 3556 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3528 7744 3556 7840
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 7098 7868 7104 7880
rect 6696 7840 7104 7868
rect 6696 7828 6702 7840
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 13464 7840 14197 7868
rect 12618 7800 12624 7812
rect 12579 7772 12624 7800
rect 12618 7760 12624 7772
rect 12676 7760 12682 7812
rect 13464 7744 13492 7840
rect 14185 7837 14197 7840
rect 14231 7837 14243 7871
rect 14185 7831 14243 7837
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 16482 7868 16488 7880
rect 14884 7840 16488 7868
rect 14884 7828 14890 7840
rect 16482 7828 16488 7840
rect 16540 7828 16546 7880
rect 2406 7732 2412 7744
rect 2367 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 3510 7732 3516 7744
rect 3471 7704 3516 7732
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 4338 7732 4344 7744
rect 4299 7704 4344 7732
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 6546 7732 6552 7744
rect 6507 7704 6552 7732
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8754 7732 8760 7744
rect 8352 7704 8760 7732
rect 8352 7692 8358 7704
rect 8754 7692 8760 7704
rect 8812 7732 8818 7744
rect 8849 7735 8907 7741
rect 8849 7732 8861 7735
rect 8812 7704 8861 7732
rect 8812 7692 8818 7704
rect 8849 7701 8861 7704
rect 8895 7701 8907 7735
rect 8849 7695 8907 7701
rect 10781 7735 10839 7741
rect 10781 7701 10793 7735
rect 10827 7732 10839 7735
rect 11422 7732 11428 7744
rect 10827 7704 11428 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 11422 7692 11428 7704
rect 11480 7692 11486 7744
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13630 7732 13636 7744
rect 13591 7704 13636 7732
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 17862 7732 17868 7744
rect 17823 7704 17868 7732
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 2314 7528 2320 7540
rect 2275 7500 2320 7528
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 5629 7531 5687 7537
rect 5629 7528 5641 7531
rect 3068 7500 5641 7528
rect 3068 7404 3096 7500
rect 5629 7497 5641 7500
rect 5675 7528 5687 7531
rect 5718 7528 5724 7540
rect 5675 7500 5724 7528
rect 5675 7497 5687 7500
rect 5629 7491 5687 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 6638 7528 6644 7540
rect 6599 7500 6644 7528
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7528 7159 7531
rect 7282 7528 7288 7540
rect 7147 7500 7288 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 7466 7528 7472 7540
rect 7427 7500 7472 7528
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 9030 7528 9036 7540
rect 8343 7500 9036 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 10192 7500 10517 7528
rect 10192 7488 10198 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 10505 7491 10563 7497
rect 8478 7420 8484 7472
rect 8536 7460 8542 7472
rect 9125 7463 9183 7469
rect 9125 7460 9137 7463
rect 8536 7432 9137 7460
rect 8536 7420 8542 7432
rect 9125 7429 9137 7432
rect 9171 7429 9183 7463
rect 9125 7423 9183 7429
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7392 2007 7395
rect 2866 7392 2872 7404
rect 1995 7364 2872 7392
rect 1995 7361 2007 7364
rect 1949 7355 2007 7361
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 3050 7392 3056 7404
rect 3011 7364 3056 7392
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9490 7392 9496 7404
rect 9079 7364 9496 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 9490 7352 9496 7364
rect 9548 7392 9554 7404
rect 9677 7395 9735 7401
rect 9677 7392 9689 7395
rect 9548 7364 9689 7392
rect 9548 7352 9554 7364
rect 9677 7361 9689 7364
rect 9723 7361 9735 7395
rect 10520 7392 10548 7491
rect 14182 7488 14188 7540
rect 14240 7528 14246 7540
rect 14277 7531 14335 7537
rect 14277 7528 14289 7531
rect 14240 7500 14289 7528
rect 14240 7488 14246 7500
rect 14277 7497 14289 7500
rect 14323 7497 14335 7531
rect 16574 7528 16580 7540
rect 16535 7500 16580 7528
rect 14277 7491 14335 7497
rect 16574 7488 16580 7500
rect 16632 7488 16638 7540
rect 19334 7488 19340 7540
rect 19392 7528 19398 7540
rect 20162 7528 20168 7540
rect 19392 7500 20168 7528
rect 19392 7488 19398 7500
rect 20162 7488 20168 7500
rect 20220 7488 20226 7540
rect 22094 7488 22100 7540
rect 22152 7528 22158 7540
rect 23198 7528 23204 7540
rect 22152 7500 23204 7528
rect 22152 7488 22158 7500
rect 23198 7488 23204 7500
rect 23256 7488 23262 7540
rect 26510 7488 26516 7540
rect 26568 7528 26574 7540
rect 27341 7531 27399 7537
rect 27341 7528 27353 7531
rect 26568 7500 27353 7528
rect 26568 7488 26574 7500
rect 27341 7497 27353 7500
rect 27387 7497 27399 7531
rect 27341 7491 27399 7497
rect 16482 7420 16488 7472
rect 16540 7460 16546 7472
rect 16853 7463 16911 7469
rect 16853 7460 16865 7463
rect 16540 7432 16865 7460
rect 16540 7420 16546 7432
rect 16853 7429 16865 7432
rect 16899 7429 16911 7463
rect 16853 7423 16911 7429
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 10520 7364 11161 7392
rect 9677 7355 9735 7361
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 11333 7395 11391 7401
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 11422 7392 11428 7404
rect 11379 7364 11428 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 2774 7284 2780 7336
rect 2832 7324 2838 7336
rect 4249 7327 4307 7333
rect 2832 7296 2877 7324
rect 2832 7284 2838 7296
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 4338 7324 4344 7336
rect 4295 7296 4344 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 4338 7284 4344 7296
rect 4396 7284 4402 7336
rect 11164 7324 11192 7355
rect 11422 7352 11428 7364
rect 11480 7352 11486 7404
rect 12802 7392 12808 7404
rect 12715 7364 12808 7392
rect 12802 7352 12808 7364
rect 12860 7392 12866 7404
rect 13722 7392 13728 7404
rect 12860 7364 13728 7392
rect 12860 7352 12866 7364
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 11882 7324 11888 7336
rect 11164 7296 11888 7324
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 13924 7324 13952 7355
rect 13504 7296 13952 7324
rect 13504 7284 13510 7296
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 2869 7259 2927 7265
rect 2869 7256 2881 7259
rect 2372 7228 2881 7256
rect 2372 7216 2378 7228
rect 2869 7225 2881 7228
rect 2915 7225 2927 7259
rect 3510 7256 3516 7268
rect 3423 7228 3516 7256
rect 2869 7219 2927 7225
rect 3510 7216 3516 7228
rect 3568 7256 3574 7268
rect 4157 7259 4215 7265
rect 4157 7256 4169 7259
rect 3568 7228 4169 7256
rect 3568 7216 3574 7228
rect 4157 7225 4169 7228
rect 4203 7256 4215 7259
rect 4516 7259 4574 7265
rect 4516 7256 4528 7259
rect 4203 7228 4528 7256
rect 4203 7225 4215 7228
rect 4157 7219 4215 7225
rect 4516 7225 4528 7228
rect 4562 7256 4574 7259
rect 4706 7256 4712 7268
rect 4562 7228 4712 7256
rect 4562 7225 4574 7228
rect 4516 7219 4574 7225
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 8665 7259 8723 7265
rect 8665 7225 8677 7259
rect 8711 7256 8723 7259
rect 9493 7259 9551 7265
rect 9493 7256 9505 7259
rect 8711 7228 9505 7256
rect 8711 7225 8723 7228
rect 8665 7219 8723 7225
rect 9493 7225 9505 7228
rect 9539 7256 9551 7259
rect 11698 7256 11704 7268
rect 9539 7228 10732 7256
rect 11659 7228 11704 7256
rect 9539 7225 9551 7228
rect 9493 7219 9551 7225
rect 2406 7188 2412 7200
rect 2367 7160 2412 7188
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 9214 7148 9220 7200
rect 9272 7188 9278 7200
rect 10704 7197 10732 7228
rect 11698 7216 11704 7228
rect 11756 7216 11762 7268
rect 13081 7259 13139 7265
rect 13081 7225 13093 7259
rect 13127 7256 13139 7259
rect 13538 7256 13544 7268
rect 13127 7228 13544 7256
rect 13127 7225 13139 7228
rect 13081 7219 13139 7225
rect 13538 7216 13544 7228
rect 13596 7256 13602 7268
rect 13633 7259 13691 7265
rect 13633 7256 13645 7259
rect 13596 7228 13645 7256
rect 13596 7216 13602 7228
rect 13633 7225 13645 7228
rect 13679 7225 13691 7259
rect 13633 7219 13691 7225
rect 9585 7191 9643 7197
rect 9585 7188 9597 7191
rect 9272 7160 9597 7188
rect 9272 7148 9278 7160
rect 9585 7157 9597 7160
rect 9631 7157 9643 7191
rect 9585 7151 9643 7157
rect 10689 7191 10747 7197
rect 10689 7157 10701 7191
rect 10735 7157 10747 7191
rect 10689 7151 10747 7157
rect 10778 7148 10784 7200
rect 10836 7188 10842 7200
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 10836 7160 11069 7188
rect 10836 7148 10842 7160
rect 11057 7157 11069 7160
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 12986 7148 12992 7200
rect 13044 7188 13050 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 13044 7160 13277 7188
rect 13044 7148 13050 7160
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13265 7151 13323 7157
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 13924 7188 13952 7296
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 26421 7327 26479 7333
rect 26421 7324 26433 7327
rect 18932 7296 26433 7324
rect 18932 7284 18938 7296
rect 26421 7293 26433 7296
rect 26467 7324 26479 7327
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26467 7296 26985 7324
rect 26467 7293 26479 7296
rect 26421 7287 26479 7293
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 26973 7287 27031 7293
rect 13998 7216 14004 7268
rect 14056 7256 14062 7268
rect 14829 7259 14887 7265
rect 14829 7256 14841 7259
rect 14056 7228 14841 7256
rect 14056 7216 14062 7228
rect 14829 7225 14841 7228
rect 14875 7225 14887 7259
rect 14829 7219 14887 7225
rect 14737 7191 14795 7197
rect 14737 7188 14749 7191
rect 13780 7160 14749 7188
rect 13780 7148 13786 7160
rect 14737 7157 14749 7160
rect 14783 7188 14795 7191
rect 15102 7188 15108 7200
rect 14783 7160 15108 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 26602 7188 26608 7200
rect 26563 7160 26608 7188
rect 26602 7148 26608 7160
rect 26660 7148 26666 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 2041 6987 2099 6993
rect 2041 6953 2053 6987
rect 2087 6984 2099 6987
rect 2406 6984 2412 6996
rect 2087 6956 2412 6984
rect 2087 6953 2099 6956
rect 2041 6947 2099 6953
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 13265 6987 13323 6993
rect 13265 6984 13277 6987
rect 12400 6956 13277 6984
rect 12400 6944 12406 6956
rect 13265 6953 13277 6956
rect 13311 6984 13323 6987
rect 13630 6984 13636 6996
rect 13311 6956 13636 6984
rect 13311 6953 13323 6956
rect 13265 6947 13323 6953
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 13998 6984 14004 6996
rect 13959 6956 14004 6984
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 2314 6916 2320 6928
rect 2275 6888 2320 6916
rect 2314 6876 2320 6888
rect 2372 6876 2378 6928
rect 4338 6876 4344 6928
rect 4396 6916 4402 6928
rect 4396 6888 5580 6916
rect 4396 6876 4402 6888
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1670 6848 1676 6860
rect 1443 6820 1676 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6848 2559 6851
rect 2682 6848 2688 6860
rect 2547 6820 2688 6848
rect 2547 6817 2559 6820
rect 2501 6811 2559 6817
rect 2682 6808 2688 6820
rect 2740 6848 2746 6860
rect 3786 6848 3792 6860
rect 2740 6820 3792 6848
rect 2740 6808 2746 6820
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4614 6848 4620 6860
rect 4111 6820 4620 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 5552 6848 5580 6888
rect 5718 6876 5724 6928
rect 5776 6916 5782 6928
rect 5966 6919 6024 6925
rect 5966 6916 5978 6919
rect 5776 6888 5978 6916
rect 5776 6876 5782 6888
rect 5966 6885 5978 6888
rect 6012 6885 6024 6919
rect 5966 6879 6024 6885
rect 17862 6876 17868 6928
rect 17920 6876 17926 6928
rect 6270 6848 6276 6860
rect 5552 6820 6276 6848
rect 5736 6789 5764 6820
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 8389 6851 8447 6857
rect 8389 6848 8401 6851
rect 8352 6820 8401 6848
rect 8352 6808 8358 6820
rect 8389 6817 8401 6820
rect 8435 6817 8447 6851
rect 8389 6811 8447 6817
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6848 10103 6851
rect 10226 6848 10232 6860
rect 10091 6820 10232 6848
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 11422 6857 11428 6860
rect 11405 6851 11428 6857
rect 11405 6848 11417 6851
rect 10336 6820 11417 6848
rect 10336 6792 10364 6820
rect 11405 6817 11417 6820
rect 11480 6848 11486 6860
rect 11480 6820 11553 6848
rect 11405 6811 11428 6817
rect 11422 6808 11428 6811
rect 11480 6808 11486 6820
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 13044 6820 13369 6848
rect 13044 6808 13050 6820
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 17880 6848 17908 6876
rect 18138 6857 18144 6860
rect 18132 6848 18144 6857
rect 17880 6820 18144 6848
rect 13357 6811 13415 6817
rect 18132 6811 18144 6820
rect 18138 6808 18144 6811
rect 18196 6808 18202 6860
rect 26510 6848 26516 6860
rect 26471 6820 26516 6848
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9364 6752 10149 6780
rect 9364 6740 9370 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10137 6743 10195 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 10686 6780 10692 6792
rect 10647 6752 10692 6780
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6749 11207 6783
rect 13446 6780 13452 6792
rect 13407 6752 13452 6780
rect 11149 6743 11207 6749
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2648 6684 2697 6712
rect 2648 6672 2654 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 4246 6712 4252 6724
rect 4207 6684 4252 6712
rect 2685 6675 2743 6681
rect 4246 6672 4252 6684
rect 4304 6672 4310 6724
rect 9674 6712 9680 6724
rect 9635 6684 9680 6712
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 3050 6644 3056 6656
rect 3011 6616 3056 6644
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 7101 6647 7159 6653
rect 7101 6613 7113 6647
rect 7147 6644 7159 6647
rect 7190 6644 7196 6656
rect 7147 6616 7196 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 8205 6647 8263 6653
rect 8205 6644 8217 6647
rect 7432 6616 8217 6644
rect 7432 6604 7438 6616
rect 8205 6613 8217 6616
rect 8251 6613 8263 6647
rect 9214 6644 9220 6656
rect 9175 6616 9220 6644
rect 8205 6607 8263 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 11164 6644 11192 6743
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 17862 6780 17868 6792
rect 17823 6752 17868 6780
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 12526 6712 12532 6724
rect 12487 6684 12532 6712
rect 12526 6672 12532 6684
rect 12584 6672 12590 6724
rect 26694 6712 26700 6724
rect 26655 6684 26700 6712
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 11514 6644 11520 6656
rect 11164 6616 11520 6644
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 12894 6644 12900 6656
rect 12855 6616 12900 6644
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 16025 6647 16083 6653
rect 16025 6644 16037 6647
rect 15252 6616 16037 6644
rect 15252 6604 15258 6616
rect 16025 6613 16037 6616
rect 16071 6644 16083 6647
rect 16482 6644 16488 6656
rect 16071 6616 16488 6644
rect 16071 6613 16083 6616
rect 16025 6607 16083 6613
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 19242 6644 19248 6656
rect 19203 6616 19248 6644
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1670 6440 1676 6452
rect 1631 6412 1676 6440
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 3053 6443 3111 6449
rect 3053 6440 3065 6443
rect 2740 6412 3065 6440
rect 2740 6400 2746 6412
rect 3053 6409 3065 6412
rect 3099 6409 3111 6443
rect 3053 6403 3111 6409
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 4157 6443 4215 6449
rect 4157 6440 4169 6443
rect 4028 6412 4169 6440
rect 4028 6400 4034 6412
rect 4157 6409 4169 6412
rect 4203 6409 4215 6443
rect 5718 6440 5724 6452
rect 5679 6412 5724 6440
rect 4157 6403 4215 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 9272 6412 9873 6440
rect 9272 6400 9278 6412
rect 9861 6409 9873 6412
rect 9907 6409 9919 6443
rect 9861 6403 9919 6409
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12342 6440 12348 6452
rect 12299 6412 12348 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 15746 6440 15752 6452
rect 15707 6412 15752 6440
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 18601 6443 18659 6449
rect 18601 6440 18613 6443
rect 17920 6412 18613 6440
rect 17920 6400 17926 6412
rect 18601 6409 18613 6412
rect 18647 6409 18659 6443
rect 18601 6403 18659 6409
rect 3786 6372 3792 6384
rect 3747 6344 3792 6372
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 4614 6372 4620 6384
rect 4575 6344 4620 6372
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 8757 6375 8815 6381
rect 8757 6341 8769 6375
rect 8803 6372 8815 6375
rect 10318 6372 10324 6384
rect 8803 6344 10324 6372
rect 8803 6341 8815 6344
rect 8757 6335 8815 6341
rect 10318 6332 10324 6344
rect 10376 6372 10382 6384
rect 10376 6344 10456 6372
rect 10376 6332 10382 6344
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2593 6307 2651 6313
rect 2593 6304 2605 6307
rect 2188 6276 2605 6304
rect 2188 6264 2194 6276
rect 2593 6273 2605 6276
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6304 9827 6307
rect 9858 6304 9864 6316
rect 9815 6276 9864 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 9858 6264 9864 6276
rect 9916 6304 9922 6316
rect 10428 6313 10456 6344
rect 10413 6307 10471 6313
rect 9916 6276 10364 6304
rect 9916 6264 9922 6276
rect 2406 6236 2412 6248
rect 2367 6208 2412 6236
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6205 2559 6239
rect 2501 6199 2559 6205
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6236 3663 6239
rect 3970 6236 3976 6248
rect 3651 6208 3976 6236
rect 3651 6205 3663 6208
rect 3605 6199 3663 6205
rect 2516 6168 2544 6199
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 7190 6236 7196 6248
rect 7151 6208 7196 6236
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 10336 6245 10364 6276
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10459 6276 10885 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10873 6273 10885 6276
rect 10919 6304 10931 6307
rect 11241 6307 11299 6313
rect 11241 6304 11253 6307
rect 10919 6276 11253 6304
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 11241 6273 11253 6276
rect 11287 6273 11299 6307
rect 11241 6267 11299 6273
rect 13357 6307 13415 6313
rect 13357 6273 13369 6307
rect 13403 6304 13415 6307
rect 13403 6276 13584 6304
rect 13403 6273 13415 6276
rect 13357 6267 13415 6273
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 11330 6236 11336 6248
rect 10367 6208 11336 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 11330 6196 11336 6208
rect 11388 6196 11394 6248
rect 13449 6239 13507 6245
rect 13449 6205 13461 6239
rect 13495 6205 13507 6239
rect 13556 6236 13584 6276
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 16482 6304 16488 6316
rect 16264 6276 16488 6304
rect 16264 6264 16270 6276
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 13722 6245 13728 6248
rect 13716 6236 13728 6245
rect 13556 6208 13728 6236
rect 13449 6199 13507 6205
rect 13716 6199 13728 6208
rect 3421 6171 3479 6177
rect 3421 6168 3433 6171
rect 2424 6140 3433 6168
rect 2424 6112 2452 6140
rect 3421 6137 3433 6140
rect 3467 6137 3479 6171
rect 7208 6168 7236 6196
rect 7622 6171 7680 6177
rect 7622 6168 7634 6171
rect 7208 6140 7634 6168
rect 3421 6131 3479 6137
rect 7622 6137 7634 6140
rect 7668 6137 7680 6171
rect 7622 6131 7680 6137
rect 12989 6171 13047 6177
rect 12989 6137 13001 6171
rect 13035 6168 13047 6171
rect 13464 6168 13492 6199
rect 13722 6196 13728 6199
rect 13780 6196 13786 6248
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 16301 6239 16359 6245
rect 16301 6236 16313 6239
rect 15804 6208 16313 6236
rect 15804 6196 15810 6208
rect 16301 6205 16313 6208
rect 16347 6205 16359 6239
rect 26510 6236 26516 6248
rect 26471 6208 26516 6236
rect 16301 6199 16359 6205
rect 26510 6196 26516 6208
rect 26568 6196 26574 6248
rect 13538 6168 13544 6180
rect 13035 6140 13400 6168
rect 13464 6140 13544 6168
rect 13035 6137 13047 6140
rect 12989 6131 13047 6137
rect 13372 6112 13400 6140
rect 13538 6128 13544 6140
rect 13596 6128 13602 6180
rect 15473 6171 15531 6177
rect 15473 6137 15485 6171
rect 15519 6168 15531 6171
rect 16390 6168 16396 6180
rect 15519 6140 16396 6168
rect 15519 6137 15531 6140
rect 15473 6131 15531 6137
rect 16390 6128 16396 6140
rect 16448 6128 16454 6180
rect 1486 6060 1492 6112
rect 1544 6100 1550 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 1544 6072 2053 6100
rect 1544 6060 1550 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2041 6063 2099 6069
rect 2406 6060 2412 6112
rect 2464 6060 2470 6112
rect 6181 6103 6239 6109
rect 6181 6069 6193 6103
rect 6227 6100 6239 6103
rect 6270 6100 6276 6112
rect 6227 6072 6276 6100
rect 6227 6069 6239 6072
rect 6181 6063 6239 6069
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 9306 6100 9312 6112
rect 9267 6072 9312 6100
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 10192 6072 10241 6100
rect 10192 6060 10198 6072
rect 10229 6069 10241 6072
rect 10275 6100 10287 6103
rect 10410 6100 10416 6112
rect 10275 6072 10416 6100
rect 10275 6069 10287 6072
rect 10229 6063 10287 6069
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 11609 6103 11667 6109
rect 11609 6100 11621 6103
rect 11572 6072 11621 6100
rect 11572 6060 11578 6072
rect 11609 6069 11621 6072
rect 11655 6069 11667 6103
rect 11609 6063 11667 6069
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 13412 6072 14841 6100
rect 13412 6060 13418 6072
rect 14829 6069 14841 6072
rect 14875 6100 14887 6103
rect 15102 6100 15108 6112
rect 14875 6072 15108 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 15102 6060 15108 6072
rect 15160 6060 15166 6112
rect 15838 6060 15844 6112
rect 15896 6100 15902 6112
rect 15933 6103 15991 6109
rect 15933 6100 15945 6103
rect 15896 6072 15945 6100
rect 15896 6060 15902 6072
rect 15933 6069 15945 6072
rect 15979 6069 15991 6103
rect 18230 6100 18236 6112
rect 18191 6072 18236 6100
rect 15933 6063 15991 6069
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 2130 5896 2136 5908
rect 2091 5868 2136 5896
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 2406 5896 2412 5908
rect 2367 5868 2412 5896
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 2832 5868 4077 5896
rect 2832 5856 2838 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 4065 5859 4123 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 10318 5856 10324 5908
rect 10376 5896 10382 5908
rect 10597 5899 10655 5905
rect 10597 5896 10609 5899
rect 10376 5868 10609 5896
rect 10376 5856 10382 5868
rect 10597 5865 10609 5868
rect 10643 5865 10655 5899
rect 12986 5896 12992 5908
rect 12947 5868 12992 5896
rect 10597 5859 10655 5865
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13538 5896 13544 5908
rect 13451 5868 13544 5896
rect 13538 5856 13544 5868
rect 13596 5896 13602 5908
rect 14274 5896 14280 5908
rect 13596 5868 14280 5896
rect 13596 5856 13602 5868
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 15657 5899 15715 5905
rect 15657 5865 15669 5899
rect 15703 5896 15715 5899
rect 16209 5899 16267 5905
rect 16209 5896 16221 5899
rect 15703 5868 16221 5896
rect 15703 5865 15715 5868
rect 15657 5859 15715 5865
rect 16209 5865 16221 5868
rect 16255 5896 16267 5899
rect 17313 5899 17371 5905
rect 17313 5896 17325 5899
rect 16255 5868 17325 5896
rect 16255 5865 16267 5868
rect 16209 5859 16267 5865
rect 17313 5865 17325 5868
rect 17359 5865 17371 5899
rect 17678 5896 17684 5908
rect 17639 5868 17684 5896
rect 17313 5859 17371 5865
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 26694 5896 26700 5908
rect 26655 5868 26700 5896
rect 26694 5856 26700 5868
rect 26752 5856 26758 5908
rect 9953 5831 10011 5837
rect 9953 5797 9965 5831
rect 9999 5828 10011 5831
rect 10134 5828 10140 5840
rect 9999 5800 10140 5828
rect 9999 5797 10011 5800
rect 9953 5791 10011 5797
rect 10134 5788 10140 5800
rect 10192 5828 10198 5840
rect 17696 5828 17724 5856
rect 10192 5800 17724 5828
rect 10192 5788 10198 5800
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 3660 5732 4445 5760
rect 3660 5720 3666 5732
rect 4433 5729 4445 5732
rect 4479 5760 4491 5763
rect 4982 5760 4988 5772
rect 4479 5732 4988 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 14366 5720 14372 5772
rect 14424 5760 14430 5772
rect 14461 5763 14519 5769
rect 14461 5760 14473 5763
rect 14424 5732 14473 5760
rect 14424 5720 14430 5732
rect 14461 5729 14473 5732
rect 14507 5729 14519 5763
rect 14461 5723 14519 5729
rect 16117 5763 16175 5769
rect 16117 5729 16129 5763
rect 16163 5760 16175 5763
rect 16482 5760 16488 5772
rect 16163 5732 16488 5760
rect 16163 5729 16175 5732
rect 16117 5723 16175 5729
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 26510 5760 26516 5772
rect 26471 5732 26516 5760
rect 26510 5720 26516 5732
rect 26568 5720 26574 5772
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3050 5692 3056 5704
rect 3011 5664 3056 5692
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3878 5692 3884 5704
rect 3791 5664 3884 5692
rect 3878 5652 3884 5664
rect 3936 5692 3942 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 3936 5664 4537 5692
rect 3936 5652 3942 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4525 5655 4583 5661
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 15562 5652 15568 5704
rect 15620 5692 15626 5704
rect 16206 5692 16212 5704
rect 15620 5664 16212 5692
rect 15620 5652 15626 5664
rect 16206 5652 16212 5664
rect 16264 5692 16270 5704
rect 16301 5695 16359 5701
rect 16301 5692 16313 5695
rect 16264 5664 16313 5692
rect 16264 5652 16270 5664
rect 16301 5661 16313 5664
rect 16347 5661 16359 5695
rect 16301 5655 16359 5661
rect 17494 5652 17500 5704
rect 17552 5692 17558 5704
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 17552 5664 17785 5692
rect 17552 5652 17558 5664
rect 17773 5661 17785 5664
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5692 17923 5695
rect 18230 5692 18236 5704
rect 17911 5664 18236 5692
rect 17911 5661 17923 5664
rect 17865 5655 17923 5661
rect 15286 5584 15292 5636
rect 15344 5624 15350 5636
rect 16666 5624 16672 5636
rect 15344 5596 16672 5624
rect 15344 5584 15350 5596
rect 16666 5584 16672 5596
rect 16724 5584 16730 5636
rect 17678 5584 17684 5636
rect 17736 5624 17742 5636
rect 17880 5624 17908 5655
rect 18230 5652 18236 5664
rect 18288 5692 18294 5704
rect 18325 5695 18383 5701
rect 18325 5692 18337 5695
rect 18288 5664 18337 5692
rect 18288 5652 18294 5664
rect 18325 5661 18337 5664
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 17736 5596 17908 5624
rect 17736 5584 17742 5596
rect 6270 5516 6276 5568
rect 6328 5556 6334 5568
rect 7374 5556 7380 5568
rect 6328 5528 7380 5556
rect 6328 5516 6334 5528
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 10226 5556 10232 5568
rect 10187 5528 10232 5556
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 15746 5556 15752 5568
rect 15707 5528 15752 5556
rect 15746 5516 15752 5528
rect 15804 5516 15810 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 2038 5352 2044 5364
rect 1999 5324 2044 5352
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 3878 5352 3884 5364
rect 3839 5324 3884 5352
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 4982 5352 4988 5364
rect 4943 5324 4988 5352
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 13265 5355 13323 5361
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13354 5352 13360 5364
rect 13311 5324 13360 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 15562 5352 15568 5364
rect 15523 5324 15568 5352
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 16390 5352 16396 5364
rect 16351 5324 16396 5352
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 18046 5352 18052 5364
rect 18007 5324 18052 5352
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 25866 5312 25872 5364
rect 25924 5352 25930 5364
rect 26237 5355 26295 5361
rect 26237 5352 26249 5355
rect 25924 5324 26249 5352
rect 25924 5312 25930 5324
rect 26237 5321 26249 5324
rect 26283 5321 26295 5355
rect 26602 5352 26608 5364
rect 26563 5324 26608 5352
rect 26237 5315 26295 5321
rect 1394 5244 1400 5296
rect 1452 5284 1458 5296
rect 1578 5284 1584 5296
rect 1452 5256 1584 5284
rect 1452 5244 1458 5256
rect 1578 5244 1584 5256
rect 1636 5244 1642 5296
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 13372 5216 13400 5312
rect 15933 5219 15991 5225
rect 4571 5188 5396 5216
rect 13372 5188 13492 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 2038 5148 2044 5160
rect 1443 5120 2044 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 2498 5148 2504 5160
rect 2455 5120 2504 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 2498 5108 2504 5120
rect 2556 5108 2562 5160
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 3421 5151 3479 5157
rect 3421 5148 3433 5151
rect 2832 5120 3433 5148
rect 2832 5108 2838 5120
rect 3421 5117 3433 5120
rect 3467 5148 3479 5151
rect 4246 5148 4252 5160
rect 3467 5120 4252 5148
rect 3467 5117 3479 5120
rect 3421 5111 3479 5117
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 5368 5089 5396 5188
rect 13354 5148 13360 5160
rect 13315 5120 13360 5148
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 13464 5148 13492 5188
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 15979 5188 16957 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16945 5185 16957 5188
rect 16991 5216 17003 5219
rect 17678 5216 17684 5228
rect 16991 5188 17684 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17678 5176 17684 5188
rect 17736 5216 17742 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 17736 5188 18613 5216
rect 17736 5176 17742 5188
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 13613 5151 13671 5157
rect 13613 5148 13625 5151
rect 13464 5120 13625 5148
rect 13613 5117 13625 5120
rect 13659 5117 13671 5151
rect 16758 5148 16764 5160
rect 16719 5120 16764 5148
rect 13613 5111 13671 5117
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 18414 5148 18420 5160
rect 18375 5120 18420 5148
rect 18414 5108 18420 5120
rect 18472 5108 18478 5160
rect 26252 5148 26280 5315
rect 26602 5312 26608 5324
rect 26660 5312 26666 5364
rect 26510 5244 26516 5296
rect 26568 5284 26574 5296
rect 26973 5287 27031 5293
rect 26973 5284 26985 5287
rect 26568 5256 26985 5284
rect 26568 5244 26574 5256
rect 26973 5253 26985 5256
rect 27019 5253 27031 5287
rect 26973 5247 27031 5253
rect 26421 5151 26479 5157
rect 26421 5148 26433 5151
rect 26252 5120 26433 5148
rect 26421 5117 26433 5120
rect 26467 5117 26479 5151
rect 26421 5111 26479 5117
rect 5353 5083 5411 5089
rect 5353 5049 5365 5083
rect 5399 5080 5411 5083
rect 5810 5080 5816 5092
rect 5399 5052 5816 5080
rect 5399 5049 5411 5052
rect 5353 5043 5411 5049
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 18506 5080 18512 5092
rect 17788 5052 18512 5080
rect 17788 5024 17816 5052
rect 18506 5040 18512 5052
rect 18564 5040 18570 5092
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 1452 4984 1593 5012
rect 1452 4972 1458 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 2682 5012 2688 5024
rect 2643 4984 2688 5012
rect 1581 4975 1639 4981
rect 2682 4972 2688 4984
rect 2740 4972 2746 5024
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3016 4984 3801 5012
rect 3016 4972 3022 4984
rect 3789 4981 3801 4984
rect 3835 5012 3847 5015
rect 4338 5012 4344 5024
rect 3835 4984 4344 5012
rect 3835 4981 3847 4984
rect 3789 4975 3847 4981
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 5718 5012 5724 5024
rect 5679 4984 5724 5012
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 14734 5012 14740 5024
rect 14695 4984 14740 5012
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 16298 5012 16304 5024
rect 16211 4984 16304 5012
rect 16298 4972 16304 4984
rect 16356 5012 16362 5024
rect 16850 5012 16856 5024
rect 16356 4984 16856 5012
rect 16356 4972 16362 4984
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 17494 5012 17500 5024
rect 17455 4984 17500 5012
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 2590 4808 2596 4820
rect 2087 4780 2596 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 2958 4808 2964 4820
rect 2871 4780 2964 4808
rect 2409 4743 2467 4749
rect 2409 4709 2421 4743
rect 2455 4740 2467 4743
rect 2884 4740 2912 4780
rect 2958 4768 2964 4780
rect 3016 4808 3022 4820
rect 4065 4811 4123 4817
rect 4065 4808 4077 4811
rect 3016 4780 4077 4808
rect 3016 4768 3022 4780
rect 4065 4777 4077 4780
rect 4111 4777 4123 4811
rect 4065 4771 4123 4777
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 5776 4780 7297 4808
rect 5776 4768 5782 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 7285 4771 7343 4777
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 12894 4808 12900 4820
rect 12759 4780 12900 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 13354 4808 13360 4820
rect 13315 4780 13360 4808
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 14366 4808 14372 4820
rect 14327 4780 14372 4808
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15746 4808 15752 4820
rect 15707 4780 15752 4808
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16485 4811 16543 4817
rect 16485 4777 16497 4811
rect 16531 4808 16543 4811
rect 16758 4808 16764 4820
rect 16531 4780 16764 4808
rect 16531 4777 16543 4780
rect 16485 4771 16543 4777
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 17678 4808 17684 4820
rect 17639 4780 17684 4808
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 18414 4808 18420 4820
rect 18187 4780 18420 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 26694 4808 26700 4820
rect 26655 4780 26700 4808
rect 26694 4768 26700 4780
rect 26752 4768 26758 4820
rect 3050 4740 3056 4752
rect 2455 4712 2912 4740
rect 3011 4712 3056 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 15657 4743 15715 4749
rect 15657 4709 15669 4743
rect 15703 4740 15715 4743
rect 15838 4740 15844 4752
rect 15703 4712 15844 4740
rect 15703 4709 15715 4712
rect 15657 4703 15715 4709
rect 15838 4700 15844 4712
rect 15896 4700 15902 4752
rect 17405 4743 17463 4749
rect 17405 4709 17417 4743
rect 17451 4740 17463 4743
rect 17586 4740 17592 4752
rect 17451 4712 17592 4740
rect 17451 4709 17463 4712
rect 17405 4703 17463 4709
rect 17586 4700 17592 4712
rect 17644 4700 17650 4752
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1578 4672 1584 4684
rect 1443 4644 1584 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1578 4632 1584 4644
rect 1636 4672 1642 4684
rect 1854 4672 1860 4684
rect 1636 4644 1860 4672
rect 1636 4632 1642 4644
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 2866 4672 2872 4684
rect 2547 4644 2872 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 3881 4675 3939 4681
rect 3881 4641 3893 4675
rect 3927 4672 3939 4675
rect 3970 4672 3976 4684
rect 3927 4644 3976 4672
rect 3927 4641 3939 4644
rect 3881 4635 3939 4641
rect 3970 4632 3976 4644
rect 4028 4672 4034 4684
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 4028 4644 4445 4672
rect 4028 4632 4034 4644
rect 4433 4641 4445 4644
rect 4479 4641 4491 4675
rect 4433 4635 4491 4641
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 6161 4675 6219 4681
rect 6161 4672 6173 4675
rect 5868 4644 6173 4672
rect 5868 4632 5874 4644
rect 6161 4641 6173 4644
rect 6207 4641 6219 4675
rect 6161 4635 6219 4641
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4672 12863 4675
rect 13078 4672 13084 4684
rect 12851 4644 13084 4672
rect 12851 4641 12863 4644
rect 12805 4635 12863 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 26510 4672 26516 4684
rect 26471 4644 26516 4672
rect 26510 4632 26516 4644
rect 26568 4632 26574 4684
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 4120 4576 4537 4604
rect 4120 4564 4126 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4706 4604 4712 4616
rect 4619 4576 4712 4604
rect 4525 4567 4583 4573
rect 4706 4564 4712 4576
rect 4764 4604 4770 4616
rect 5718 4604 5724 4616
rect 4764 4576 5724 4604
rect 4764 4564 4770 4576
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 1670 4428 1676 4480
rect 1728 4468 1734 4480
rect 2685 4471 2743 4477
rect 2685 4468 2697 4471
rect 1728 4440 2697 4468
rect 1728 4428 1734 4440
rect 2685 4437 2697 4440
rect 2731 4437 2743 4471
rect 5920 4468 5948 4567
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 12897 4607 12955 4613
rect 12897 4604 12909 4607
rect 12768 4576 12909 4604
rect 12768 4564 12774 4576
rect 12897 4573 12909 4576
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15436 4576 15853 4604
rect 15436 4564 15442 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 6270 4468 6276 4480
rect 5920 4440 6276 4468
rect 2685 4431 2743 4437
rect 6270 4428 6276 4440
rect 6328 4428 6334 4480
rect 12342 4468 12348 4480
rect 12303 4440 12348 4468
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 3970 4264 3976 4276
rect 3931 4236 3976 4264
rect 3970 4224 3976 4236
rect 4028 4224 4034 4276
rect 5445 4267 5503 4273
rect 5445 4233 5457 4267
rect 5491 4264 5503 4267
rect 5718 4264 5724 4276
rect 5491 4236 5724 4264
rect 5491 4233 5503 4236
rect 5445 4227 5503 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 12253 4267 12311 4273
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12894 4264 12900 4276
rect 12299 4236 12900 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12894 4224 12900 4236
rect 12952 4224 12958 4276
rect 13078 4264 13084 4276
rect 13039 4236 13084 4264
rect 13078 4224 13084 4236
rect 13136 4224 13142 4276
rect 15378 4264 15384 4276
rect 15339 4236 15384 4264
rect 15378 4224 15384 4236
rect 15436 4224 15442 4276
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 16117 4267 16175 4273
rect 16117 4264 16129 4267
rect 15804 4236 16129 4264
rect 15804 4224 15810 4236
rect 16117 4233 16129 4236
rect 16163 4233 16175 4267
rect 16117 4227 16175 4233
rect 26510 4224 26516 4276
rect 26568 4264 26574 4276
rect 27341 4267 27399 4273
rect 27341 4264 27353 4267
rect 26568 4236 27353 4264
rect 26568 4224 26574 4236
rect 27341 4233 27353 4236
rect 27387 4233 27399 4267
rect 27341 4227 27399 4233
rect 15838 4196 15844 4208
rect 15192 4168 15844 4196
rect 1946 4128 1952 4140
rect 1412 4100 1952 4128
rect 1412 4069 1440 4100
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 3418 4128 3424 4140
rect 3379 4100 3424 4128
rect 3418 4088 3424 4100
rect 3476 4128 3482 4140
rect 4614 4128 4620 4140
rect 3476 4100 4384 4128
rect 4575 4100 4620 4128
rect 3476 4088 3482 4100
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4029 1455 4063
rect 1397 4023 1455 4029
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 2501 4063 2559 4069
rect 2501 4060 2513 4063
rect 2455 4032 2513 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 2501 4029 2513 4032
rect 2547 4060 2559 4063
rect 3436 4060 3464 4088
rect 4356 4069 4384 4100
rect 4614 4088 4620 4100
rect 4672 4128 4678 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4672 4100 4997 4128
rect 4672 4088 4678 4100
rect 4985 4097 4997 4100
rect 5031 4128 5043 4131
rect 5810 4128 5816 4140
rect 5031 4100 5816 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5810 4088 5816 4100
rect 5868 4128 5874 4140
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5868 4100 5917 4128
rect 5868 4088 5874 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4128 15071 4131
rect 15192 4128 15220 4168
rect 15838 4156 15844 4168
rect 15896 4156 15902 4208
rect 15059 4100 15220 4128
rect 15059 4097 15071 4100
rect 15013 4091 15071 4097
rect 2547 4032 3464 4060
rect 4341 4063 4399 4069
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 8478 4060 8484 4072
rect 7699 4032 8484 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 15841 4063 15899 4069
rect 15841 4029 15853 4063
rect 15887 4060 15899 4063
rect 16482 4060 16488 4072
rect 15887 4032 16488 4060
rect 15887 4029 15899 4032
rect 15841 4023 15899 4029
rect 16482 4020 16488 4032
rect 16540 4020 16546 4072
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 26421 4063 26479 4069
rect 26421 4060 26433 4063
rect 26384 4032 26433 4060
rect 26384 4020 26390 4032
rect 26421 4029 26433 4032
rect 26467 4060 26479 4063
rect 26973 4063 27031 4069
rect 26973 4060 26985 4063
rect 26467 4032 26985 4060
rect 26467 4029 26479 4032
rect 26421 4023 26479 4029
rect 26973 4029 26985 4032
rect 27019 4029 27031 4063
rect 26973 4023 27031 4029
rect 2866 3952 2872 4004
rect 2924 3992 2930 4004
rect 3145 3995 3203 4001
rect 3145 3992 3157 3995
rect 2924 3964 3157 3992
rect 2924 3952 2930 3964
rect 3145 3961 3157 3964
rect 3191 3992 3203 3995
rect 4522 3992 4528 4004
rect 3191 3964 4528 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 7929 3995 7987 4001
rect 7929 3992 7941 3995
rect 5684 3964 7941 3992
rect 5684 3952 5690 3964
rect 7929 3961 7941 3964
rect 7975 3961 7987 3995
rect 7929 3955 7987 3961
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2774 3924 2780 3936
rect 2731 3896 2780 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 3881 3927 3939 3933
rect 3881 3924 3893 3927
rect 3752 3896 3893 3924
rect 3752 3884 3758 3896
rect 3881 3893 3893 3896
rect 3927 3924 3939 3927
rect 4430 3924 4436 3936
rect 3927 3896 4436 3924
rect 3927 3893 3939 3896
rect 3881 3887 3939 3893
rect 4430 3884 4436 3896
rect 4488 3884 4494 3936
rect 6270 3924 6276 3936
rect 6231 3896 6276 3924
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 12710 3924 12716 3936
rect 12671 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 26602 3924 26608 3936
rect 26563 3896 26608 3924
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 1949 3723 2007 3729
rect 1949 3720 1961 3723
rect 1912 3692 1961 3720
rect 1912 3680 1918 3692
rect 1949 3689 1961 3692
rect 1995 3689 2007 3723
rect 1949 3683 2007 3689
rect 3145 3723 3203 3729
rect 3145 3689 3157 3723
rect 3191 3720 3203 3723
rect 3234 3720 3240 3732
rect 3191 3692 3240 3720
rect 3191 3689 3203 3692
rect 3145 3683 3203 3689
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4062 3720 4068 3732
rect 3927 3692 4068 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4433 3723 4491 3729
rect 4433 3689 4445 3723
rect 4479 3720 4491 3723
rect 4522 3720 4528 3732
rect 4479 3692 4528 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 14090 3720 14096 3732
rect 13412 3692 14096 3720
rect 13412 3680 13418 3692
rect 14090 3680 14096 3692
rect 14148 3720 14154 3732
rect 14918 3720 14924 3732
rect 14148 3692 14924 3720
rect 14148 3680 14154 3692
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 26694 3720 26700 3732
rect 26655 3692 26700 3720
rect 26694 3680 26700 3692
rect 26752 3680 26758 3732
rect 8478 3612 8484 3664
rect 8536 3652 8542 3664
rect 8665 3655 8723 3661
rect 8665 3652 8677 3655
rect 8536 3624 8677 3652
rect 8536 3612 8542 3624
rect 8665 3621 8677 3624
rect 8711 3652 8723 3655
rect 11514 3652 11520 3664
rect 8711 3624 11520 3652
rect 8711 3621 8723 3624
rect 8665 3615 8723 3621
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3584 1455 3587
rect 2222 3584 2228 3596
rect 1443 3556 2228 3584
rect 1443 3553 1455 3556
rect 1397 3547 1455 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2501 3587 2559 3593
rect 2501 3553 2513 3587
rect 2547 3584 2559 3587
rect 2682 3584 2688 3596
rect 2547 3556 2688 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 2682 3544 2688 3556
rect 2740 3544 2746 3596
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 4798 3584 4804 3596
rect 4571 3556 4804 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 9769 3587 9827 3593
rect 9769 3553 9781 3587
rect 9815 3584 9827 3587
rect 9950 3584 9956 3596
rect 9815 3556 9956 3584
rect 9815 3553 9827 3556
rect 9769 3547 9827 3553
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 11072 3593 11100 3624
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3553 11115 3587
rect 11057 3547 11115 3553
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 11313 3587 11371 3593
rect 11313 3584 11325 3587
rect 11204 3556 11325 3584
rect 11204 3544 11210 3556
rect 11313 3553 11325 3556
rect 11359 3553 11371 3587
rect 11313 3547 11371 3553
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 14516 3556 15301 3584
rect 14516 3544 14522 3556
rect 15289 3553 15301 3556
rect 15335 3584 15347 3587
rect 16482 3584 16488 3596
rect 15335 3556 16488 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 25314 3584 25320 3596
rect 25275 3556 25320 3584
rect 25314 3544 25320 3556
rect 25372 3544 25378 3596
rect 26513 3587 26571 3593
rect 26513 3553 26525 3587
rect 26559 3553 26571 3587
rect 26513 3547 26571 3553
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 4672 3488 4717 3516
rect 4672 3476 4678 3488
rect 25038 3476 25044 3528
rect 25096 3516 25102 3528
rect 26528 3516 26556 3547
rect 27338 3516 27344 3528
rect 25096 3488 27344 3516
rect 25096 3476 25102 3488
rect 27338 3476 27344 3488
rect 27396 3476 27402 3528
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 4338 3340 4344 3392
rect 4396 3380 4402 3392
rect 5077 3383 5135 3389
rect 5077 3380 5089 3383
rect 4396 3352 5089 3380
rect 4396 3340 4402 3352
rect 5077 3349 5089 3352
rect 5123 3349 5135 3383
rect 5077 3343 5135 3349
rect 9953 3383 10011 3389
rect 9953 3349 9965 3383
rect 9999 3380 10011 3383
rect 11790 3380 11796 3392
rect 9999 3352 11796 3380
rect 9999 3349 10011 3352
rect 9953 3343 10011 3349
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 12434 3380 12440 3392
rect 12395 3352 12440 3380
rect 12434 3340 12440 3352
rect 12492 3340 12498 3392
rect 15473 3383 15531 3389
rect 15473 3349 15485 3383
rect 15519 3380 15531 3383
rect 15838 3380 15844 3392
rect 15519 3352 15844 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 25498 3380 25504 3392
rect 25459 3352 25504 3380
rect 25498 3340 25504 3352
rect 25556 3340 25562 3392
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 2222 3176 2228 3188
rect 2183 3148 2228 3176
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 2590 3176 2596 3188
rect 2551 3148 2596 3176
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 3605 3179 3663 3185
rect 3605 3145 3617 3179
rect 3651 3176 3663 3179
rect 4614 3176 4620 3188
rect 3651 3148 4620 3176
rect 3651 3145 3663 3148
rect 3605 3139 3663 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 4798 3176 4804 3188
rect 4759 3148 4804 3176
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5258 3176 5264 3188
rect 5219 3148 5264 3176
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 6546 3176 6552 3188
rect 6227 3148 6552 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 3973 3111 4031 3117
rect 3973 3077 3985 3111
rect 4019 3108 4031 3111
rect 4522 3108 4528 3120
rect 4019 3080 4528 3108
rect 4019 3077 4031 3080
rect 3973 3071 4031 3077
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 4632 3108 4660 3136
rect 5718 3108 5724 3120
rect 4632 3080 5724 3108
rect 5718 3068 5724 3080
rect 5776 3068 5782 3120
rect 3234 3040 3240 3052
rect 2792 3012 3240 3040
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 1486 2972 1492 2984
rect 1443 2944 1492 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 1486 2932 1492 2944
rect 1544 2972 1550 2984
rect 2038 2972 2044 2984
rect 1544 2944 2044 2972
rect 1544 2932 1550 2944
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2792 2981 2820 3012
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 2777 2975 2835 2981
rect 2777 2941 2789 2975
rect 2823 2941 2835 2975
rect 2777 2935 2835 2941
rect 3053 2975 3111 2981
rect 3053 2941 3065 2975
rect 3099 2972 3111 2975
rect 3510 2972 3516 2984
rect 3099 2944 3516 2972
rect 3099 2941 3111 2944
rect 3053 2935 3111 2941
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 4065 2975 4123 2981
rect 4065 2941 4077 2975
rect 4111 2972 4123 2975
rect 5258 2972 5264 2984
rect 4111 2944 5264 2972
rect 4111 2941 4123 2944
rect 4065 2935 4123 2941
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2972 5411 2975
rect 6196 2972 6224 3139
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 9950 3176 9956 3188
rect 9911 3148 9956 3176
rect 9950 3136 9956 3148
rect 10008 3176 10014 3188
rect 10505 3179 10563 3185
rect 10505 3176 10517 3179
rect 10008 3148 10517 3176
rect 10008 3136 10014 3148
rect 10505 3145 10517 3148
rect 10551 3145 10563 3179
rect 10505 3139 10563 3145
rect 11609 3179 11667 3185
rect 11609 3145 11621 3179
rect 11655 3176 11667 3179
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11655 3148 11897 3176
rect 11655 3145 11667 3148
rect 11609 3139 11667 3145
rect 11885 3145 11897 3148
rect 11931 3176 11943 3179
rect 12434 3176 12440 3188
rect 11931 3148 12440 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 14458 3176 14464 3188
rect 14419 3148 14464 3176
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 25130 3176 25136 3188
rect 25091 3148 25136 3176
rect 25130 3136 25136 3148
rect 25188 3136 25194 3188
rect 25314 3136 25320 3188
rect 25372 3176 25378 3188
rect 25869 3179 25927 3185
rect 25869 3176 25881 3179
rect 25372 3148 25881 3176
rect 25372 3136 25378 3148
rect 25869 3145 25881 3148
rect 25915 3145 25927 3179
rect 26602 3176 26608 3188
rect 26563 3148 26608 3176
rect 25869 3139 25927 3145
rect 26602 3136 26608 3148
rect 26660 3136 26666 3188
rect 27338 3176 27344 3188
rect 27299 3148 27344 3176
rect 27338 3136 27344 3148
rect 27396 3136 27402 3188
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 8573 3043 8631 3049
rect 8573 3040 8585 3043
rect 8536 3012 8585 3040
rect 8536 3000 8542 3012
rect 8573 3009 8585 3012
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 11204 3012 12173 3040
rect 11204 3000 11210 3012
rect 12161 3009 12173 3012
rect 12207 3040 12219 3043
rect 12342 3040 12348 3052
rect 12207 3012 12348 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12710 2981 12716 2984
rect 5399 2944 6224 2972
rect 11241 2975 11299 2981
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11609 2975 11667 2981
rect 11609 2972 11621 2975
rect 11287 2944 11621 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11609 2941 11621 2944
rect 11655 2941 11667 2975
rect 11609 2935 11667 2941
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2941 12495 2975
rect 12704 2972 12716 2981
rect 12671 2944 12716 2972
rect 12437 2935 12495 2941
rect 12704 2935 12716 2944
rect 12768 2972 12774 2984
rect 14734 2972 14740 2984
rect 12768 2944 14740 2972
rect 474 2864 480 2916
rect 532 2904 538 2916
rect 1673 2907 1731 2913
rect 1673 2904 1685 2907
rect 532 2876 1685 2904
rect 532 2864 538 2876
rect 1673 2873 1685 2876
rect 1719 2873 1731 2907
rect 1673 2867 1731 2873
rect 4341 2907 4399 2913
rect 4341 2873 4353 2907
rect 4387 2904 4399 2907
rect 4522 2904 4528 2916
rect 4387 2876 4528 2904
rect 4387 2873 4399 2876
rect 4341 2867 4399 2873
rect 4522 2864 4528 2876
rect 4580 2864 4586 2916
rect 5534 2864 5540 2916
rect 5592 2904 5598 2916
rect 5629 2907 5687 2913
rect 5629 2904 5641 2907
rect 5592 2876 5641 2904
rect 5592 2864 5598 2876
rect 5629 2873 5641 2876
rect 5675 2873 5687 2907
rect 8818 2907 8876 2913
rect 8818 2904 8830 2907
rect 5629 2867 5687 2873
rect 8404 2876 8830 2904
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8404 2845 8432 2876
rect 8818 2873 8830 2876
rect 8864 2904 8876 2907
rect 11057 2907 11115 2913
rect 11057 2904 11069 2907
rect 8864 2876 11069 2904
rect 8864 2873 8876 2876
rect 8818 2867 8876 2873
rect 11057 2873 11069 2876
rect 11103 2904 11115 2907
rect 11146 2904 11152 2916
rect 11103 2876 11152 2904
rect 11103 2873 11115 2876
rect 11057 2867 11115 2873
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 12452 2904 12480 2935
rect 12710 2932 12716 2935
rect 12768 2932 12774 2944
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 14918 2972 14924 2984
rect 14879 2944 14924 2972
rect 14918 2932 14924 2944
rect 14976 2932 14982 2984
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18141 2975 18199 2981
rect 18141 2972 18153 2975
rect 18012 2944 18153 2972
rect 18012 2932 18018 2944
rect 18141 2941 18153 2944
rect 18187 2972 18199 2975
rect 18693 2975 18751 2981
rect 18693 2972 18705 2975
rect 18187 2944 18705 2972
rect 18187 2941 18199 2944
rect 18141 2935 18199 2941
rect 18693 2941 18705 2944
rect 18739 2941 18751 2975
rect 18693 2935 18751 2941
rect 25130 2932 25136 2984
rect 25188 2972 25194 2984
rect 25317 2975 25375 2981
rect 25317 2972 25329 2975
rect 25188 2944 25329 2972
rect 25188 2932 25194 2944
rect 25317 2941 25329 2944
rect 25363 2941 25375 2975
rect 26418 2972 26424 2984
rect 26379 2944 26424 2972
rect 25317 2935 25375 2941
rect 26418 2932 26424 2944
rect 26476 2972 26482 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26476 2944 26985 2972
rect 26476 2932 26482 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 27522 2972 27528 2984
rect 27483 2944 27528 2972
rect 26973 2935 27031 2941
rect 27522 2932 27528 2944
rect 27580 2972 27586 2984
rect 28077 2975 28135 2981
rect 28077 2972 28089 2975
rect 27580 2944 28089 2972
rect 27580 2932 27586 2944
rect 28077 2941 28089 2944
rect 28123 2941 28135 2975
rect 28077 2935 28135 2941
rect 12618 2904 12624 2916
rect 11440 2876 12296 2904
rect 12452 2876 12624 2904
rect 11440 2845 11468 2876
rect 8389 2839 8447 2845
rect 8389 2836 8401 2839
rect 8352 2808 8401 2836
rect 8352 2796 8358 2808
rect 8389 2805 8401 2808
rect 8435 2805 8447 2839
rect 8389 2799 8447 2805
rect 11425 2839 11483 2845
rect 11425 2805 11437 2839
rect 11471 2805 11483 2839
rect 12268 2836 12296 2876
rect 12618 2864 12624 2876
rect 12676 2864 12682 2916
rect 14752 2904 14780 2932
rect 15194 2913 15200 2916
rect 15166 2907 15200 2913
rect 15166 2904 15178 2907
rect 14752 2876 15178 2904
rect 15166 2873 15178 2876
rect 15252 2904 15258 2916
rect 15252 2876 15314 2904
rect 15166 2867 15200 2873
rect 15194 2864 15200 2867
rect 15252 2864 15258 2876
rect 12802 2836 12808 2848
rect 12268 2808 12808 2836
rect 11425 2799 11483 2805
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 13814 2836 13820 2848
rect 13775 2808 13820 2836
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 15286 2796 15292 2848
rect 15344 2836 15350 2848
rect 16301 2839 16359 2845
rect 16301 2836 16313 2839
rect 15344 2808 16313 2836
rect 15344 2796 15350 2808
rect 16301 2805 16313 2808
rect 16347 2805 16359 2839
rect 18322 2836 18328 2848
rect 18283 2808 18328 2836
rect 16301 2799 16359 2805
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 25498 2836 25504 2848
rect 25459 2808 25504 2836
rect 25498 2796 25504 2808
rect 25556 2796 25562 2848
rect 27706 2836 27712 2848
rect 27667 2808 27712 2836
rect 27706 2796 27712 2808
rect 27764 2796 27770 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 2038 2592 2044 2644
rect 2096 2632 2102 2644
rect 2225 2635 2283 2641
rect 2225 2632 2237 2635
rect 2096 2604 2237 2632
rect 2096 2592 2102 2604
rect 2225 2601 2237 2604
rect 2271 2601 2283 2635
rect 2225 2595 2283 2601
rect 2406 2592 2412 2644
rect 2464 2632 2470 2644
rect 2593 2635 2651 2641
rect 2593 2632 2605 2635
rect 2464 2604 2605 2632
rect 2464 2592 2470 2604
rect 2593 2601 2605 2604
rect 2639 2601 2651 2635
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 2593 2595 2651 2601
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 5718 2632 5724 2644
rect 5679 2604 5724 2632
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 11606 2632 11612 2644
rect 11567 2604 11612 2632
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 12066 2632 12072 2644
rect 12027 2604 12072 2632
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12805 2635 12863 2641
rect 12805 2632 12817 2635
rect 12492 2604 12817 2632
rect 12492 2592 12498 2604
rect 12805 2601 12817 2604
rect 12851 2632 12863 2635
rect 14090 2632 14096 2644
rect 12851 2604 14096 2632
rect 12851 2601 12863 2604
rect 12805 2595 12863 2601
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 14458 2632 14464 2644
rect 14419 2604 14464 2632
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 15194 2592 15200 2604
rect 15252 2632 15258 2644
rect 15252 2604 15761 2632
rect 15252 2592 15258 2604
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2496 1547 2499
rect 2424 2496 2452 2592
rect 1535 2468 2452 2496
rect 2777 2499 2835 2505
rect 1535 2465 1547 2468
rect 1489 2459 1547 2465
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 3344 2496 3372 2592
rect 4338 2524 4344 2576
rect 4396 2564 4402 2576
rect 6270 2564 6276 2576
rect 4396 2536 6276 2564
rect 4396 2524 4402 2536
rect 6270 2524 6276 2536
rect 6328 2524 6334 2576
rect 6733 2567 6791 2573
rect 6733 2533 6745 2567
rect 6779 2564 6791 2567
rect 7438 2567 7496 2573
rect 7438 2564 7450 2567
rect 6779 2536 7450 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 7438 2533 7450 2536
rect 7484 2564 7496 2567
rect 8202 2564 8208 2576
rect 7484 2536 8208 2564
rect 7484 2533 7496 2536
rect 7438 2527 7496 2533
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 11514 2564 11520 2576
rect 11195 2536 11520 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 4614 2505 4620 2508
rect 2823 2468 3372 2496
rect 3881 2499 3939 2505
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 3881 2465 3893 2499
rect 3927 2496 3939 2499
rect 4608 2496 4620 2505
rect 3927 2468 4620 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4608 2459 4620 2468
rect 4614 2456 4620 2459
rect 4672 2456 4678 2508
rect 6288 2496 6316 2524
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 6288 2468 7205 2496
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 12084 2496 12112 2592
rect 15733 2573 15761 2604
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 16853 2635 16911 2641
rect 16853 2632 16865 2635
rect 16632 2604 16865 2632
rect 16632 2592 16638 2604
rect 16853 2601 16865 2604
rect 16899 2601 16911 2635
rect 19610 2632 19616 2644
rect 19571 2604 19616 2632
rect 16853 2595 16911 2601
rect 19610 2592 19616 2604
rect 19668 2592 19674 2644
rect 23014 2632 23020 2644
rect 22975 2604 23020 2632
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 27062 2632 27068 2644
rect 27023 2604 27068 2632
rect 27062 2592 27068 2604
rect 27120 2592 27126 2644
rect 15718 2567 15776 2573
rect 15718 2533 15730 2567
rect 15764 2533 15776 2567
rect 15718 2527 15776 2533
rect 11471 2468 12112 2496
rect 13173 2499 13231 2505
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 13173 2465 13185 2499
rect 13219 2465 13231 2499
rect 14274 2496 14280 2508
rect 14187 2468 14280 2496
rect 13173 2459 13231 2465
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 2498 2428 2504 2440
rect 1811 2400 2504 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 4338 2428 4344 2440
rect 4299 2400 4344 2428
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 13188 2428 13216 2459
rect 14274 2456 14280 2468
rect 14332 2496 14338 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14332 2468 14841 2496
rect 14332 2456 14338 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 14918 2456 14924 2508
rect 14976 2496 14982 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 14976 2468 15485 2496
rect 14976 2456 14982 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2496 18383 2499
rect 18414 2496 18420 2508
rect 18371 2468 18420 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18414 2456 18420 2468
rect 18472 2496 18478 2508
rect 18877 2499 18935 2505
rect 18877 2496 18889 2499
rect 18472 2468 18889 2496
rect 18472 2456 18478 2468
rect 18877 2465 18889 2468
rect 18923 2465 18935 2499
rect 19426 2496 19432 2508
rect 19387 2468 19432 2496
rect 18877 2459 18935 2465
rect 19426 2456 19432 2468
rect 19484 2496 19490 2508
rect 19981 2499 20039 2505
rect 19981 2496 19993 2499
rect 19484 2468 19993 2496
rect 19484 2456 19490 2468
rect 19981 2465 19993 2468
rect 20027 2465 20039 2499
rect 22830 2496 22836 2508
rect 22791 2468 22836 2496
rect 19981 2459 20039 2465
rect 22830 2456 22836 2468
rect 22888 2496 22894 2508
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 22888 2468 23397 2496
rect 22888 2456 22894 2468
rect 23385 2465 23397 2468
rect 23431 2465 23443 2499
rect 24578 2496 24584 2508
rect 24539 2468 24584 2496
rect 23385 2459 23443 2465
rect 24578 2456 24584 2468
rect 24636 2496 24642 2508
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24636 2468 25145 2496
rect 24636 2456 24642 2468
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25682 2496 25688 2508
rect 25595 2468 25688 2496
rect 25133 2459 25191 2465
rect 25682 2456 25688 2468
rect 25740 2496 25746 2508
rect 26237 2499 26295 2505
rect 26237 2496 26249 2499
rect 25740 2468 26249 2496
rect 25740 2456 25746 2468
rect 26237 2465 26249 2468
rect 26283 2465 26295 2499
rect 26237 2459 26295 2465
rect 26786 2456 26792 2508
rect 26844 2496 26850 2508
rect 26881 2499 26939 2505
rect 26881 2496 26893 2499
rect 26844 2468 26893 2496
rect 26844 2456 26850 2468
rect 26881 2465 26893 2468
rect 26927 2496 26939 2499
rect 27433 2499 27491 2505
rect 27433 2496 27445 2499
rect 26927 2468 27445 2496
rect 26927 2465 26939 2468
rect 26881 2459 26939 2465
rect 27433 2465 27445 2468
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 13817 2431 13875 2437
rect 13817 2428 13829 2431
rect 13188 2400 13829 2428
rect 13817 2397 13829 2400
rect 13863 2428 13875 2431
rect 15102 2428 15108 2440
rect 13863 2400 15108 2428
rect 13863 2397 13875 2400
rect 13817 2391 13875 2397
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 13357 2363 13415 2369
rect 13357 2329 13369 2363
rect 13403 2360 13415 2363
rect 14918 2360 14924 2372
rect 13403 2332 14924 2360
rect 13403 2329 13415 2332
rect 13357 2323 13415 2329
rect 14918 2320 14924 2332
rect 14976 2320 14982 2372
rect 2958 2292 2964 2304
rect 2919 2264 2964 2292
rect 2958 2252 2964 2264
rect 3016 2252 3022 2304
rect 7834 2252 7840 2304
rect 7892 2292 7898 2304
rect 8570 2292 8576 2304
rect 7892 2264 8576 2292
rect 7892 2252 7898 2264
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 9953 2295 10011 2301
rect 9953 2261 9965 2295
rect 9999 2292 10011 2295
rect 10778 2292 10784 2304
rect 9999 2264 10784 2292
rect 9999 2261 10011 2264
rect 9953 2255 10011 2261
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 18506 2292 18512 2304
rect 18467 2264 18512 2292
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 24762 2292 24768 2304
rect 24723 2264 24768 2292
rect 24762 2252 24768 2264
rect 24820 2252 24826 2304
rect 25866 2292 25872 2304
rect 25827 2264 25872 2292
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
rect 19058 552 19064 604
rect 19116 592 19122 604
rect 19150 592 19156 604
rect 19116 564 19156 592
rect 19116 552 19122 564
rect 19150 552 19156 564
rect 19208 552 19214 604
<< via1 >>
rect 4068 22312 4120 22364
rect 2964 22176 3016 22228
rect 13176 22176 13228 22228
rect 12532 22108 12584 22160
rect 24860 22108 24912 22160
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 25320 21632 25372 21684
rect 25688 21632 25740 21684
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 14188 21020 14240 21072
rect 25780 21020 25832 21072
rect 3884 20952 3936 21004
rect 13176 20952 13228 21004
rect 20168 20952 20220 21004
rect 21548 20995 21600 21004
rect 21548 20961 21557 20995
rect 21557 20961 21591 20995
rect 21591 20961 21600 20995
rect 21548 20952 21600 20961
rect 3148 20884 3200 20936
rect 25688 20884 25740 20936
rect 8208 20816 8260 20868
rect 5172 20748 5224 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 9588 20544 9640 20596
rect 11336 20544 11388 20596
rect 19432 20544 19484 20596
rect 21548 20587 21600 20596
rect 21548 20553 21557 20587
rect 21557 20553 21591 20587
rect 21591 20553 21600 20587
rect 21548 20544 21600 20553
rect 22008 20544 22060 20596
rect 20628 20519 20680 20528
rect 20628 20485 20637 20519
rect 20637 20485 20671 20519
rect 20671 20485 20680 20519
rect 20628 20476 20680 20485
rect 23848 20519 23900 20528
rect 23848 20485 23857 20519
rect 23857 20485 23891 20519
rect 23891 20485 23900 20519
rect 23848 20476 23900 20485
rect 8576 20340 8628 20392
rect 12716 20340 12768 20392
rect 12716 20247 12768 20256
rect 12716 20213 12725 20247
rect 12725 20213 12759 20247
rect 12759 20213 12768 20247
rect 12716 20204 12768 20213
rect 16488 20247 16540 20256
rect 16488 20213 16497 20247
rect 16497 20213 16531 20247
rect 16531 20213 16540 20247
rect 16488 20204 16540 20213
rect 18236 20247 18288 20256
rect 18236 20213 18245 20247
rect 18245 20213 18279 20247
rect 18279 20213 18288 20247
rect 18236 20204 18288 20213
rect 18972 20340 19024 20392
rect 22284 20383 22336 20392
rect 22284 20349 22293 20383
rect 22293 20349 22327 20383
rect 22327 20349 22336 20383
rect 22284 20340 22336 20349
rect 23664 20383 23716 20392
rect 23664 20349 23673 20383
rect 23673 20349 23707 20383
rect 23707 20349 23716 20383
rect 23664 20340 23716 20349
rect 20168 20315 20220 20324
rect 20168 20281 20177 20315
rect 20177 20281 20211 20315
rect 20211 20281 20220 20315
rect 20168 20272 20220 20281
rect 20720 20272 20772 20324
rect 18880 20204 18932 20256
rect 21916 20247 21968 20256
rect 21916 20213 21925 20247
rect 21925 20213 21959 20247
rect 21959 20213 21968 20247
rect 21916 20204 21968 20213
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 18604 20043 18656 20052
rect 18604 20009 18613 20043
rect 18613 20009 18647 20043
rect 18647 20009 18656 20043
rect 18604 20000 18656 20009
rect 21548 20000 21600 20052
rect 17316 19907 17368 19916
rect 17316 19873 17325 19907
rect 17325 19873 17359 19907
rect 17359 19873 17368 19907
rect 17316 19864 17368 19873
rect 19432 19864 19484 19916
rect 20720 19864 20772 19916
rect 17500 19771 17552 19780
rect 17500 19737 17509 19771
rect 17509 19737 17543 19771
rect 17543 19737 17552 19771
rect 17500 19728 17552 19737
rect 19708 19771 19760 19780
rect 19708 19737 19717 19771
rect 19717 19737 19751 19771
rect 19751 19737 19760 19771
rect 19708 19728 19760 19737
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 17316 19499 17368 19508
rect 17316 19465 17325 19499
rect 17325 19465 17359 19499
rect 17359 19465 17368 19499
rect 17316 19456 17368 19465
rect 15752 19320 15804 19372
rect 16488 19320 16540 19372
rect 17408 19388 17460 19440
rect 17776 19388 17828 19440
rect 19064 19320 19116 19372
rect 14280 19252 14332 19304
rect 14556 19252 14608 19304
rect 19432 19184 19484 19236
rect 19800 19116 19852 19168
rect 20720 19116 20772 19168
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 19340 15988 19392 16040
rect 21364 15988 21416 16040
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 11796 14535 11848 14544
rect 11796 14501 11805 14535
rect 11805 14501 11839 14535
rect 11839 14501 11848 14535
rect 11796 14492 11848 14501
rect 11888 14467 11940 14476
rect 11888 14433 11897 14467
rect 11897 14433 11931 14467
rect 11931 14433 11940 14467
rect 11888 14424 11940 14433
rect 12164 14356 12216 14408
rect 12440 14220 12492 14272
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 11796 14016 11848 14068
rect 11888 14016 11940 14068
rect 2688 13812 2740 13864
rect 10784 13744 10836 13796
rect 12164 13880 12216 13932
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 13912 13855 13964 13864
rect 13912 13821 13946 13855
rect 13946 13821 13964 13855
rect 13912 13812 13964 13821
rect 1676 13719 1728 13728
rect 1676 13685 1685 13719
rect 1685 13685 1719 13719
rect 1719 13685 1728 13719
rect 1676 13676 1728 13685
rect 4896 13676 4948 13728
rect 10232 13719 10284 13728
rect 10232 13685 10241 13719
rect 10241 13685 10275 13719
rect 10275 13685 10284 13719
rect 10232 13676 10284 13685
rect 15016 13719 15068 13728
rect 15016 13685 15025 13719
rect 15025 13685 15059 13719
rect 15059 13685 15068 13719
rect 15016 13676 15068 13685
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 1676 13472 1728 13524
rect 2504 13472 2556 13524
rect 2780 13472 2832 13524
rect 11888 13472 11940 13524
rect 9496 13404 9548 13456
rect 12256 13404 12308 13456
rect 2688 13336 2740 13388
rect 4528 13336 4580 13388
rect 5264 13379 5316 13388
rect 5264 13345 5298 13379
rect 5298 13345 5316 13379
rect 5264 13336 5316 13345
rect 9956 13379 10008 13388
rect 9956 13345 9990 13379
rect 9990 13345 10008 13379
rect 9956 13336 10008 13345
rect 11796 13336 11848 13388
rect 12900 13336 12952 13388
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 4988 13311 5040 13320
rect 4988 13277 4997 13311
rect 4997 13277 5031 13311
rect 5031 13277 5040 13311
rect 4988 13268 5040 13277
rect 7656 13268 7708 13320
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 1860 13132 1912 13184
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 10784 13132 10836 13184
rect 13636 13132 13688 13184
rect 14924 13132 14976 13184
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 2872 12928 2924 12980
rect 2596 12860 2648 12912
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 3516 12928 3568 12980
rect 4528 12971 4580 12980
rect 4528 12937 4537 12971
rect 4537 12937 4571 12971
rect 4571 12937 4580 12971
rect 4528 12928 4580 12937
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 17960 12928 18012 12980
rect 9956 12860 10008 12912
rect 10140 12860 10192 12912
rect 12716 12860 12768 12912
rect 3608 12835 3660 12844
rect 1676 12724 1728 12776
rect 2780 12724 2832 12776
rect 3332 12767 3384 12776
rect 3332 12733 3341 12767
rect 3341 12733 3375 12767
rect 3375 12733 3384 12767
rect 3332 12724 3384 12733
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 5264 12792 5316 12844
rect 7656 12835 7708 12844
rect 4528 12724 4580 12776
rect 4896 12767 4948 12776
rect 4896 12733 4905 12767
rect 4905 12733 4939 12767
rect 4939 12733 4948 12767
rect 4896 12724 4948 12733
rect 4436 12699 4488 12708
rect 4436 12665 4445 12699
rect 4445 12665 4479 12699
rect 4479 12665 4488 12699
rect 5080 12724 5132 12776
rect 4436 12656 4488 12665
rect 3332 12588 3384 12640
rect 4068 12631 4120 12640
rect 4068 12597 4077 12631
rect 4077 12597 4111 12631
rect 4111 12597 4120 12631
rect 4068 12588 4120 12597
rect 7656 12801 7665 12835
rect 7665 12801 7699 12835
rect 7699 12801 7708 12835
rect 7656 12792 7708 12801
rect 9680 12792 9732 12844
rect 10232 12792 10284 12844
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 12900 12792 12952 12844
rect 12440 12724 12492 12776
rect 13084 12724 13136 12776
rect 14924 12767 14976 12776
rect 14924 12733 14933 12767
rect 14933 12733 14967 12767
rect 14967 12733 14976 12767
rect 14924 12724 14976 12733
rect 15016 12724 15068 12776
rect 6828 12588 6880 12640
rect 7196 12588 7248 12640
rect 10508 12631 10560 12640
rect 10508 12597 10517 12631
rect 10517 12597 10551 12631
rect 10551 12597 10560 12631
rect 10508 12588 10560 12597
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12440 12588 12492 12597
rect 16396 12588 16448 12640
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 1860 12384 1912 12436
rect 3608 12384 3660 12436
rect 4528 12427 4580 12436
rect 4528 12393 4537 12427
rect 4537 12393 4571 12427
rect 4571 12393 4580 12427
rect 4528 12384 4580 12393
rect 4988 12427 5040 12436
rect 4988 12393 4997 12427
rect 4997 12393 5031 12427
rect 5031 12393 5040 12427
rect 4988 12384 5040 12393
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 10508 12384 10560 12436
rect 10784 12427 10836 12436
rect 10784 12393 10793 12427
rect 10793 12393 10827 12427
rect 10827 12393 10836 12427
rect 10784 12384 10836 12393
rect 11428 12384 11480 12436
rect 12440 12384 12492 12436
rect 12900 12384 12952 12436
rect 13084 12427 13136 12436
rect 13084 12393 13093 12427
rect 13093 12393 13127 12427
rect 13127 12393 13136 12427
rect 13084 12384 13136 12393
rect 13728 12384 13780 12436
rect 2044 12316 2096 12368
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 6368 12316 6420 12368
rect 5816 12291 5868 12300
rect 2780 12248 2832 12257
rect 5816 12257 5825 12291
rect 5825 12257 5859 12291
rect 5859 12257 5868 12291
rect 5816 12248 5868 12257
rect 10692 12248 10744 12300
rect 12440 12248 12492 12300
rect 13544 12248 13596 12300
rect 14924 12248 14976 12300
rect 16948 12316 17000 12368
rect 16580 12248 16632 12300
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 4068 12180 4120 12232
rect 9036 12180 9088 12232
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 12348 12223 12400 12232
rect 10232 12180 10284 12189
rect 12348 12189 12357 12223
rect 12357 12189 12391 12223
rect 12391 12189 12400 12223
rect 12348 12180 12400 12189
rect 13820 12223 13872 12232
rect 13820 12189 13829 12223
rect 13829 12189 13863 12223
rect 13863 12189 13872 12223
rect 13820 12180 13872 12189
rect 26240 12112 26292 12164
rect 26516 12112 26568 12164
rect 11704 12087 11756 12096
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 12808 12044 12860 12096
rect 15476 12044 15528 12096
rect 16488 12044 16540 12096
rect 18236 12044 18288 12096
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 2504 11840 2556 11892
rect 2780 11883 2832 11892
rect 2780 11849 2789 11883
rect 2789 11849 2823 11883
rect 2823 11849 2832 11883
rect 2780 11840 2832 11849
rect 3608 11840 3660 11892
rect 4068 11840 4120 11892
rect 6368 11840 6420 11892
rect 9404 11883 9456 11892
rect 9404 11849 9413 11883
rect 9413 11849 9447 11883
rect 9447 11849 9456 11883
rect 9404 11840 9456 11849
rect 9588 11883 9640 11892
rect 9588 11849 9597 11883
rect 9597 11849 9631 11883
rect 9631 11849 9640 11883
rect 9588 11840 9640 11849
rect 11428 11883 11480 11892
rect 11428 11849 11437 11883
rect 11437 11849 11471 11883
rect 11471 11849 11480 11883
rect 11428 11840 11480 11849
rect 12440 11883 12492 11892
rect 12440 11849 12449 11883
rect 12449 11849 12483 11883
rect 12483 11849 12492 11883
rect 16580 11883 16632 11892
rect 12440 11840 12492 11849
rect 16580 11849 16589 11883
rect 16589 11849 16623 11883
rect 16623 11849 16632 11883
rect 16580 11840 16632 11849
rect 18236 11883 18288 11892
rect 18236 11849 18245 11883
rect 18245 11849 18279 11883
rect 18279 11849 18288 11883
rect 18236 11840 18288 11849
rect 18696 11840 18748 11892
rect 2688 11704 2740 11756
rect 5816 11772 5868 11824
rect 6736 11772 6788 11824
rect 12348 11772 12400 11824
rect 10232 11704 10284 11756
rect 12900 11704 12952 11756
rect 9404 11636 9456 11688
rect 9772 11636 9824 11688
rect 12164 11636 12216 11688
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 13452 11636 13504 11688
rect 13820 11636 13872 11688
rect 16948 11679 17000 11688
rect 16948 11645 16957 11679
rect 16957 11645 16991 11679
rect 16991 11645 17000 11679
rect 16948 11636 17000 11645
rect 18512 11636 18564 11688
rect 18696 11679 18748 11688
rect 18696 11645 18730 11679
rect 18730 11645 18748 11679
rect 18696 11636 18748 11645
rect 26424 11679 26476 11688
rect 26424 11645 26433 11679
rect 26433 11645 26467 11679
rect 26467 11645 26476 11679
rect 26424 11636 26476 11645
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 2504 11500 2556 11552
rect 3332 11568 3384 11620
rect 9036 11611 9088 11620
rect 9036 11577 9045 11611
rect 9045 11577 9079 11611
rect 9079 11577 9088 11611
rect 9036 11568 9088 11577
rect 13544 11611 13596 11620
rect 13544 11577 13553 11611
rect 13553 11577 13587 11611
rect 13587 11577 13596 11611
rect 13544 11568 13596 11577
rect 3424 11500 3476 11552
rect 9956 11543 10008 11552
rect 9956 11509 9965 11543
rect 9965 11509 9999 11543
rect 9999 11509 10008 11543
rect 9956 11500 10008 11509
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 13084 11500 13136 11552
rect 13728 11500 13780 11552
rect 19432 11500 19484 11552
rect 26608 11543 26660 11552
rect 26608 11509 26617 11543
rect 26617 11509 26651 11543
rect 26651 11509 26660 11543
rect 26608 11500 26660 11509
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 2872 11296 2924 11348
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 6920 11296 6972 11348
rect 10232 11339 10284 11348
rect 10232 11305 10241 11339
rect 10241 11305 10275 11339
rect 10275 11305 10284 11339
rect 10232 11296 10284 11305
rect 12440 11296 12492 11348
rect 12900 11339 12952 11348
rect 12900 11305 12909 11339
rect 12909 11305 12943 11339
rect 12943 11305 12952 11339
rect 12900 11296 12952 11305
rect 13544 11296 13596 11348
rect 14004 11296 14056 11348
rect 7104 11228 7156 11280
rect 12164 11271 12216 11280
rect 12164 11237 12173 11271
rect 12173 11237 12207 11271
rect 12207 11237 12216 11271
rect 12164 11228 12216 11237
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 4620 11160 4672 11212
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 13268 11203 13320 11212
rect 13268 11169 13277 11203
rect 13277 11169 13311 11203
rect 13311 11169 13320 11203
rect 13268 11160 13320 11169
rect 17316 11160 17368 11212
rect 17684 11203 17736 11212
rect 17684 11169 17693 11203
rect 17693 11169 17727 11203
rect 17727 11169 17736 11203
rect 17684 11160 17736 11169
rect 26516 11203 26568 11212
rect 26516 11169 26525 11203
rect 26525 11169 26559 11203
rect 26559 11169 26568 11203
rect 26516 11160 26568 11169
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 2412 11024 2464 11076
rect 3608 11092 3660 11144
rect 4344 11092 4396 11144
rect 4528 11135 4580 11144
rect 4528 11101 4537 11135
rect 4537 11101 4571 11135
rect 4571 11101 4580 11135
rect 4528 11092 4580 11101
rect 4896 11092 4948 11144
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 17408 11092 17460 11144
rect 18236 11092 18288 11144
rect 9956 11067 10008 11076
rect 9956 11033 9965 11067
rect 9965 11033 9999 11067
rect 9999 11033 10008 11067
rect 9956 11024 10008 11033
rect 10416 11024 10468 11076
rect 16488 11067 16540 11076
rect 16488 11033 16497 11067
rect 16497 11033 16531 11067
rect 16531 11033 16540 11067
rect 16488 11024 16540 11033
rect 26700 11067 26752 11076
rect 26700 11033 26709 11067
rect 26709 11033 26743 11067
rect 26743 11033 26752 11067
rect 26700 11024 26752 11033
rect 16764 10956 16816 11008
rect 18420 10999 18472 11008
rect 18420 10965 18429 10999
rect 18429 10965 18463 10999
rect 18463 10965 18472 10999
rect 18420 10956 18472 10965
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2044 10795 2096 10804
rect 2044 10761 2053 10795
rect 2053 10761 2087 10795
rect 2087 10761 2096 10795
rect 2044 10752 2096 10761
rect 2412 10795 2464 10804
rect 2412 10761 2421 10795
rect 2421 10761 2455 10795
rect 2455 10761 2464 10795
rect 2412 10752 2464 10761
rect 2780 10752 2832 10804
rect 6920 10752 6972 10804
rect 13268 10752 13320 10804
rect 13544 10795 13596 10804
rect 13544 10761 13553 10795
rect 13553 10761 13587 10795
rect 13587 10761 13596 10795
rect 13544 10752 13596 10761
rect 26516 10795 26568 10804
rect 26516 10761 26525 10795
rect 26525 10761 26559 10795
rect 26559 10761 26568 10795
rect 26516 10752 26568 10761
rect 4896 10616 4948 10668
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 10876 10616 10928 10668
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 16580 10616 16632 10668
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 17776 10659 17828 10668
rect 17776 10625 17785 10659
rect 17785 10625 17819 10659
rect 17819 10625 17828 10659
rect 17776 10616 17828 10625
rect 18236 10616 18288 10668
rect 18696 10616 18748 10668
rect 2044 10548 2096 10600
rect 10784 10480 10836 10532
rect 3424 10412 3476 10464
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 3700 10412 3752 10421
rect 4436 10412 4488 10464
rect 4620 10455 4672 10464
rect 4620 10421 4629 10455
rect 4629 10421 4663 10455
rect 4663 10421 4672 10455
rect 4620 10412 4672 10421
rect 4896 10412 4948 10464
rect 7104 10455 7156 10464
rect 7104 10421 7113 10455
rect 7113 10421 7147 10455
rect 7147 10421 7156 10455
rect 7104 10412 7156 10421
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 16764 10591 16816 10600
rect 16764 10557 16773 10591
rect 16773 10557 16807 10591
rect 16807 10557 16816 10591
rect 16764 10548 16816 10557
rect 18328 10548 18380 10600
rect 17040 10480 17092 10532
rect 11336 10412 11388 10464
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 16948 10412 17000 10464
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 18420 10455 18472 10464
rect 18420 10421 18429 10455
rect 18429 10421 18463 10455
rect 18463 10421 18472 10455
rect 18420 10412 18472 10421
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 3424 10208 3476 10260
rect 4528 10208 4580 10260
rect 6920 10251 6972 10260
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 8116 10208 8168 10260
rect 10876 10208 10928 10260
rect 13452 10208 13504 10260
rect 14004 10208 14056 10260
rect 14924 10208 14976 10260
rect 16856 10208 16908 10260
rect 9864 10140 9916 10192
rect 17224 10140 17276 10192
rect 18144 10208 18196 10260
rect 18696 10251 18748 10260
rect 18696 10217 18705 10251
rect 18705 10217 18739 10251
rect 18739 10217 18748 10251
rect 18696 10208 18748 10217
rect 26700 10251 26752 10260
rect 26700 10217 26709 10251
rect 26709 10217 26743 10251
rect 26743 10217 26752 10251
rect 26700 10208 26752 10217
rect 21364 10140 21416 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 4804 10072 4856 10124
rect 8208 10072 8260 10124
rect 14924 10115 14976 10124
rect 14924 10081 14933 10115
rect 14933 10081 14967 10115
rect 14967 10081 14976 10115
rect 14924 10072 14976 10081
rect 15660 10072 15712 10124
rect 15844 10072 15896 10124
rect 18052 10115 18104 10124
rect 18052 10081 18061 10115
rect 18061 10081 18095 10115
rect 18095 10081 18104 10115
rect 18052 10072 18104 10081
rect 26516 10115 26568 10124
rect 26516 10081 26525 10115
rect 26525 10081 26559 10115
rect 26559 10081 26568 10115
rect 26516 10072 26568 10081
rect 4896 10004 4948 10056
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 17040 10004 17092 10056
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 17408 10004 17460 10056
rect 18696 10004 18748 10056
rect 2872 9936 2924 9988
rect 2320 9868 2372 9920
rect 2964 9868 3016 9920
rect 16488 9868 16540 9920
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 1400 9664 1452 9716
rect 4252 9664 4304 9716
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 4896 9707 4948 9716
rect 4896 9673 4905 9707
rect 4905 9673 4939 9707
rect 4939 9673 4948 9707
rect 4896 9664 4948 9673
rect 7104 9664 7156 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 3148 9596 3200 9648
rect 4804 9596 4856 9648
rect 8116 9596 8168 9648
rect 9680 9664 9732 9716
rect 10784 9707 10836 9716
rect 10784 9673 10793 9707
rect 10793 9673 10827 9707
rect 10827 9673 10836 9707
rect 10784 9664 10836 9673
rect 11520 9664 11572 9716
rect 11980 9664 12032 9716
rect 10600 9639 10652 9648
rect 10600 9605 10609 9639
rect 10609 9605 10643 9639
rect 10643 9605 10652 9639
rect 10600 9596 10652 9605
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 10876 9528 10928 9580
rect 12072 9596 12124 9648
rect 11152 9503 11204 9512
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 7104 9435 7156 9444
rect 7104 9401 7138 9435
rect 7138 9401 7156 9435
rect 7104 9392 7156 9401
rect 9496 9392 9548 9444
rect 9864 9392 9916 9444
rect 11796 9528 11848 9580
rect 14004 9571 14056 9580
rect 14004 9537 14013 9571
rect 14013 9537 14047 9571
rect 14047 9537 14056 9571
rect 14004 9528 14056 9537
rect 18696 9664 18748 9716
rect 19524 9664 19576 9716
rect 19800 9664 19852 9716
rect 17960 9596 18012 9648
rect 17040 9460 17092 9512
rect 17316 9460 17368 9512
rect 17408 9392 17460 9444
rect 18512 9571 18564 9580
rect 18512 9537 18521 9571
rect 18521 9537 18555 9571
rect 18555 9537 18564 9571
rect 18512 9528 18564 9537
rect 18696 9571 18748 9580
rect 18696 9537 18705 9571
rect 18705 9537 18739 9571
rect 18739 9537 18748 9571
rect 18696 9528 18748 9537
rect 18420 9503 18472 9512
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 26516 9503 26568 9512
rect 26516 9469 26525 9503
rect 26525 9469 26559 9503
rect 26559 9469 26568 9503
rect 26516 9460 26568 9469
rect 19156 9392 19208 9444
rect 8300 9324 8352 9376
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 15384 9367 15436 9376
rect 15384 9333 15393 9367
rect 15393 9333 15427 9367
rect 15427 9333 15436 9367
rect 15384 9324 15436 9333
rect 15844 9324 15896 9376
rect 16488 9324 16540 9376
rect 16672 9324 16724 9376
rect 17224 9324 17276 9376
rect 18052 9367 18104 9376
rect 18052 9333 18061 9367
rect 18061 9333 18095 9367
rect 18095 9333 18104 9367
rect 18052 9324 18104 9333
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 10876 9163 10928 9172
rect 10876 9129 10885 9163
rect 10885 9129 10919 9163
rect 10919 9129 10928 9163
rect 10876 9120 10928 9129
rect 11336 9120 11388 9172
rect 11612 9120 11664 9172
rect 12164 9120 12216 9172
rect 14004 9163 14056 9172
rect 14004 9129 14013 9163
rect 14013 9129 14047 9163
rect 14047 9129 14056 9163
rect 14004 9120 14056 9129
rect 17776 9163 17828 9172
rect 17776 9129 17785 9163
rect 17785 9129 17819 9163
rect 17819 9129 17828 9163
rect 17776 9120 17828 9129
rect 18972 9120 19024 9172
rect 26700 9163 26752 9172
rect 26700 9129 26709 9163
rect 26709 9129 26743 9163
rect 26743 9129 26752 9163
rect 26700 9120 26752 9129
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 2504 9027 2556 9036
rect 2504 8993 2513 9027
rect 2513 8993 2547 9027
rect 2547 8993 2556 9027
rect 2504 8984 2556 8993
rect 6276 9052 6328 9104
rect 6828 9052 6880 9104
rect 16212 9095 16264 9104
rect 16212 9061 16221 9095
rect 16221 9061 16255 9095
rect 16255 9061 16264 9095
rect 16212 9052 16264 9061
rect 16856 9095 16908 9104
rect 16856 9061 16865 9095
rect 16865 9061 16899 9095
rect 16899 9061 16908 9095
rect 16856 9052 16908 9061
rect 17040 9052 17092 9104
rect 5816 8984 5868 9036
rect 11520 8984 11572 9036
rect 18512 8984 18564 9036
rect 19616 9052 19668 9104
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 11796 8959 11848 8968
rect 11796 8925 11805 8959
rect 11805 8925 11839 8959
rect 11839 8925 11848 8959
rect 11796 8916 11848 8925
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 17408 8916 17460 8968
rect 18696 8916 18748 8968
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 12256 8848 12308 8900
rect 2688 8823 2740 8832
rect 2688 8789 2697 8823
rect 2697 8789 2731 8823
rect 2731 8789 2740 8823
rect 2688 8780 2740 8789
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 9496 8780 9548 8832
rect 14372 8780 14424 8832
rect 14924 8780 14976 8832
rect 17960 8780 18012 8832
rect 18328 8780 18380 8832
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 2504 8576 2556 8585
rect 5816 8619 5868 8628
rect 5816 8585 5825 8619
rect 5825 8585 5859 8619
rect 5859 8585 5868 8619
rect 5816 8576 5868 8585
rect 7932 8576 7984 8628
rect 11612 8619 11664 8628
rect 11612 8585 11621 8619
rect 11621 8585 11655 8619
rect 11655 8585 11664 8619
rect 11612 8576 11664 8585
rect 16488 8576 16540 8628
rect 17132 8576 17184 8628
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 18512 8619 18564 8628
rect 18512 8585 18521 8619
rect 18521 8585 18555 8619
rect 18555 8585 18564 8619
rect 18512 8576 18564 8585
rect 18972 8576 19024 8628
rect 19892 8576 19944 8628
rect 26608 8619 26660 8628
rect 26608 8585 26617 8619
rect 26617 8585 26651 8619
rect 26651 8585 26660 8619
rect 26608 8576 26660 8585
rect 6276 8508 6328 8560
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 3148 8440 3200 8492
rect 3516 8440 3568 8492
rect 11520 8508 11572 8560
rect 14372 8508 14424 8560
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 18328 8483 18380 8492
rect 7656 8415 7708 8424
rect 7656 8381 7665 8415
rect 7665 8381 7699 8415
rect 7699 8381 7708 8415
rect 7656 8372 7708 8381
rect 9220 8415 9272 8424
rect 9220 8381 9229 8415
rect 9229 8381 9263 8415
rect 9263 8381 9272 8415
rect 9220 8372 9272 8381
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 7288 8279 7340 8288
rect 2780 8236 2832 8245
rect 7288 8245 7297 8279
rect 7297 8245 7331 8279
rect 7331 8245 7340 8279
rect 7288 8236 7340 8245
rect 9588 8304 9640 8356
rect 14096 8372 14148 8424
rect 14832 8415 14884 8424
rect 14832 8381 14841 8415
rect 14841 8381 14875 8415
rect 14875 8381 14884 8415
rect 14832 8372 14884 8381
rect 18328 8449 18337 8483
rect 18337 8449 18371 8483
rect 18371 8449 18380 8483
rect 19248 8508 19300 8560
rect 26516 8508 26568 8560
rect 27712 8551 27764 8560
rect 27712 8517 27721 8551
rect 27721 8517 27755 8551
rect 27755 8517 27764 8551
rect 27712 8508 27764 8517
rect 18328 8440 18380 8449
rect 19432 8440 19484 8492
rect 15384 8372 15436 8424
rect 26424 8415 26476 8424
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 8484 8236 8536 8288
rect 11796 8236 11848 8288
rect 12532 8236 12584 8288
rect 12624 8236 12676 8288
rect 17408 8304 17460 8356
rect 19616 8304 19668 8356
rect 16304 8236 16356 8288
rect 16580 8236 16632 8288
rect 18880 8279 18932 8288
rect 18880 8245 18889 8279
rect 18889 8245 18923 8279
rect 18923 8245 18932 8279
rect 18880 8236 18932 8245
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 2780 8032 2832 8084
rect 2872 8075 2924 8084
rect 2872 8041 2881 8075
rect 2881 8041 2915 8075
rect 2915 8041 2924 8075
rect 2872 8032 2924 8041
rect 3976 8032 4028 8084
rect 7288 8032 7340 8084
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 14188 8032 14240 8084
rect 14832 8075 14884 8084
rect 14832 8041 14841 8075
rect 14841 8041 14875 8075
rect 14875 8041 14884 8075
rect 14832 8032 14884 8041
rect 16396 8032 16448 8084
rect 18880 8032 18932 8084
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 7472 7964 7524 8016
rect 2320 7896 2372 7948
rect 3884 7896 3936 7948
rect 9036 7939 9088 7948
rect 9036 7905 9045 7939
rect 9045 7905 9079 7939
rect 9079 7905 9088 7939
rect 9036 7896 9088 7905
rect 11704 7896 11756 7948
rect 14004 7939 14056 7948
rect 14004 7905 14013 7939
rect 14013 7905 14047 7939
rect 14047 7905 14056 7939
rect 14004 7896 14056 7905
rect 16580 7896 16632 7948
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 1400 7828 1452 7880
rect 2688 7828 2740 7880
rect 6644 7828 6696 7880
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 12624 7803 12676 7812
rect 12624 7769 12633 7803
rect 12633 7769 12667 7803
rect 12667 7769 12676 7803
rect 12624 7760 12676 7769
rect 14832 7828 14884 7880
rect 16488 7871 16540 7880
rect 16488 7837 16497 7871
rect 16497 7837 16531 7871
rect 16531 7837 16540 7871
rect 16488 7828 16540 7837
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 4344 7735 4396 7744
rect 4344 7701 4353 7735
rect 4353 7701 4387 7735
rect 4387 7701 4396 7735
rect 4344 7692 4396 7701
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 8300 7692 8352 7744
rect 8760 7692 8812 7744
rect 11428 7692 11480 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 17868 7735 17920 7744
rect 17868 7701 17877 7735
rect 17877 7701 17911 7735
rect 17911 7701 17920 7735
rect 17868 7692 17920 7701
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 2320 7531 2372 7540
rect 2320 7497 2329 7531
rect 2329 7497 2363 7531
rect 2363 7497 2372 7531
rect 2320 7488 2372 7497
rect 5724 7488 5776 7540
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 7288 7488 7340 7540
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 9036 7488 9088 7540
rect 10140 7488 10192 7540
rect 8484 7420 8536 7472
rect 2872 7352 2924 7404
rect 3056 7395 3108 7404
rect 3056 7361 3065 7395
rect 3065 7361 3099 7395
rect 3099 7361 3108 7395
rect 3056 7352 3108 7361
rect 9496 7352 9548 7404
rect 14188 7488 14240 7540
rect 16580 7531 16632 7540
rect 16580 7497 16589 7531
rect 16589 7497 16623 7531
rect 16623 7497 16632 7531
rect 16580 7488 16632 7497
rect 19340 7488 19392 7540
rect 20168 7488 20220 7540
rect 22100 7488 22152 7540
rect 23204 7488 23256 7540
rect 26516 7488 26568 7540
rect 16488 7420 16540 7472
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 4344 7284 4396 7336
rect 11428 7352 11480 7404
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 13728 7395 13780 7404
rect 12808 7352 12860 7361
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 11888 7284 11940 7336
rect 13452 7284 13504 7336
rect 2320 7216 2372 7268
rect 3516 7259 3568 7268
rect 3516 7225 3525 7259
rect 3525 7225 3559 7259
rect 3559 7225 3568 7259
rect 3516 7216 3568 7225
rect 4712 7216 4764 7268
rect 11704 7259 11756 7268
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 9220 7148 9272 7200
rect 11704 7225 11713 7259
rect 11713 7225 11747 7259
rect 11747 7225 11756 7259
rect 11704 7216 11756 7225
rect 13544 7216 13596 7268
rect 10784 7148 10836 7200
rect 12992 7148 13044 7200
rect 13728 7148 13780 7200
rect 18880 7284 18932 7336
rect 14004 7216 14056 7268
rect 15108 7148 15160 7200
rect 26608 7191 26660 7200
rect 26608 7157 26617 7191
rect 26617 7157 26651 7191
rect 26651 7157 26660 7191
rect 26608 7148 26660 7157
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 2412 6944 2464 6996
rect 12348 6944 12400 6996
rect 13636 6944 13688 6996
rect 14004 6987 14056 6996
rect 14004 6953 14013 6987
rect 14013 6953 14047 6987
rect 14047 6953 14056 6987
rect 14004 6944 14056 6953
rect 2320 6919 2372 6928
rect 2320 6885 2329 6919
rect 2329 6885 2363 6919
rect 2363 6885 2372 6919
rect 2320 6876 2372 6885
rect 4344 6876 4396 6928
rect 1676 6808 1728 6860
rect 2688 6808 2740 6860
rect 3792 6808 3844 6860
rect 4620 6808 4672 6860
rect 5724 6876 5776 6928
rect 17868 6876 17920 6928
rect 6276 6808 6328 6860
rect 8300 6808 8352 6860
rect 10232 6808 10284 6860
rect 11428 6851 11480 6860
rect 11428 6817 11451 6851
rect 11451 6817 11480 6851
rect 11428 6808 11480 6817
rect 12992 6808 13044 6860
rect 18144 6851 18196 6860
rect 18144 6817 18178 6851
rect 18178 6817 18196 6851
rect 18144 6808 18196 6817
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 9312 6740 9364 6792
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 13452 6783 13504 6792
rect 2596 6672 2648 6724
rect 4252 6715 4304 6724
rect 4252 6681 4261 6715
rect 4261 6681 4295 6715
rect 4295 6681 4304 6715
rect 4252 6672 4304 6681
rect 9680 6715 9732 6724
rect 9680 6681 9689 6715
rect 9689 6681 9723 6715
rect 9723 6681 9732 6715
rect 9680 6672 9732 6681
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 7196 6604 7248 6656
rect 7380 6604 7432 6656
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 17868 6783 17920 6792
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 12532 6715 12584 6724
rect 12532 6681 12541 6715
rect 12541 6681 12575 6715
rect 12575 6681 12584 6715
rect 12532 6672 12584 6681
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 11520 6604 11572 6656
rect 12900 6647 12952 6656
rect 12900 6613 12909 6647
rect 12909 6613 12943 6647
rect 12943 6613 12952 6647
rect 12900 6604 12952 6613
rect 15200 6604 15252 6656
rect 16488 6604 16540 6656
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 2688 6400 2740 6452
rect 3976 6400 4028 6452
rect 5724 6443 5776 6452
rect 5724 6409 5733 6443
rect 5733 6409 5767 6443
rect 5767 6409 5776 6443
rect 5724 6400 5776 6409
rect 9220 6400 9272 6452
rect 12348 6400 12400 6452
rect 15752 6443 15804 6452
rect 15752 6409 15761 6443
rect 15761 6409 15795 6443
rect 15795 6409 15804 6443
rect 15752 6400 15804 6409
rect 17868 6400 17920 6452
rect 3792 6375 3844 6384
rect 3792 6341 3801 6375
rect 3801 6341 3835 6375
rect 3835 6341 3844 6375
rect 3792 6332 3844 6341
rect 4620 6375 4672 6384
rect 4620 6341 4629 6375
rect 4629 6341 4663 6375
rect 4663 6341 4672 6375
rect 4620 6332 4672 6341
rect 10324 6332 10376 6384
rect 2136 6264 2188 6316
rect 9864 6264 9916 6316
rect 2412 6239 2464 6248
rect 2412 6205 2421 6239
rect 2421 6205 2455 6239
rect 2455 6205 2464 6239
rect 2412 6196 2464 6205
rect 3976 6196 4028 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 11336 6196 11388 6248
rect 16212 6264 16264 6316
rect 16488 6307 16540 6316
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 13728 6239 13780 6248
rect 13728 6205 13762 6239
rect 13762 6205 13780 6239
rect 13728 6196 13780 6205
rect 15752 6196 15804 6248
rect 26516 6239 26568 6248
rect 26516 6205 26525 6239
rect 26525 6205 26559 6239
rect 26559 6205 26568 6239
rect 26516 6196 26568 6205
rect 13544 6128 13596 6180
rect 16396 6171 16448 6180
rect 16396 6137 16405 6171
rect 16405 6137 16439 6171
rect 16439 6137 16448 6171
rect 16396 6128 16448 6137
rect 1492 6060 1544 6112
rect 2412 6060 2464 6112
rect 6276 6060 6328 6112
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 10140 6060 10192 6112
rect 10416 6060 10468 6112
rect 11520 6060 11572 6112
rect 13360 6060 13412 6112
rect 15108 6060 15160 6112
rect 15844 6060 15896 6112
rect 18236 6103 18288 6112
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 2780 5899 2832 5908
rect 2780 5865 2789 5899
rect 2789 5865 2823 5899
rect 2823 5865 2832 5899
rect 2780 5856 2832 5865
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 10324 5856 10376 5908
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 13544 5899 13596 5908
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 14280 5899 14332 5908
rect 13544 5856 13596 5865
rect 14280 5865 14289 5899
rect 14289 5865 14323 5899
rect 14323 5865 14332 5899
rect 14280 5856 14332 5865
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 26700 5899 26752 5908
rect 26700 5865 26709 5899
rect 26709 5865 26743 5899
rect 26743 5865 26752 5899
rect 26700 5856 26752 5865
rect 10140 5788 10192 5840
rect 3608 5720 3660 5772
rect 4988 5720 5040 5772
rect 14372 5720 14424 5772
rect 16488 5720 16540 5772
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3884 5695 3936 5704
rect 3884 5661 3893 5695
rect 3893 5661 3927 5695
rect 3927 5661 3936 5695
rect 3884 5652 3936 5661
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 15568 5652 15620 5704
rect 16212 5652 16264 5704
rect 17500 5652 17552 5704
rect 15292 5584 15344 5636
rect 16672 5584 16724 5636
rect 17684 5584 17736 5636
rect 18236 5652 18288 5704
rect 6276 5516 6328 5568
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 15752 5559 15804 5568
rect 15752 5525 15761 5559
rect 15761 5525 15795 5559
rect 15795 5525 15804 5559
rect 15752 5516 15804 5525
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 2044 5355 2096 5364
rect 2044 5321 2053 5355
rect 2053 5321 2087 5355
rect 2087 5321 2096 5355
rect 2044 5312 2096 5321
rect 3884 5355 3936 5364
rect 3884 5321 3893 5355
rect 3893 5321 3927 5355
rect 3927 5321 3936 5355
rect 3884 5312 3936 5321
rect 4988 5355 5040 5364
rect 4988 5321 4997 5355
rect 4997 5321 5031 5355
rect 5031 5321 5040 5355
rect 4988 5312 5040 5321
rect 13360 5312 13412 5364
rect 15568 5355 15620 5364
rect 15568 5321 15577 5355
rect 15577 5321 15611 5355
rect 15611 5321 15620 5355
rect 15568 5312 15620 5321
rect 16396 5355 16448 5364
rect 16396 5321 16405 5355
rect 16405 5321 16439 5355
rect 16439 5321 16448 5355
rect 16396 5312 16448 5321
rect 18052 5355 18104 5364
rect 18052 5321 18061 5355
rect 18061 5321 18095 5355
rect 18095 5321 18104 5355
rect 18052 5312 18104 5321
rect 25872 5312 25924 5364
rect 26608 5355 26660 5364
rect 1400 5244 1452 5296
rect 1584 5244 1636 5296
rect 2044 5108 2096 5160
rect 2504 5151 2556 5160
rect 2504 5117 2513 5151
rect 2513 5117 2547 5151
rect 2547 5117 2556 5151
rect 2504 5108 2556 5117
rect 2780 5108 2832 5160
rect 4252 5151 4304 5160
rect 4252 5117 4261 5151
rect 4261 5117 4295 5151
rect 4295 5117 4304 5151
rect 4252 5108 4304 5117
rect 13360 5151 13412 5160
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 17684 5176 17736 5228
rect 16764 5151 16816 5160
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 18420 5151 18472 5160
rect 18420 5117 18429 5151
rect 18429 5117 18463 5151
rect 18463 5117 18472 5151
rect 18420 5108 18472 5117
rect 26608 5321 26617 5355
rect 26617 5321 26651 5355
rect 26651 5321 26660 5355
rect 26608 5312 26660 5321
rect 26516 5244 26568 5296
rect 5816 5040 5868 5092
rect 18512 5083 18564 5092
rect 18512 5049 18521 5083
rect 18521 5049 18555 5083
rect 18555 5049 18564 5083
rect 18512 5040 18564 5049
rect 1400 4972 1452 5024
rect 2688 5015 2740 5024
rect 2688 4981 2697 5015
rect 2697 4981 2731 5015
rect 2731 4981 2740 5015
rect 2688 4972 2740 4981
rect 2964 4972 3016 5024
rect 4344 5015 4396 5024
rect 4344 4981 4353 5015
rect 4353 4981 4387 5015
rect 4387 4981 4396 5015
rect 4344 4972 4396 4981
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 14740 5015 14792 5024
rect 14740 4981 14749 5015
rect 14749 4981 14783 5015
rect 14783 4981 14792 5015
rect 14740 4972 14792 4981
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16856 5015 16908 5024
rect 16304 4972 16356 4981
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 17500 5015 17552 5024
rect 17500 4981 17509 5015
rect 17509 4981 17543 5015
rect 17543 4981 17552 5015
rect 17500 4972 17552 4981
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 2596 4768 2648 4820
rect 2964 4768 3016 4820
rect 5724 4768 5776 4820
rect 12900 4768 12952 4820
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 14372 4811 14424 4820
rect 14372 4777 14381 4811
rect 14381 4777 14415 4811
rect 14415 4777 14424 4811
rect 14372 4768 14424 4777
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 16764 4768 16816 4820
rect 17684 4811 17736 4820
rect 17684 4777 17693 4811
rect 17693 4777 17727 4811
rect 17727 4777 17736 4811
rect 17684 4768 17736 4777
rect 18420 4768 18472 4820
rect 26700 4811 26752 4820
rect 26700 4777 26709 4811
rect 26709 4777 26743 4811
rect 26743 4777 26752 4811
rect 26700 4768 26752 4777
rect 3056 4743 3108 4752
rect 3056 4709 3065 4743
rect 3065 4709 3099 4743
rect 3099 4709 3108 4743
rect 3056 4700 3108 4709
rect 15844 4700 15896 4752
rect 17592 4700 17644 4752
rect 1584 4632 1636 4684
rect 1860 4632 1912 4684
rect 2872 4632 2924 4684
rect 3976 4632 4028 4684
rect 5816 4632 5868 4684
rect 13084 4632 13136 4684
rect 26516 4675 26568 4684
rect 26516 4641 26525 4675
rect 26525 4641 26559 4675
rect 26559 4641 26568 4675
rect 26516 4632 26568 4641
rect 4068 4564 4120 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 5724 4564 5776 4616
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 1676 4428 1728 4480
rect 12716 4564 12768 4616
rect 15384 4564 15436 4616
rect 6276 4428 6328 4480
rect 12348 4471 12400 4480
rect 12348 4437 12357 4471
rect 12357 4437 12391 4471
rect 12391 4437 12400 4471
rect 12348 4428 12400 4437
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 3976 4267 4028 4276
rect 3976 4233 3985 4267
rect 3985 4233 4019 4267
rect 4019 4233 4028 4267
rect 3976 4224 4028 4233
rect 5724 4224 5776 4276
rect 12900 4224 12952 4276
rect 13084 4267 13136 4276
rect 13084 4233 13093 4267
rect 13093 4233 13127 4267
rect 13127 4233 13136 4267
rect 13084 4224 13136 4233
rect 15384 4267 15436 4276
rect 15384 4233 15393 4267
rect 15393 4233 15427 4267
rect 15427 4233 15436 4267
rect 15384 4224 15436 4233
rect 15752 4224 15804 4276
rect 26516 4224 26568 4276
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 3424 4131 3476 4140
rect 3424 4097 3433 4131
rect 3433 4097 3467 4131
rect 3467 4097 3476 4131
rect 4620 4131 4672 4140
rect 3424 4088 3476 4097
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 5816 4088 5868 4140
rect 15844 4156 15896 4208
rect 8484 4063 8536 4072
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 8484 4020 8536 4029
rect 16488 4020 16540 4072
rect 26332 4020 26384 4072
rect 2872 3952 2924 4004
rect 4528 3952 4580 4004
rect 5632 3952 5684 4004
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 2780 3884 2832 3936
rect 3700 3884 3752 3936
rect 4436 3927 4488 3936
rect 4436 3893 4445 3927
rect 4445 3893 4479 3927
rect 4479 3893 4488 3927
rect 4436 3884 4488 3893
rect 6276 3927 6328 3936
rect 6276 3893 6285 3927
rect 6285 3893 6319 3927
rect 6319 3893 6328 3927
rect 6276 3884 6328 3893
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 26608 3927 26660 3936
rect 26608 3893 26617 3927
rect 26617 3893 26651 3927
rect 26651 3893 26660 3927
rect 26608 3884 26660 3893
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 1860 3680 1912 3732
rect 3240 3680 3292 3732
rect 4068 3723 4120 3732
rect 4068 3689 4077 3723
rect 4077 3689 4111 3723
rect 4111 3689 4120 3723
rect 4068 3680 4120 3689
rect 4528 3680 4580 3732
rect 13360 3680 13412 3732
rect 14096 3680 14148 3732
rect 14924 3723 14976 3732
rect 14924 3689 14933 3723
rect 14933 3689 14967 3723
rect 14967 3689 14976 3723
rect 14924 3680 14976 3689
rect 26700 3723 26752 3732
rect 26700 3689 26709 3723
rect 26709 3689 26743 3723
rect 26743 3689 26752 3723
rect 26700 3680 26752 3689
rect 8484 3612 8536 3664
rect 2228 3544 2280 3596
rect 2688 3544 2740 3596
rect 4804 3544 4856 3596
rect 9956 3544 10008 3596
rect 11520 3612 11572 3664
rect 11152 3544 11204 3596
rect 14464 3544 14516 3596
rect 16488 3544 16540 3596
rect 25320 3587 25372 3596
rect 25320 3553 25329 3587
rect 25329 3553 25363 3587
rect 25363 3553 25372 3587
rect 25320 3544 25372 3553
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 25044 3476 25096 3528
rect 27344 3476 27396 3528
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 4344 3340 4396 3392
rect 11796 3340 11848 3392
rect 12440 3383 12492 3392
rect 12440 3349 12449 3383
rect 12449 3349 12483 3383
rect 12483 3349 12492 3383
rect 12440 3340 12492 3349
rect 15844 3340 15896 3392
rect 25504 3383 25556 3392
rect 25504 3349 25513 3383
rect 25513 3349 25547 3383
rect 25547 3349 25556 3383
rect 25504 3340 25556 3349
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 2596 3179 2648 3188
rect 2596 3145 2605 3179
rect 2605 3145 2639 3179
rect 2639 3145 2648 3179
rect 2596 3136 2648 3145
rect 4620 3136 4672 3188
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 4528 3068 4580 3120
rect 5724 3068 5776 3120
rect 1492 2932 1544 2984
rect 2044 2932 2096 2984
rect 3240 3000 3292 3052
rect 3516 2932 3568 2984
rect 5264 2932 5316 2984
rect 6552 3136 6604 3188
rect 9956 3179 10008 3188
rect 9956 3145 9965 3179
rect 9965 3145 9999 3179
rect 9999 3145 10008 3179
rect 9956 3136 10008 3145
rect 12440 3136 12492 3188
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 25136 3179 25188 3188
rect 25136 3145 25145 3179
rect 25145 3145 25179 3179
rect 25179 3145 25188 3179
rect 25136 3136 25188 3145
rect 25320 3136 25372 3188
rect 26608 3179 26660 3188
rect 26608 3145 26617 3179
rect 26617 3145 26651 3179
rect 26651 3145 26660 3179
rect 26608 3136 26660 3145
rect 27344 3179 27396 3188
rect 27344 3145 27353 3179
rect 27353 3145 27387 3179
rect 27387 3145 27396 3179
rect 27344 3136 27396 3145
rect 8484 3000 8536 3052
rect 11152 3000 11204 3052
rect 12348 3000 12400 3052
rect 12716 2975 12768 2984
rect 12716 2941 12750 2975
rect 12750 2941 12768 2975
rect 14740 2975 14792 2984
rect 480 2864 532 2916
rect 4528 2864 4580 2916
rect 5540 2864 5592 2916
rect 8300 2796 8352 2848
rect 11152 2864 11204 2916
rect 12716 2932 12768 2941
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 14924 2975 14976 2984
rect 14924 2941 14933 2975
rect 14933 2941 14967 2975
rect 14967 2941 14976 2975
rect 14924 2932 14976 2941
rect 17960 2932 18012 2984
rect 25136 2932 25188 2984
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 27528 2975 27580 2984
rect 27528 2941 27537 2975
rect 27537 2941 27571 2975
rect 27571 2941 27580 2975
rect 27528 2932 27580 2941
rect 12624 2864 12676 2916
rect 15200 2907 15252 2916
rect 15200 2873 15212 2907
rect 15212 2873 15252 2907
rect 15200 2864 15252 2873
rect 12808 2796 12860 2848
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 15292 2796 15344 2848
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 25504 2839 25556 2848
rect 25504 2805 25513 2839
rect 25513 2805 25547 2839
rect 25547 2805 25556 2839
rect 25504 2796 25556 2805
rect 27712 2839 27764 2848
rect 27712 2805 27721 2839
rect 27721 2805 27755 2839
rect 27755 2805 27764 2839
rect 27712 2796 27764 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 2044 2592 2096 2644
rect 2412 2592 2464 2644
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 11612 2635 11664 2644
rect 11612 2601 11621 2635
rect 11621 2601 11655 2635
rect 11655 2601 11664 2635
rect 11612 2592 11664 2601
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12072 2592 12124 2601
rect 12440 2592 12492 2644
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 14464 2635 14516 2644
rect 14464 2601 14473 2635
rect 14473 2601 14507 2635
rect 14507 2601 14516 2635
rect 14464 2592 14516 2601
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 4344 2524 4396 2576
rect 6276 2567 6328 2576
rect 6276 2533 6285 2567
rect 6285 2533 6319 2567
rect 6319 2533 6328 2567
rect 6276 2524 6328 2533
rect 8208 2524 8260 2576
rect 11520 2524 11572 2576
rect 4620 2499 4672 2508
rect 4620 2465 4654 2499
rect 4654 2465 4672 2499
rect 4620 2456 4672 2465
rect 16580 2592 16632 2644
rect 19616 2635 19668 2644
rect 19616 2601 19625 2635
rect 19625 2601 19659 2635
rect 19659 2601 19668 2635
rect 19616 2592 19668 2601
rect 23020 2635 23072 2644
rect 23020 2601 23029 2635
rect 23029 2601 23063 2635
rect 23063 2601 23072 2635
rect 23020 2592 23072 2601
rect 27068 2635 27120 2644
rect 27068 2601 27077 2635
rect 27077 2601 27111 2635
rect 27111 2601 27120 2635
rect 27068 2592 27120 2601
rect 14280 2499 14332 2508
rect 2504 2388 2556 2440
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 14924 2456 14976 2508
rect 18420 2456 18472 2508
rect 19432 2499 19484 2508
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 22836 2499 22888 2508
rect 22836 2465 22845 2499
rect 22845 2465 22879 2499
rect 22879 2465 22888 2499
rect 22836 2456 22888 2465
rect 24584 2499 24636 2508
rect 24584 2465 24593 2499
rect 24593 2465 24627 2499
rect 24627 2465 24636 2499
rect 24584 2456 24636 2465
rect 25688 2499 25740 2508
rect 25688 2465 25697 2499
rect 25697 2465 25731 2499
rect 25731 2465 25740 2499
rect 25688 2456 25740 2465
rect 26792 2456 26844 2508
rect 15108 2388 15160 2440
rect 14924 2320 14976 2372
rect 2964 2295 3016 2304
rect 2964 2261 2973 2295
rect 2973 2261 3007 2295
rect 3007 2261 3016 2295
rect 2964 2252 3016 2261
rect 7840 2252 7892 2304
rect 8576 2295 8628 2304
rect 8576 2261 8585 2295
rect 8585 2261 8619 2295
rect 8619 2261 8628 2295
rect 8576 2252 8628 2261
rect 10784 2252 10836 2304
rect 18512 2295 18564 2304
rect 18512 2261 18521 2295
rect 18521 2261 18555 2295
rect 18555 2261 18564 2295
rect 18512 2252 18564 2261
rect 24768 2295 24820 2304
rect 24768 2261 24777 2295
rect 24777 2261 24811 2295
rect 24811 2261 24820 2295
rect 24768 2252 24820 2261
rect 25872 2295 25924 2304
rect 25872 2261 25881 2295
rect 25881 2261 25915 2295
rect 25915 2261 25924 2295
rect 25872 2252 25924 2261
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
rect 19064 552 19116 604
rect 19156 552 19208 604
<< metal2 >>
rect 754 23520 810 24000
rect 2226 23520 2282 24000
rect 2962 23624 3018 23633
rect 2962 23559 3018 23568
rect 768 20369 796 23520
rect 754 20360 810 20369
rect 754 20295 810 20304
rect 2240 19825 2268 23520
rect 2778 23080 2834 23089
rect 2778 23015 2834 23024
rect 2226 19816 2282 19825
rect 2226 19751 2282 19760
rect 2792 19530 2820 23015
rect 2976 22234 3004 23559
rect 3698 23520 3754 24000
rect 5170 23520 5226 24000
rect 6734 23520 6790 24000
rect 8206 23520 8262 24000
rect 9678 23520 9734 24000
rect 11242 23520 11298 24000
rect 12714 23520 12770 24000
rect 14186 23520 14242 24000
rect 15750 23520 15806 24000
rect 17222 23520 17278 24000
rect 18694 23520 18750 24000
rect 20166 23520 20222 24000
rect 21730 23520 21786 24000
rect 23202 23520 23258 24000
rect 24674 23520 24730 24000
rect 25502 23624 25558 23633
rect 25502 23559 25558 23568
rect 2964 22228 3016 22234
rect 2964 22170 3016 22176
rect 3148 20936 3200 20942
rect 3148 20878 3200 20884
rect 2792 19502 2912 19530
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 2318 14648 2374 14657
rect 2318 14583 2374 14592
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1688 13530 1716 13670
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1490 13288 1546 13297
rect 1490 13223 1546 13232
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1412 9722 1440 10066
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1412 7886 1440 8978
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1504 6848 1532 13223
rect 1688 12782 1716 13466
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12850 1900 13126
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1872 12442 1900 12786
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 2056 12374 2084 12786
rect 2044 12368 2096 12374
rect 2042 12336 2044 12345
rect 2096 12336 2098 12345
rect 2042 12271 2098 12280
rect 1582 11656 1638 11665
rect 1582 11591 1638 11600
rect 1596 11558 1624 11591
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1582 11112 1638 11121
rect 1582 11047 1638 11056
rect 1596 10810 1624 11047
rect 2042 10840 2098 10849
rect 1584 10804 1636 10810
rect 2042 10775 2044 10784
rect 1584 10746 1636 10752
rect 2096 10775 2098 10784
rect 2044 10746 2096 10752
rect 2056 10606 2084 10746
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 1582 10432 1638 10441
rect 1582 10367 1638 10376
rect 1596 10266 1624 10367
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 2332 9926 2360 14583
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2516 11898 2544 13466
rect 2700 13394 2728 13806
rect 2792 13530 2820 19343
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2884 13410 2912 19502
rect 2962 15328 3018 15337
rect 2962 15263 3018 15272
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2792 13382 2912 13410
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2516 11558 2544 11834
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2424 10810 2452 11018
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2502 10568 2558 10577
rect 2502 10503 2558 10512
rect 2320 9920 2372 9926
rect 1582 9888 1638 9897
rect 2320 9862 2372 9868
rect 1582 9823 1638 9832
rect 1596 9654 1624 9823
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1582 9344 1638 9353
rect 1582 9279 1638 9288
rect 1596 9178 1624 9279
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 2516 9042 2544 10503
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 1582 8664 1638 8673
rect 2516 8634 2544 8978
rect 1582 8599 1584 8608
rect 1636 8599 1638 8608
rect 2504 8628 2556 8634
rect 1584 8570 1636 8576
rect 2504 8570 2556 8576
rect 2042 8528 2098 8537
rect 2042 8463 2044 8472
rect 2096 8463 2098 8472
rect 2044 8434 2096 8440
rect 1950 8256 2006 8265
rect 1950 8191 2006 8200
rect 1412 6820 1532 6848
rect 1676 6860 1728 6866
rect 1412 5302 1440 6820
rect 1676 6802 1728 6808
rect 1584 6656 1636 6662
rect 1688 6633 1716 6802
rect 1584 6598 1636 6604
rect 1674 6624 1730 6633
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1400 5296 1452 5302
rect 1400 5238 1452 5244
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 480 2916 532 2922
rect 480 2858 532 2864
rect 492 480 520 2858
rect 1412 921 1440 4966
rect 1504 2990 1532 6054
rect 1596 5681 1624 6598
rect 1674 6559 1730 6568
rect 1688 6458 1716 6559
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1584 5296 1636 5302
rect 1584 5238 1636 5244
rect 1596 4690 1624 5238
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1584 4480 1636 4486
rect 1582 4448 1584 4457
rect 1676 4480 1728 4486
rect 1636 4448 1638 4457
rect 1676 4422 1728 4428
rect 1582 4383 1638 4392
rect 1584 3936 1636 3942
rect 1582 3904 1584 3913
rect 1636 3904 1638 3913
rect 1582 3839 1638 3848
rect 1584 3392 1636 3398
rect 1582 3360 1584 3369
rect 1636 3360 1638 3369
rect 1582 3295 1638 3304
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1490 2816 1546 2825
rect 1490 2751 1546 2760
rect 1398 912 1454 921
rect 1398 847 1454 856
rect 1504 480 1532 2751
rect 478 0 534 480
rect 1490 0 1546 480
rect 1688 377 1716 4422
rect 1872 3738 1900 4626
rect 1964 4146 1992 8191
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2332 7546 2360 7890
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2424 7290 2452 7686
rect 2608 7562 2636 12854
rect 2792 12782 2820 13382
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2884 12986 2912 13262
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2792 11898 2820 12242
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2686 11792 2742 11801
rect 2686 11727 2688 11736
rect 2740 11727 2742 11736
rect 2688 11698 2740 11704
rect 2884 11354 2912 12174
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10810 2820 11154
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2792 10266 2820 10746
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2884 9994 2912 11086
rect 2976 10010 3004 15263
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3068 12238 3096 13262
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3054 12064 3110 12073
rect 3054 11999 3110 12008
rect 3068 10713 3096 11999
rect 3054 10704 3110 10713
rect 3054 10639 3110 10648
rect 2872 9988 2924 9994
rect 2976 9982 3096 10010
rect 2872 9930 2924 9936
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 8129 2728 8774
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2686 8120 2742 8129
rect 2792 8090 2820 8230
rect 2686 8055 2742 8064
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2688 7880 2740 7886
rect 2686 7848 2688 7857
rect 2740 7848 2742 7857
rect 2686 7783 2742 7792
rect 2332 7274 2452 7290
rect 2320 7268 2452 7274
rect 2372 7262 2452 7268
rect 2516 7534 2636 7562
rect 2320 7210 2372 7216
rect 2332 6934 2360 7210
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2424 7002 2452 7142
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2148 6225 2176 6258
rect 2424 6254 2452 6938
rect 2412 6248 2464 6254
rect 2134 6216 2190 6225
rect 2412 6190 2464 6196
rect 2516 6202 2544 7534
rect 2594 7440 2650 7449
rect 2594 7375 2650 7384
rect 2608 6730 2636 7375
rect 2792 7342 2820 8026
rect 2884 7410 2912 8026
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2700 6458 2728 6802
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2516 6174 2636 6202
rect 2134 6151 2190 6160
rect 2042 5944 2098 5953
rect 2148 5914 2176 6151
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5914 2452 6054
rect 2042 5879 2098 5888
rect 2136 5908 2188 5914
rect 2056 5370 2084 5879
rect 2136 5850 2188 5856
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2608 5794 2636 6174
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2424 5766 2636 5794
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2056 5166 2084 5306
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2226 4992 2282 5001
rect 2226 4927 2282 4936
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2240 3602 2268 4927
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2240 3194 2268 3538
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2056 2650 2084 2926
rect 2424 2650 2452 5766
rect 2792 5658 2820 5850
rect 2608 5630 2820 5658
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2502 5264 2558 5273
rect 2502 5199 2558 5208
rect 2516 5166 2544 5199
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2608 4826 2636 5630
rect 2780 5160 2832 5166
rect 2686 5128 2742 5137
rect 2780 5102 2832 5108
rect 2686 5063 2742 5072
rect 2700 5030 2728 5063
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2792 4162 2820 5102
rect 2884 4808 2912 5646
rect 2976 5030 3004 9862
rect 3068 7528 3096 9982
rect 3160 9654 3188 20878
rect 3712 19961 3740 23520
rect 4066 22400 4122 22409
rect 4066 22335 4068 22344
rect 4120 22335 4122 22344
rect 4068 22306 4120 22312
rect 3974 21856 4030 21865
rect 3974 21791 4030 21800
rect 3882 21312 3938 21321
rect 3882 21247 3938 21256
rect 3896 21010 3924 21247
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 3882 20632 3938 20641
rect 3882 20567 3938 20576
rect 3698 19952 3754 19961
rect 3698 19887 3754 19896
rect 3422 18320 3478 18329
rect 3422 18255 3478 18264
rect 3698 18320 3754 18329
rect 3698 18255 3754 18264
rect 3238 14104 3294 14113
rect 3238 14039 3294 14048
rect 3252 11665 3280 14039
rect 3332 12776 3384 12782
rect 3330 12744 3332 12753
rect 3384 12744 3386 12753
rect 3330 12679 3386 12688
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 12481 3372 12582
rect 3330 12472 3386 12481
rect 3330 12407 3386 12416
rect 3238 11656 3294 11665
rect 3436 11642 3464 18255
rect 3514 14920 3570 14929
rect 3514 14855 3570 14864
rect 3528 12986 3556 14855
rect 3712 13512 3740 18255
rect 3896 15065 3924 20567
rect 3882 15056 3938 15065
rect 3882 14991 3938 15000
rect 3712 13484 3832 13512
rect 3698 13424 3754 13433
rect 3698 13359 3754 13368
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3514 12880 3570 12889
rect 3514 12815 3570 12824
rect 3608 12844 3660 12850
rect 3528 12209 3556 12815
rect 3608 12786 3660 12792
rect 3620 12442 3648 12786
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3514 12200 3570 12209
rect 3514 12135 3570 12144
rect 3620 11898 3648 12378
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3238 11591 3294 11600
rect 3332 11620 3384 11626
rect 3436 11614 3556 11642
rect 3332 11562 3384 11568
rect 3238 11112 3294 11121
rect 3238 11047 3294 11056
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3160 9178 3188 9590
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3160 8498 3188 9114
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3068 7500 3188 7528
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3068 6662 3096 7346
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 5710 3096 6598
rect 3160 6089 3188 7500
rect 3146 6080 3202 6089
rect 3146 6015 3202 6024
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2964 4820 3016 4826
rect 2884 4780 2964 4808
rect 2964 4762 3016 4768
rect 3068 4758 3096 5646
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2700 4134 2820 4162
rect 2700 3602 2728 4134
rect 2884 4010 2912 4626
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2700 3482 2728 3538
rect 2608 3454 2728 3482
rect 2608 3194 2636 3454
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2700 2689 2728 3334
rect 2686 2680 2742 2689
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2412 2644 2464 2650
rect 2686 2615 2742 2624
rect 2412 2586 2464 2592
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 2516 480 2544 2382
rect 2792 1465 2820 3878
rect 3252 3738 3280 11047
rect 3344 8129 3372 11562
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3436 11354 3464 11494
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3528 10962 3556 11614
rect 3620 11150 3648 11834
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3528 10934 3648 10962
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10305 3464 10406
rect 3422 10296 3478 10305
rect 3422 10231 3424 10240
rect 3476 10231 3478 10240
rect 3424 10202 3476 10208
rect 3330 8120 3386 8129
rect 3330 8055 3386 8064
rect 3330 7032 3386 7041
rect 3330 6967 3386 6976
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3252 3058 3280 3674
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3344 2650 3372 6967
rect 3436 4146 3464 10202
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3528 7750 3556 8434
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7274 3556 7686
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3620 5778 3648 10934
rect 3712 10470 3740 13359
rect 3804 12617 3832 13484
rect 3988 12730 4016 21791
rect 5184 20806 5212 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 6748 20505 6776 23520
rect 8220 20874 8248 23520
rect 8208 20868 8260 20874
rect 8208 20810 8260 20816
rect 9692 20618 9720 23520
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 9600 20602 9720 20618
rect 9588 20596 9720 20602
rect 9640 20590 9720 20596
rect 9588 20538 9640 20544
rect 6734 20496 6790 20505
rect 6734 20431 6790 20440
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 4066 20088 4122 20097
rect 4066 20023 4122 20032
rect 4080 14521 4108 20023
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 7838 16960 7894 16969
rect 7838 16895 7894 16904
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 4618 16008 4674 16017
rect 4618 15943 4674 15952
rect 4342 15872 4398 15881
rect 4342 15807 4398 15816
rect 4066 14512 4122 14521
rect 4066 14447 4122 14456
rect 3988 12702 4200 12730
rect 4068 12640 4120 12646
rect 3790 12608 3846 12617
rect 3790 12543 3846 12552
rect 3974 12608 4030 12617
rect 4068 12582 4120 12588
rect 3974 12543 4030 12552
rect 3790 12472 3846 12481
rect 3790 12407 3846 12416
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3712 3942 3740 10406
rect 3804 6866 3832 12407
rect 3882 8936 3938 8945
rect 3882 8871 3938 8880
rect 3896 7954 3924 8871
rect 3988 8090 4016 12543
rect 4080 12238 4108 12582
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4080 11898 4108 12174
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4172 11778 4200 12702
rect 4080 11750 4200 11778
rect 4080 8945 4108 11750
rect 4356 11150 4384 15807
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4540 12986 4568 13330
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4436 12708 4488 12714
rect 4436 12650 4488 12656
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4448 10849 4476 12650
rect 4540 12442 4568 12718
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4632 11218 4660 15943
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4908 12782 4936 13670
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 5000 12442 5028 13262
rect 5078 12880 5134 12889
rect 5276 12850 5304 13330
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 5078 12815 5134 12824
rect 5264 12844 5316 12850
rect 5092 12782 5120 12815
rect 5264 12786 5316 12792
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 6380 12374 6408 13126
rect 7668 12850 7696 13262
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 6828 12640 6880 12646
rect 7196 12640 7248 12646
rect 6880 12588 6960 12594
rect 6828 12582 6960 12588
rect 7196 12582 7248 12588
rect 6840 12566 6960 12582
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5828 11830 5856 12242
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 6380 11898 6408 12310
rect 6734 12064 6790 12073
rect 6734 11999 6790 12008
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6748 11830 6776 11999
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6748 11218 6776 11766
rect 6932 11354 6960 12566
rect 7208 12442 7236 12582
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7208 12345 7236 12378
rect 7194 12336 7250 12345
rect 7194 12271 7250 12280
rect 7668 12073 7696 12786
rect 7654 12064 7710 12073
rect 7654 11999 7710 12008
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4434 10840 4490 10849
rect 4434 10775 4490 10784
rect 4540 10554 4568 11086
rect 4448 10526 4568 10554
rect 4448 10470 4476 10526
rect 4632 10470 4660 11154
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4802 10704 4858 10713
rect 4908 10674 4936 11086
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 6748 10792 6776 11154
rect 6920 10804 6972 10810
rect 6748 10764 6920 10792
rect 6920 10746 6972 10752
rect 4802 10639 4858 10648
rect 4896 10668 4948 10674
rect 4436 10464 4488 10470
rect 4620 10464 4672 10470
rect 4436 10406 4488 10412
rect 4526 10432 4582 10441
rect 4250 10160 4306 10169
rect 4250 10095 4306 10104
rect 4264 9722 4292 10095
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4066 8936 4122 8945
rect 4066 8871 4122 8880
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3988 6458 4016 8026
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4356 7342 4384 7686
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4356 6934 4384 7278
rect 4344 6928 4396 6934
rect 4250 6896 4306 6905
rect 4344 6870 4396 6876
rect 4250 6831 4306 6840
rect 4264 6730 4292 6831
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3792 6384 3844 6390
rect 3790 6352 3792 6361
rect 3844 6352 3846 6361
rect 3790 6287 3846 6296
rect 3988 6254 4016 6394
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3896 5370 3924 5646
rect 4250 5536 4306 5545
rect 4250 5471 4306 5480
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 4264 5166 4292 5471
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4356 4729 4384 4966
rect 4342 4720 4398 4729
rect 3976 4684 4028 4690
rect 4342 4655 4398 4664
rect 3976 4626 4028 4632
rect 3988 4282 4016 4626
rect 4068 4616 4120 4622
rect 4448 4593 4476 10406
rect 4620 10406 4672 10412
rect 4526 10367 4582 10376
rect 4540 10266 4568 10367
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4540 9722 4568 10202
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4068 4558 4120 4564
rect 4434 4584 4490 4593
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 4080 3738 4108 4558
rect 4434 4519 4490 4528
rect 4540 4010 4568 9658
rect 4632 8265 4660 10406
rect 4816 10130 4844 10639
rect 4896 10610 4948 10616
rect 4908 10470 4936 10610
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4816 9654 4844 10066
rect 4908 10062 4936 10406
rect 6932 10266 6960 10746
rect 7116 10470 7144 11222
rect 7562 10840 7618 10849
rect 7562 10775 7618 10784
rect 7576 10577 7604 10775
rect 7562 10568 7618 10577
rect 7562 10503 7618 10512
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6932 10146 6960 10202
rect 6840 10118 6960 10146
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 9722 4936 9998
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4618 8256 4674 8265
rect 4618 8191 4674 8200
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4632 6390 4660 6802
rect 4620 6384 4672 6390
rect 4618 6352 4620 6361
rect 4672 6352 4674 6361
rect 4618 6287 4674 6296
rect 4724 5710 4752 7210
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4724 4622 4752 5646
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4448 3641 4476 3878
rect 4540 3738 4568 3946
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4434 3632 4490 3641
rect 4434 3567 4490 3576
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2976 2145 3004 2246
rect 2962 2136 3018 2145
rect 2962 2071 3018 2080
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3528 480 3556 2926
rect 4356 2582 4384 3334
rect 4540 3126 4568 3674
rect 4632 3534 4660 4082
rect 4816 3602 4844 9590
rect 6840 9586 6868 10118
rect 7116 9722 7144 10406
rect 7852 9897 7880 16895
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7838 9888 7894 9897
rect 7838 9823 7894 9832
rect 7470 9752 7526 9761
rect 7104 9716 7156 9722
rect 7470 9687 7526 9696
rect 7104 9658 7156 9664
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6840 9110 6868 9522
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5828 8634 5856 8978
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 6288 8566 6316 9046
rect 7116 8838 7144 9386
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 7116 7886 7144 8774
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 8090 7328 8230
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5736 6934 5764 7482
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 5736 6458 5764 6870
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 6288 6118 6316 6802
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 4986 5808 5042 5817
rect 4986 5743 4988 5752
rect 5040 5743 5042 5752
rect 4988 5714 5040 5720
rect 5000 5370 5028 5714
rect 6288 5574 6316 6054
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4826 5764 4966
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5736 4622 5764 4762
rect 5828 4690 5856 5034
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5736 4282 5764 4558
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5828 4146 5856 4626
rect 6288 4486 6316 5510
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4632 3194 4660 3470
rect 4816 3194 4844 3538
rect 5262 3496 5318 3505
rect 5262 3431 5318 3440
rect 5276 3194 5304 3431
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 5276 2990 5304 3130
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4356 2446 4384 2518
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4540 480 4568 2858
rect 5552 2825 5580 2858
rect 5538 2816 5594 2825
rect 5538 2751 5594 2760
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4632 1601 4660 2450
rect 4618 1592 4674 1601
rect 4618 1527 4674 1536
rect 5644 480 5672 3946
rect 6288 3942 6316 4422
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5736 2650 5764 3062
rect 6288 2961 6316 3878
rect 6564 3194 6592 7686
rect 6656 7546 6684 7822
rect 7300 7546 7328 8026
rect 7484 8022 7512 9687
rect 8128 9654 8156 10202
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8220 10010 8248 10066
rect 8220 9982 8340 10010
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8312 9382 8340 9982
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 7930 8664 7986 8673
rect 7930 8599 7932 8608
rect 7984 8599 7986 8608
rect 7932 8570 7984 8576
rect 7944 8498 7972 8570
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7668 8090 7696 8366
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7484 7546 7512 7958
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 8312 6866 8340 7686
rect 8496 7478 8524 8230
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7208 6254 7236 6598
rect 7392 6254 7420 6598
rect 7196 6248 7248 6254
rect 7194 6216 7196 6225
rect 7380 6248 7432 6254
rect 7248 6216 7250 6225
rect 7380 6190 7432 6196
rect 7194 6151 7250 6160
rect 7392 5574 7420 6190
rect 8312 5914 8340 6802
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 8484 4072 8536 4078
rect 8482 4040 8484 4049
rect 8536 4040 8538 4049
rect 8482 3975 8538 3984
rect 8588 3913 8616 20334
rect 9218 18864 9274 18873
rect 9218 18799 9274 18808
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9048 11665 9076 12174
rect 9034 11656 9090 11665
rect 9034 11591 9036 11600
rect 9088 11591 9090 11600
rect 9036 11562 9088 11568
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8772 7750 8800 9318
rect 9232 8430 9260 18799
rect 9494 16552 9550 16561
rect 9494 16487 9550 16496
rect 9508 13462 9536 16487
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 12918 9996 13330
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9402 12200 9458 12209
rect 9402 12135 9458 12144
rect 9416 11898 9444 12135
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9588 11892 9640 11898
rect 9692 11880 9720 12786
rect 10152 12458 10180 12854
rect 10244 12850 10272 13670
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10152 12430 10272 12458
rect 10520 12442 10548 12582
rect 10244 12238 10272 12430
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 9640 11852 9720 11880
rect 9588 11834 9640 11840
rect 9416 11694 9444 11834
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9722 9720 9998
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 8838 9536 9386
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9508 8498 9536 8774
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9048 7857 9076 7890
rect 9034 7848 9090 7857
rect 9034 7783 9090 7792
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 9048 7546 9076 7783
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9232 7449 9260 8366
rect 9218 7440 9274 7449
rect 9508 7410 9536 8434
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9218 7375 9274 7384
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 8666 7304 8722 7313
rect 8666 7239 8722 7248
rect 8574 3904 8630 3913
rect 8574 3839 8630 3848
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 8496 3058 8524 3606
rect 8574 3088 8630 3097
rect 8484 3052 8536 3058
rect 8574 3023 8630 3032
rect 8484 2994 8536 3000
rect 8496 2961 8524 2994
rect 6274 2952 6330 2961
rect 6274 2887 6330 2896
rect 8482 2952 8538 2961
rect 8482 2887 8538 2896
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 6288 2582 6316 2887
rect 8300 2848 8352 2854
rect 8220 2796 8300 2802
rect 8220 2790 8352 2796
rect 8220 2774 8340 2790
rect 8220 2582 8248 2774
rect 6276 2576 6328 2582
rect 6276 2518 6328 2524
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8588 2310 8616 3023
rect 7840 2304 7892 2310
rect 7668 2252 7840 2258
rect 7668 2246 7892 2252
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 7668 2230 7880 2246
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 6642 1592 6698 1601
rect 6642 1527 6698 1536
rect 6656 480 6684 1527
rect 7668 480 7696 2230
rect 8680 480 8708 7239
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 6662 9260 7142
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 6458 9260 6598
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9324 6118 9352 6734
rect 9600 6712 9628 8298
rect 9784 8242 9812 11630
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11082 9996 11494
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9876 9450 9904 10134
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9968 8673 9996 10610
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 9761 10088 10406
rect 10046 9752 10102 9761
rect 10046 9687 10102 9696
rect 9954 8664 10010 8673
rect 9954 8599 10010 8608
rect 9784 8214 9904 8242
rect 9770 8120 9826 8129
rect 9770 8055 9826 8064
rect 9680 6724 9732 6730
rect 9600 6684 9680 6712
rect 9680 6666 9732 6672
rect 9784 6225 9812 8055
rect 9876 6322 9904 8214
rect 10152 7546 10180 12174
rect 10244 11762 10272 12174
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10244 11354 10272 11698
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9770 6216 9826 6225
rect 9770 6151 9826 6160
rect 9312 6112 9364 6118
rect 9310 6080 9312 6089
rect 10140 6112 10192 6118
rect 9364 6080 9366 6089
rect 10140 6054 10192 6060
rect 9310 6015 9366 6024
rect 9324 5681 9352 6015
rect 10152 5953 10180 6054
rect 10138 5944 10194 5953
rect 10138 5879 10194 5888
rect 10152 5846 10180 5879
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 9310 5672 9366 5681
rect 9310 5607 9366 5616
rect 10244 5574 10272 6802
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 6390 10364 6734
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 10336 5914 10364 6326
rect 10428 6118 10456 11018
rect 10612 9654 10640 21966
rect 11256 21434 11284 23520
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 11256 21406 11376 21434
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 11348 20602 11376 21406
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 12070 18864 12126 18873
rect 12070 18799 12126 18808
rect 11978 18048 12034 18057
rect 10956 17980 11252 18000
rect 11978 17983 12034 17992
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 11796 14544 11848 14550
rect 11794 14512 11796 14521
rect 11848 14512 11850 14521
rect 11794 14447 11850 14456
rect 11888 14476 11940 14482
rect 11808 14074 11836 14447
rect 11888 14418 11940 14424
rect 11900 14074 11928 14418
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10796 13190 10824 13738
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11900 13530 11928 14010
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11808 13297 11836 13330
rect 11794 13288 11850 13297
rect 11794 13223 11850 13232
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 12850 10824 13126
rect 11808 12986 11836 13223
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10796 12442 10824 12786
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10704 11558 10732 12242
rect 11440 11898 11468 12378
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10704 7970 10732 11494
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 11716 11121 11744 12038
rect 11702 11112 11758 11121
rect 11702 11047 11758 11056
rect 11992 10985 12020 17983
rect 11978 10976 12034 10985
rect 11978 10911 12034 10920
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 10796 9722 10824 10474
rect 10888 10266 10916 10610
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10888 9178 10916 9522
rect 11152 9512 11204 9518
rect 11150 9480 11152 9489
rect 11204 9480 11206 9489
rect 11150 9415 11206 9424
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 11348 9178 11376 10406
rect 11992 9722 12020 10911
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 10782 7984 10838 7993
rect 10704 7942 10782 7970
rect 10782 7919 10838 7928
rect 10796 7206 10824 7919
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10690 7032 10746 7041
rect 10796 7018 10824 7142
rect 10746 6990 10824 7018
rect 10690 6967 10746 6976
rect 10704 6798 10732 6967
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10888 6361 10916 9114
rect 11532 9042 11560 9658
rect 12084 9654 12112 18799
rect 12544 18193 12572 22102
rect 12728 20398 12756 23520
rect 13176 22228 13228 22234
rect 13176 22170 13228 22176
rect 13188 21978 13216 22170
rect 13188 21950 13308 21978
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12728 19417 12756 20198
rect 12714 19408 12770 19417
rect 12714 19343 12770 19352
rect 12530 18184 12586 18193
rect 12530 18119 12586 18128
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12176 13938 12204 14350
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12268 12986 12296 13398
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12452 12782 12480 14214
rect 12898 13424 12954 13433
rect 12898 13359 12900 13368
rect 12952 13359 12954 13368
rect 12900 13330 12952 13336
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12728 12918 12756 13262
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12442 12480 12582
rect 12912 12442 12940 12786
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13096 12442 13124 12718
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12360 11830 12388 12174
rect 12452 11898 12480 12242
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12348 11824 12400 11830
rect 12346 11792 12348 11801
rect 12400 11792 12402 11801
rect 12346 11727 12402 11736
rect 12360 11701 12388 11727
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11286 12204 11630
rect 12452 11354 12480 11834
rect 12820 11694 12848 12038
rect 12912 11762 12940 12378
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12912 11354 12940 11494
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 13096 10674 13124 11494
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11532 8566 11560 8978
rect 11624 8634 11652 9114
rect 11808 8974 11836 9522
rect 12176 9178 12204 9998
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 13188 9081 13216 20946
rect 13280 11218 13308 21950
rect 14200 21298 14228 23520
rect 14200 21270 14320 21298
rect 14188 21072 14240 21078
rect 14188 21014 14240 21020
rect 13450 17776 13506 17785
rect 13450 17711 13506 17720
rect 13464 13002 13492 17711
rect 14002 14376 14058 14385
rect 14002 14311 14058 14320
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13648 13190 13676 13806
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13464 12974 13676 13002
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13556 11937 13584 12242
rect 13542 11928 13598 11937
rect 13542 11863 13598 11872
rect 13452 11688 13504 11694
rect 13556 11665 13584 11863
rect 13452 11630 13504 11636
rect 13542 11656 13598 11665
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13280 11121 13308 11154
rect 13464 11150 13492 11630
rect 13542 11591 13544 11600
rect 13596 11591 13598 11600
rect 13544 11562 13596 11568
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13452 11144 13504 11150
rect 13266 11112 13322 11121
rect 13452 11086 13504 11092
rect 13266 11047 13322 11056
rect 13280 10810 13308 11047
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13464 10266 13492 11086
rect 13556 10849 13584 11290
rect 13542 10840 13598 10849
rect 13542 10775 13544 10784
rect 13596 10775 13598 10784
rect 13544 10746 13596 10752
rect 13556 10715 13584 10746
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13174 9072 13230 9081
rect 13174 9007 13230 9016
rect 13542 9072 13598 9081
rect 13542 9007 13598 9016
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11808 8294 11836 8910
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11440 7410 11468 7686
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 11440 6866 11468 7346
rect 11716 7313 11744 7890
rect 11888 7336 11940 7342
rect 11702 7304 11758 7313
rect 11888 7278 11940 7284
rect 11702 7239 11704 7248
rect 11756 7239 11758 7248
rect 11704 7210 11756 7216
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 10874 6352 10930 6361
rect 10874 6287 10930 6296
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 10416 6112 10468 6118
rect 11348 6089 11376 6190
rect 11532 6118 11560 6598
rect 11520 6112 11572 6118
rect 10416 6054 10468 6060
rect 11334 6080 11390 6089
rect 10956 6012 11252 6032
rect 11520 6054 11572 6060
rect 11334 6015 11390 6024
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 5273 10272 5510
rect 10230 5264 10286 5273
rect 10230 5199 10286 5208
rect 10244 5001 10272 5199
rect 10230 4992 10286 5001
rect 10230 4927 10286 4936
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 9770 3904 9826 3913
rect 9770 3839 9826 3848
rect 9784 480 9812 3839
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 11532 3670 11560 6054
rect 11900 5001 11928 7278
rect 11886 4992 11942 5001
rect 11886 4927 11942 4936
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 9968 3194 9996 3538
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 11164 3058 11192 3538
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11164 2922 11192 2994
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 11532 2582 11560 3606
rect 12268 3505 12296 8842
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12360 6458 12388 6938
rect 12544 6730 12572 8230
rect 12636 7857 12664 8230
rect 12622 7848 12678 7857
rect 12622 7783 12624 7792
rect 12676 7783 12678 7792
rect 12624 7754 12676 7760
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12820 7041 12848 7346
rect 13464 7342 13492 7686
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13556 7274 13584 9007
rect 13648 8514 13676 12974
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13740 11558 13768 12378
rect 13820 12232 13872 12238
rect 13924 12220 13952 13806
rect 13872 12192 13952 12220
rect 13820 12174 13872 12180
rect 13832 11694 13860 12174
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 14016 11354 14044 14311
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14016 9586 14044 10202
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14016 9178 14044 9522
rect 14004 9172 14056 9178
rect 14056 9132 14136 9160
rect 14004 9114 14056 9120
rect 13648 8486 13768 8514
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 12806 7032 12862 7041
rect 12806 6967 12862 6976
rect 13004 6866 13032 7142
rect 13648 7002 13676 7686
rect 13740 7410 13768 8486
rect 14108 8430 14136 9132
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14200 8090 14228 21014
rect 14292 19310 14320 21270
rect 15764 19378 15792 23520
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 16486 20360 16542 20369
rect 16486 20295 16542 20304
rect 16500 20262 16528 20295
rect 16488 20256 16540 20262
rect 17236 20244 17264 23520
rect 18234 20360 18290 20369
rect 18234 20295 18290 20304
rect 18248 20262 18276 20295
rect 18236 20256 18288 20262
rect 17236 20216 17448 20244
rect 16488 20198 16540 20204
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 17328 19514 17356 19858
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17420 19446 17448 20216
rect 18236 20198 18288 20204
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18616 19961 18644 19994
rect 18602 19952 18658 19961
rect 18602 19887 18658 19896
rect 17498 19816 17554 19825
rect 17498 19751 17500 19760
rect 17552 19751 17554 19760
rect 17500 19722 17552 19728
rect 17408 19440 17460 19446
rect 17408 19382 17460 19388
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14384 8566 14412 8774
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 14016 7274 14044 7890
rect 14200 7721 14228 8026
rect 14186 7712 14242 7721
rect 14186 7647 14242 7656
rect 14200 7546 14228 7647
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12912 4826 12940 6598
rect 13004 5914 13032 6802
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13464 6202 13492 6734
rect 13740 6254 13768 7142
rect 14016 7002 14044 7210
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 13372 6174 13492 6202
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13544 6180 13596 6186
rect 13372 6118 13400 6174
rect 13544 6122 13596 6128
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13372 5370 13400 6054
rect 13556 5914 13584 6122
rect 14278 5944 14334 5953
rect 13544 5908 13596 5914
rect 14278 5879 14280 5888
rect 13544 5850 13596 5856
rect 14332 5879 14334 5888
rect 14280 5850 14332 5856
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13556 5250 13584 5850
rect 14384 5778 14412 8502
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 13372 5222 13584 5250
rect 13372 5166 13400 5222
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13372 4826 13400 5102
rect 14384 4826 14412 5714
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12360 4049 12388 4422
rect 12346 4040 12402 4049
rect 12346 3975 12402 3984
rect 12728 3942 12756 4558
rect 12912 4282 12940 4762
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13096 4321 13124 4626
rect 13082 4312 13138 4321
rect 12900 4276 12952 4282
rect 13082 4247 13084 4256
rect 12900 4218 12952 4224
rect 13136 4247 13138 4256
rect 13084 4218 13136 4224
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12254 3496 12310 3505
rect 12254 3431 12310 3440
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 11610 2816 11666 2825
rect 11610 2751 11666 2760
rect 11624 2650 11652 2751
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10796 480 10824 2246
rect 11808 480 11836 3334
rect 12452 3194 12480 3334
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12728 3074 12756 3878
rect 13372 3738 13400 4762
rect 14370 4584 14426 4593
rect 14370 4519 14426 4528
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 12360 3058 12756 3074
rect 12348 3052 12756 3058
rect 12400 3046 12756 3052
rect 12348 2994 12400 3000
rect 12728 2990 12756 3046
rect 12716 2984 12768 2990
rect 12070 2952 12126 2961
rect 12070 2887 12126 2896
rect 12452 2922 12664 2938
rect 12716 2926 12768 2932
rect 13818 2952 13874 2961
rect 12452 2916 12676 2922
rect 12452 2910 12624 2916
rect 12084 2650 12112 2887
rect 12452 2650 12480 2910
rect 13818 2887 13874 2896
rect 12624 2858 12676 2864
rect 13832 2854 13860 2887
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13910 2816 13966 2825
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12820 480 12848 2790
rect 13910 2751 13966 2760
rect 13924 480 13952 2751
rect 14108 2650 14136 3674
rect 14278 3088 14334 3097
rect 14278 3023 14334 3032
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14292 2514 14320 3023
rect 14384 2961 14412 4519
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14476 3194 14504 3538
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14370 2952 14426 2961
rect 14370 2887 14426 2896
rect 14462 2816 14518 2825
rect 14462 2751 14518 2760
rect 14476 2650 14504 2751
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14568 2553 14596 19246
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 15750 17096 15806 17105
rect 15750 17031 15806 17040
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14936 12782 14964 13126
rect 15028 12782 15056 13670
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14936 12306 14964 12718
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14936 10266 14964 12242
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14936 8838 14964 10066
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 15396 8430 15424 9318
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 14844 8090 14872 8366
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14844 7886 14872 8026
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 6882 15148 7142
rect 15120 6854 15240 6882
rect 15212 6662 15240 6854
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15120 5930 15148 6054
rect 15120 5902 15424 5930
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5545 15332 5578
rect 15290 5536 15346 5545
rect 15290 5471 15346 5480
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14752 2990 14780 4966
rect 15396 4622 15424 5902
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 4321 15332 4422
rect 15290 4312 15346 4321
rect 15396 4282 15424 4558
rect 15290 4247 15346 4256
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14936 2990 14964 3674
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14554 2544 14610 2553
rect 14280 2508 14332 2514
rect 14936 2514 14964 2926
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 15212 2650 15240 2858
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15304 2530 15332 2790
rect 15488 2689 15516 12038
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15672 9897 15700 10066
rect 15658 9888 15714 9897
rect 15658 9823 15714 9832
rect 15764 6769 15792 17031
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 16408 11880 16436 12582
rect 16500 12102 16528 19314
rect 17682 13152 17738 13161
rect 17682 13087 17738 13096
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16592 11898 16620 12242
rect 16580 11892 16632 11898
rect 16408 11852 16580 11880
rect 16408 11801 16436 11852
rect 16580 11834 16632 11840
rect 16394 11792 16450 11801
rect 16394 11727 16450 11736
rect 16960 11694 16988 12310
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 17696 11218 17724 13087
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 16500 10690 16528 11018
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16500 10674 16620 10690
rect 16500 10668 16632 10674
rect 16500 10662 16580 10668
rect 16580 10610 16632 10616
rect 16776 10606 16804 10950
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 17052 10538 17080 10610
rect 17040 10532 17092 10538
rect 17040 10474 17092 10480
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15856 9382 15884 10066
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 16408 9625 16436 10406
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9761 16528 9862
rect 16486 9752 16542 9761
rect 16486 9687 16542 9696
rect 16394 9616 16450 9625
rect 16394 9551 16450 9560
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16210 9208 16266 9217
rect 16210 9143 16266 9152
rect 16224 9110 16252 9143
rect 16212 9104 16264 9110
rect 16264 9052 16436 9058
rect 16212 9046 16436 9052
rect 16224 9030 16436 9046
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 16316 8294 16344 8910
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16408 8090 16436 9030
rect 16500 8634 16528 9318
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16592 7954 16620 8230
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 16500 7478 16528 7822
rect 16592 7546 16620 7890
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 15750 6760 15806 6769
rect 15750 6695 15806 6704
rect 15764 6458 15792 6695
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15764 6254 15792 6394
rect 16500 6361 16528 6598
rect 16486 6352 16542 6361
rect 16212 6316 16264 6322
rect 16486 6287 16488 6296
rect 16212 6258 16264 6264
rect 16540 6287 16542 6296
rect 16488 6258 16540 6264
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15580 5370 15608 5646
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15764 4826 15792 5510
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15764 4282 15792 4762
rect 15856 4758 15884 6054
rect 16224 5710 16252 6258
rect 16396 6180 16448 6186
rect 16396 6122 16448 6128
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16302 5672 16358 5681
rect 16302 5607 16358 5616
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 16316 5030 16344 5607
rect 16408 5370 16436 6122
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16500 5545 16528 5714
rect 16684 5642 16712 9318
rect 16868 9110 16896 10202
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16486 5536 16542 5545
rect 16486 5471 16542 5480
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 15844 4752 15896 4758
rect 15844 4694 15896 4700
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15856 4214 15884 4694
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 16500 4078 16528 5471
rect 16762 5264 16818 5273
rect 16762 5199 16818 5208
rect 16776 5166 16804 5199
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16776 4826 16804 5102
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16868 4593 16896 4966
rect 16854 4584 16910 4593
rect 16854 4519 16910 4528
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16960 3641 16988 10406
rect 17052 10062 17080 10474
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17052 9518 17080 9998
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17052 9110 17080 9454
rect 17236 9382 17264 10134
rect 17328 10062 17356 11154
rect 17408 11144 17460 11150
rect 17788 11098 17816 19382
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17408 11086 17460 11092
rect 17420 10470 17448 11086
rect 17696 11070 17816 11098
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 10056 17368 10062
rect 17314 10024 17316 10033
rect 17408 10056 17460 10062
rect 17368 10024 17370 10033
rect 17408 9998 17460 10004
rect 17314 9959 17370 9968
rect 17420 9908 17448 9998
rect 17328 9880 17448 9908
rect 17328 9518 17356 9880
rect 17696 9636 17724 11070
rect 17972 10713 18000 12922
rect 18708 12481 18736 23520
rect 20180 21162 20208 23520
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 20088 21134 20208 21162
rect 19430 20632 19486 20641
rect 19430 20567 19432 20576
rect 19484 20567 19486 20576
rect 19432 20538 19484 20544
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18786 19408 18842 19417
rect 18786 19343 18842 19352
rect 18694 12472 18750 12481
rect 18694 12407 18750 12416
rect 18418 12336 18474 12345
rect 18418 12271 18474 12280
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18248 11898 18276 12038
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18248 11150 18276 11834
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 17774 10704 17830 10713
rect 17774 10639 17776 10648
rect 17828 10639 17830 10648
rect 17958 10704 18014 10713
rect 18248 10674 18276 11086
rect 18432 11014 18460 12271
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11694 18552 12038
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18708 11694 18736 11834
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 17958 10639 18014 10648
rect 18236 10668 18288 10674
rect 17776 10610 17828 10616
rect 18236 10610 18288 10616
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18144 10260 18196 10266
rect 18064 10220 18144 10248
rect 18064 10130 18092 10220
rect 18144 10202 18196 10208
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17960 9648 18012 9654
rect 17696 9608 17960 9636
rect 17960 9590 18012 9596
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17144 4729 17172 8570
rect 17328 5409 17356 9454
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17420 8974 17448 9386
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18064 9217 18092 9318
rect 18050 9208 18106 9217
rect 17776 9172 17828 9178
rect 18050 9143 18106 9152
rect 17776 9114 17828 9120
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17420 8634 17448 8910
rect 17788 8634 17816 9114
rect 18340 8838 18368 10542
rect 18432 10470 18460 10950
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18420 10464 18472 10470
rect 18418 10432 18420 10441
rect 18472 10432 18474 10441
rect 18418 10367 18474 10376
rect 18708 10266 18736 10610
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18708 10062 18736 10202
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18418 9752 18474 9761
rect 18708 9722 18736 9998
rect 18418 9687 18474 9696
rect 18696 9716 18748 9722
rect 18432 9518 18460 9687
rect 18696 9658 18748 9664
rect 18510 9616 18566 9625
rect 18510 9551 18512 9560
rect 18564 9551 18566 9560
rect 18696 9580 18748 9586
rect 18512 9522 18564 9528
rect 18696 9522 18748 9528
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17314 5400 17370 5409
rect 17314 5335 17370 5344
rect 17328 4865 17356 5335
rect 17420 5137 17448 8298
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17880 6934 17908 7686
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17682 6488 17738 6497
rect 17880 6458 17908 6734
rect 17682 6423 17738 6432
rect 17868 6452 17920 6458
rect 17498 6080 17554 6089
rect 17498 6015 17554 6024
rect 17512 5710 17540 6015
rect 17696 5914 17724 6423
rect 17868 6394 17920 6400
rect 17880 5953 17908 6394
rect 17866 5944 17922 5953
rect 17684 5908 17736 5914
rect 17604 5868 17684 5896
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17406 5128 17462 5137
rect 17406 5063 17462 5072
rect 17512 5030 17540 5646
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17314 4856 17370 4865
rect 17314 4791 17370 4800
rect 17130 4720 17186 4729
rect 17130 4655 17186 4664
rect 16946 3632 17002 3641
rect 16488 3596 16540 3602
rect 16540 3556 16620 3584
rect 16946 3567 17002 3576
rect 16488 3538 16540 3544
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15474 2680 15530 2689
rect 15474 2615 15530 2624
rect 14554 2479 14610 2488
rect 14924 2508 14976 2514
rect 14280 2450 14332 2456
rect 14924 2450 14976 2456
rect 15120 2502 15332 2530
rect 15120 2446 15148 2502
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 14924 2372 14976 2378
rect 14924 2314 14976 2320
rect 14936 480 14964 2314
rect 15856 1442 15884 3334
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 16592 2650 16620 3556
rect 17512 3097 17540 4966
rect 17604 4758 17632 5868
rect 17866 5879 17922 5888
rect 17684 5850 17736 5856
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17696 5234 17724 5578
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17696 4826 17724 5170
rect 17776 5024 17828 5030
rect 17774 4992 17776 5001
rect 17828 4992 17830 5001
rect 17774 4927 17830 4936
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17592 4752 17644 4758
rect 17592 4694 17644 4700
rect 17498 3088 17554 3097
rect 17498 3023 17554 3032
rect 17972 2990 18000 8774
rect 18524 8634 18552 8978
rect 18708 8974 18736 9522
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18326 8528 18382 8537
rect 18326 8463 18328 8472
rect 18380 8463 18382 8472
rect 18328 8434 18380 8440
rect 18418 7984 18474 7993
rect 18418 7919 18474 7928
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18156 6746 18184 6802
rect 18156 6718 18276 6746
rect 18248 6118 18276 6718
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 5710 18276 6054
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18050 5536 18106 5545
rect 18050 5471 18106 5480
rect 18064 5370 18092 5471
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 18432 5166 18460 7919
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18432 4826 18460 5102
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18524 4457 18552 5034
rect 18510 4448 18566 4457
rect 18510 4383 18566 4392
rect 18800 4185 18828 19343
rect 18892 8378 18920 20198
rect 18984 19360 19012 20334
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19064 19372 19116 19378
rect 18984 19332 19064 19360
rect 19116 19332 19196 19360
rect 19064 19314 19116 19320
rect 18970 15056 19026 15065
rect 18970 14991 19026 15000
rect 18984 9178 19012 14991
rect 19062 12472 19118 12481
rect 19062 12407 19118 12416
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18984 8634 19012 9114
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18892 8350 19012 8378
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18892 8090 18920 8230
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18878 7440 18934 7449
rect 18878 7375 18934 7384
rect 18892 7342 18920 7375
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18786 4176 18842 4185
rect 18786 4111 18842 4120
rect 18984 4026 19012 8350
rect 18064 3998 19012 4026
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 16946 2816 17002 2825
rect 16946 2751 17002 2760
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 15856 1414 15976 1442
rect 15948 480 15976 1414
rect 16960 480 16988 2751
rect 18064 480 18092 3998
rect 19076 3641 19104 12407
rect 19168 9625 19196 19332
rect 19444 19242 19472 19858
rect 19706 19816 19762 19825
rect 19706 19751 19708 19760
rect 19760 19751 19762 19760
rect 19708 19722 19760 19728
rect 19432 19236 19484 19242
rect 19432 19178 19484 19184
rect 19800 19168 19852 19174
rect 19800 19110 19852 19116
rect 19340 16040 19392 16046
rect 19338 16008 19340 16017
rect 19392 16008 19394 16017
rect 19338 15943 19394 15952
rect 19338 12472 19394 12481
rect 19338 12407 19394 12416
rect 19246 9752 19302 9761
rect 19246 9687 19302 9696
rect 19154 9616 19210 9625
rect 19154 9551 19210 9560
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 19168 4049 19196 9386
rect 19260 8566 19288 9687
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19352 7546 19380 12407
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 8974 19472 11494
rect 19812 9722 19840 19110
rect 20088 12481 20116 21134
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 20180 20330 20208 20946
rect 21560 20602 21588 20946
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 20628 20528 20680 20534
rect 20626 20496 20628 20505
rect 20680 20496 20682 20505
rect 20626 20431 20682 20440
rect 21744 20369 21772 23520
rect 23216 20641 23244 23520
rect 23202 20632 23258 20641
rect 22008 20596 22060 20602
rect 23202 20567 23258 20576
rect 22008 20538 22060 20544
rect 22020 20369 22048 20538
rect 23848 20528 23900 20534
rect 23846 20496 23848 20505
rect 23900 20496 23902 20505
rect 23846 20431 23902 20440
rect 22284 20392 22336 20398
rect 21730 20360 21786 20369
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 20720 20324 20772 20330
rect 21730 20295 21786 20304
rect 22006 20360 22062 20369
rect 23664 20392 23716 20398
rect 22284 20334 22336 20340
rect 23662 20360 23664 20369
rect 23716 20360 23718 20369
rect 22006 20295 22062 20304
rect 20720 20266 20772 20272
rect 20732 19922 20760 20266
rect 21916 20256 21968 20262
rect 21914 20224 21916 20233
rect 21968 20224 21970 20233
rect 20956 20156 21252 20176
rect 22020 20210 22048 20295
rect 22020 20182 22140 20210
rect 21914 20159 21970 20168
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21560 19961 21588 19994
rect 21546 19952 21602 19961
rect 20720 19916 20772 19922
rect 21546 19887 21602 19896
rect 20720 19858 20772 19864
rect 20732 19174 20760 19858
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20074 12472 20130 12481
rect 20074 12407 20130 12416
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19444 8498 19472 8910
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19444 8090 19472 8434
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 6361 19288 6598
rect 19246 6352 19302 6361
rect 19246 6287 19302 6296
rect 19154 4040 19210 4049
rect 19154 3975 19210 3984
rect 18418 3632 18474 3641
rect 18418 3567 18474 3576
rect 19062 3632 19118 3641
rect 19062 3567 19118 3576
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 1674 368 1730 377
rect 1674 303 1730 312
rect 2502 0 2558 480
rect 3514 0 3570 480
rect 4526 0 4582 480
rect 5630 0 5686 480
rect 6642 0 6698 480
rect 7654 0 7710 480
rect 8666 0 8722 480
rect 9770 0 9826 480
rect 10782 0 10838 480
rect 11794 0 11850 480
rect 12806 0 12862 480
rect 13910 0 13966 480
rect 14922 0 14978 480
rect 15934 0 15990 480
rect 16946 0 17002 480
rect 18050 0 18106 480
rect 18340 377 18368 2790
rect 18432 2514 18460 3567
rect 19430 2680 19486 2689
rect 19430 2615 19486 2624
rect 19444 2514 19472 2615
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19154 2408 19210 2417
rect 19154 2343 19210 2352
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18524 1465 18552 2246
rect 18510 1456 18566 1465
rect 18510 1391 18566 1400
rect 19168 610 19196 2343
rect 19536 1442 19564 9658
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19628 8673 19656 9046
rect 19614 8664 19670 8673
rect 19614 8599 19670 8608
rect 19892 8628 19944 8634
rect 19628 8362 19656 8599
rect 19892 8570 19944 8576
rect 19904 8401 19932 8570
rect 19890 8392 19946 8401
rect 19616 8356 19668 8362
rect 19890 8327 19946 8336
rect 19616 8298 19668 8304
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 19614 3496 19670 3505
rect 19614 3431 19670 3440
rect 19628 2650 19656 3431
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 20180 2417 20208 7482
rect 20166 2408 20222 2417
rect 20166 2343 20222 2352
rect 19536 1414 20116 1442
rect 19064 604 19116 610
rect 19064 546 19116 552
rect 19156 604 19208 610
rect 19156 546 19208 552
rect 19076 480 19104 546
rect 20088 480 20116 1414
rect 20732 1306 20760 19110
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21376 15881 21404 15982
rect 21362 15872 21418 15881
rect 20956 15804 21252 15824
rect 21362 15807 21418 15816
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 21362 14648 21418 14657
rect 21362 14583 21418 14592
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 21376 10198 21404 14583
rect 21364 10192 21416 10198
rect 21364 10134 21416 10140
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 22112 7546 22140 20182
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 20732 1278 21128 1306
rect 21100 480 21128 1278
rect 22296 626 22324 20334
rect 23662 20295 23718 20304
rect 24688 19825 24716 23520
rect 24858 22400 24914 22409
rect 24858 22335 24914 22344
rect 24872 22166 24900 22335
rect 24860 22160 24912 22166
rect 24860 22102 24912 22108
rect 25320 21684 25372 21690
rect 25320 21626 25372 21632
rect 24674 19816 24730 19825
rect 24674 19751 24730 19760
rect 25042 19408 25098 19417
rect 25042 19343 25098 19352
rect 25056 14929 25084 19343
rect 25042 14920 25098 14929
rect 25042 14855 25098 14864
rect 25042 13968 25098 13977
rect 25042 13903 25098 13912
rect 25056 7993 25084 13903
rect 25332 13025 25360 21626
rect 25410 20088 25466 20097
rect 25410 20023 25466 20032
rect 25424 14385 25452 20023
rect 25410 14376 25466 14385
rect 25410 14311 25466 14320
rect 25318 13016 25374 13025
rect 25318 12951 25374 12960
rect 25318 12880 25374 12889
rect 25318 12815 25374 12824
rect 25042 7984 25098 7993
rect 25042 7919 25098 7928
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23018 2816 23074 2825
rect 23018 2751 23074 2760
rect 23032 2650 23060 2751
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 22834 2544 22890 2553
rect 22834 2479 22836 2488
rect 22888 2479 22890 2488
rect 22836 2450 22888 2456
rect 22204 598 22324 626
rect 22204 480 22232 598
rect 23216 480 23244 7482
rect 25332 6497 25360 12815
rect 25516 11665 25544 23559
rect 26238 23520 26294 24000
rect 27710 23520 27766 24000
rect 29182 23520 29238 24000
rect 25686 23080 25742 23089
rect 25686 23015 25742 23024
rect 25700 21690 25728 23015
rect 26252 21978 26280 23520
rect 26252 21950 26372 21978
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25686 21584 25742 21593
rect 25686 21519 25742 21528
rect 25700 20942 25728 21519
rect 25778 21312 25834 21321
rect 25778 21247 25834 21256
rect 25792 21078 25820 21247
rect 25780 21072 25832 21078
rect 25780 21014 25832 21020
rect 25688 20936 25740 20942
rect 25688 20878 25740 20884
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 25594 20360 25650 20369
rect 25594 20295 25650 20304
rect 25502 11656 25558 11665
rect 25502 11591 25558 11600
rect 25608 9761 25636 20295
rect 26344 19961 26372 21950
rect 27724 20233 27752 23520
rect 29196 20505 29224 23520
rect 29182 20496 29238 20505
rect 29182 20431 29238 20440
rect 27710 20224 27766 20233
rect 27710 20159 27766 20168
rect 26330 19952 26386 19961
rect 26330 19887 26386 19896
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 25778 17096 25834 17105
rect 25778 17031 25834 17040
rect 25686 16144 25742 16153
rect 25686 16079 25742 16088
rect 25700 13433 25728 16079
rect 25686 13424 25742 13433
rect 25686 13359 25742 13368
rect 25594 9752 25650 9761
rect 25594 9687 25650 9696
rect 25792 8673 25820 17031
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 25870 15464 25926 15473
rect 25870 15399 25926 15408
rect 25778 8664 25834 8673
rect 25778 8599 25834 8608
rect 25884 6882 25912 15399
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 27526 14512 27582 14521
rect 27526 14447 27582 14456
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 26146 12744 26202 12753
rect 26146 12679 26202 12688
rect 26160 12186 26188 12679
rect 26160 12170 26280 12186
rect 26160 12164 26292 12170
rect 26160 12158 26240 12164
rect 26240 12106 26292 12112
rect 26516 12164 26568 12170
rect 26516 12106 26568 12112
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26436 11121 26464 11630
rect 26528 11218 26556 12106
rect 26606 11656 26662 11665
rect 26606 11591 26662 11600
rect 26620 11558 26648 11591
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26516 11212 26568 11218
rect 26516 11154 26568 11160
rect 26422 11112 26478 11121
rect 26422 11047 26478 11056
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 26528 10810 26556 11154
rect 26698 11112 26754 11121
rect 26698 11047 26700 11056
rect 26752 11047 26754 11056
rect 26700 11018 26752 11024
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26330 10704 26386 10713
rect 26330 10639 26386 10648
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 25792 6854 25912 6882
rect 25318 6488 25374 6497
rect 25318 6423 25374 6432
rect 24398 5400 24454 5409
rect 24398 5335 24454 5344
rect 24412 5001 24440 5335
rect 25792 5273 25820 6854
rect 25870 6760 25926 6769
rect 25870 6695 25926 6704
rect 25884 5370 25912 6695
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 25872 5364 25924 5370
rect 25872 5306 25924 5312
rect 25778 5264 25834 5273
rect 25778 5199 25834 5208
rect 24398 4992 24454 5001
rect 24398 4927 24454 4936
rect 25686 4448 25742 4457
rect 25686 4383 25742 4392
rect 24214 4176 24270 4185
rect 24214 4111 24270 4120
rect 24228 480 24256 4111
rect 25318 4040 25374 4049
rect 25318 3975 25374 3984
rect 25134 3632 25190 3641
rect 25332 3602 25360 3975
rect 25134 3567 25190 3576
rect 25320 3596 25372 3602
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 25056 2961 25084 3470
rect 25148 3194 25176 3567
rect 25320 3538 25372 3544
rect 25332 3194 25360 3538
rect 25504 3392 25556 3398
rect 25504 3334 25556 3340
rect 25136 3188 25188 3194
rect 25136 3130 25188 3136
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 25148 2990 25176 3130
rect 25516 3097 25544 3334
rect 25502 3088 25558 3097
rect 25502 3023 25558 3032
rect 25136 2984 25188 2990
rect 25042 2952 25098 2961
rect 25136 2926 25188 2932
rect 25042 2887 25098 2896
rect 25504 2848 25556 2854
rect 25226 2816 25282 2825
rect 25226 2751 25282 2760
rect 25502 2816 25504 2825
rect 25556 2816 25558 2825
rect 25502 2751 25558 2760
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24596 2417 24624 2450
rect 24582 2408 24638 2417
rect 24582 2343 24638 2352
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24780 1737 24808 2246
rect 24766 1728 24822 1737
rect 24766 1663 24822 1672
rect 25240 480 25268 2751
rect 25700 2514 25728 4383
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 26344 4078 26372 10639
rect 26698 10432 26754 10441
rect 26698 10367 26754 10376
rect 26712 10266 26740 10367
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26528 9518 26556 10066
rect 26698 9888 26754 9897
rect 26698 9823 26754 9832
rect 26516 9512 26568 9518
rect 26514 9480 26516 9489
rect 26568 9480 26570 9489
rect 26514 9415 26570 9424
rect 26606 9344 26662 9353
rect 26606 9279 26662 9288
rect 26422 9072 26478 9081
rect 26422 9007 26478 9016
rect 26516 9036 26568 9042
rect 26436 8430 26464 9007
rect 26516 8978 26568 8984
rect 26528 8945 26556 8978
rect 26514 8936 26570 8945
rect 26514 8871 26570 8880
rect 26528 8566 26556 8871
rect 26620 8634 26648 9279
rect 26712 9178 26740 9823
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26698 8664 26754 8673
rect 26608 8628 26660 8634
rect 26698 8599 26754 8608
rect 26608 8570 26660 8576
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26514 8392 26570 8401
rect 26514 8327 26570 8336
rect 26528 7954 26556 8327
rect 26712 8090 26740 8599
rect 27540 8430 27568 14447
rect 27712 8560 27764 8566
rect 27712 8502 27764 8508
rect 27528 8424 27580 8430
rect 27724 8401 27752 8502
rect 27528 8366 27580 8372
rect 27710 8392 27766 8401
rect 27710 8327 27766 8336
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 26528 7546 26556 7890
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 26698 7440 26754 7449
rect 26698 7375 26754 7384
rect 26608 7200 26660 7206
rect 26608 7142 26660 7148
rect 26620 7041 26648 7142
rect 26606 7032 26662 7041
rect 26606 6967 26662 6976
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26528 6254 26556 6802
rect 26712 6730 26740 7375
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26698 6352 26754 6361
rect 26698 6287 26754 6296
rect 26516 6248 26568 6254
rect 26514 6216 26516 6225
rect 26568 6216 26570 6225
rect 26514 6151 26570 6160
rect 26712 5914 26740 6287
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 26514 5808 26570 5817
rect 26514 5743 26516 5752
rect 26568 5743 26570 5752
rect 26516 5714 26568 5720
rect 26528 5302 26556 5714
rect 26606 5672 26662 5681
rect 26606 5607 26662 5616
rect 26620 5370 26648 5607
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26516 5296 26568 5302
rect 26516 5238 26568 5244
rect 26698 5128 26754 5137
rect 26698 5063 26754 5072
rect 26712 4826 26740 5063
rect 26790 4992 26846 5001
rect 26790 4927 26846 4936
rect 26700 4820 26752 4826
rect 26700 4762 26752 4768
rect 26514 4720 26570 4729
rect 26514 4655 26516 4664
rect 26568 4655 26570 4664
rect 26516 4626 26568 4632
rect 26422 4584 26478 4593
rect 26422 4519 26478 4528
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26330 3496 26386 3505
rect 26330 3431 26386 3440
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 25688 2508 25740 2514
rect 25688 2450 25740 2456
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25884 2009 25912 2246
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 25870 2000 25926 2009
rect 25870 1935 25926 1944
rect 26344 480 26372 3431
rect 26436 2990 26464 4519
rect 26528 4282 26556 4626
rect 26606 4448 26662 4457
rect 26606 4383 26662 4392
rect 26516 4276 26568 4282
rect 26516 4218 26568 4224
rect 26620 3942 26648 4383
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26698 3904 26754 3913
rect 26698 3839 26754 3848
rect 26712 3738 26740 3839
rect 26700 3732 26752 3738
rect 26700 3674 26752 3680
rect 26606 3360 26662 3369
rect 26606 3295 26662 3304
rect 26620 3194 26648 3295
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26804 2514 26832 4927
rect 27344 3528 27396 3534
rect 27344 3470 27396 3476
rect 27356 3194 27384 3470
rect 27344 3188 27396 3194
rect 27344 3130 27396 3136
rect 27342 3088 27398 3097
rect 27342 3023 27398 3032
rect 27066 2680 27122 2689
rect 27066 2615 27068 2624
rect 27120 2615 27122 2624
rect 27068 2586 27120 2592
rect 26792 2508 26844 2514
rect 26792 2450 26844 2456
rect 27356 480 27384 3023
rect 27528 2984 27580 2990
rect 27526 2952 27528 2961
rect 27580 2952 27582 2961
rect 27526 2887 27582 2896
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 28354 2816 28410 2825
rect 27724 921 27752 2790
rect 28354 2751 28410 2760
rect 27710 912 27766 921
rect 27710 847 27766 856
rect 28368 480 28396 2751
rect 29366 1728 29422 1737
rect 29366 1663 29422 1672
rect 29380 480 29408 1663
rect 18326 368 18382 377
rect 18326 303 18382 312
rect 19062 0 19118 480
rect 20074 0 20130 480
rect 21086 0 21142 480
rect 22190 0 22246 480
rect 23202 0 23258 480
rect 24214 0 24270 480
rect 25226 0 25282 480
rect 26330 0 26386 480
rect 27342 0 27398 480
rect 28354 0 28410 480
rect 29366 0 29422 480
<< via2 >>
rect 2962 23568 3018 23624
rect 754 20304 810 20360
rect 2778 23024 2834 23080
rect 2226 19760 2282 19816
rect 25502 23568 25558 23624
rect 2778 19352 2834 19408
rect 2318 14592 2374 14648
rect 1490 13232 1546 13288
rect 2042 12316 2044 12336
rect 2044 12316 2096 12336
rect 2096 12316 2098 12336
rect 2042 12280 2098 12316
rect 1582 11600 1638 11656
rect 1582 11056 1638 11112
rect 2042 10804 2098 10840
rect 2042 10784 2044 10804
rect 2044 10784 2096 10804
rect 2096 10784 2098 10804
rect 1582 10376 1638 10432
rect 2962 15272 3018 15328
rect 2502 10512 2558 10568
rect 1582 9832 1638 9888
rect 1582 9288 1638 9344
rect 1582 8628 1638 8664
rect 1582 8608 1584 8628
rect 1584 8608 1636 8628
rect 1636 8608 1638 8628
rect 2042 8492 2098 8528
rect 2042 8472 2044 8492
rect 2044 8472 2096 8492
rect 2096 8472 2098 8492
rect 1950 8200 2006 8256
rect 1674 6568 1730 6624
rect 1582 5616 1638 5672
rect 1582 4428 1584 4448
rect 1584 4428 1636 4448
rect 1636 4428 1638 4448
rect 1582 4392 1638 4428
rect 1582 3884 1584 3904
rect 1584 3884 1636 3904
rect 1636 3884 1638 3904
rect 1582 3848 1638 3884
rect 1582 3340 1584 3360
rect 1584 3340 1636 3360
rect 1636 3340 1638 3360
rect 1582 3304 1638 3340
rect 1490 2760 1546 2816
rect 1398 856 1454 912
rect 2686 11756 2742 11792
rect 2686 11736 2688 11756
rect 2688 11736 2740 11756
rect 2740 11736 2742 11756
rect 3054 12008 3110 12064
rect 3054 10648 3110 10704
rect 2686 8064 2742 8120
rect 2686 7828 2688 7848
rect 2688 7828 2740 7848
rect 2740 7828 2742 7848
rect 2686 7792 2742 7828
rect 2134 6160 2190 6216
rect 2594 7384 2650 7440
rect 2042 5888 2098 5944
rect 2226 4936 2282 4992
rect 2502 5208 2558 5264
rect 2686 5072 2742 5128
rect 4066 22364 4122 22400
rect 4066 22344 4068 22364
rect 4068 22344 4120 22364
rect 4120 22344 4122 22364
rect 3974 21800 4030 21856
rect 3882 21256 3938 21312
rect 3882 20576 3938 20632
rect 3698 19896 3754 19952
rect 3422 18264 3478 18320
rect 3698 18264 3754 18320
rect 3238 14048 3294 14104
rect 3330 12724 3332 12744
rect 3332 12724 3384 12744
rect 3384 12724 3386 12744
rect 3330 12688 3386 12724
rect 3330 12416 3386 12472
rect 3238 11600 3294 11656
rect 3514 14864 3570 14920
rect 3882 15000 3938 15056
rect 3698 13368 3754 13424
rect 3514 12824 3570 12880
rect 3514 12144 3570 12200
rect 3238 11056 3294 11112
rect 3146 6024 3202 6080
rect 2686 2624 2742 2680
rect 3422 10260 3478 10296
rect 3422 10240 3424 10260
rect 3424 10240 3476 10260
rect 3476 10240 3478 10260
rect 3330 8064 3386 8120
rect 3330 6976 3386 7032
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 6734 20440 6790 20496
rect 4066 20032 4122 20088
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 7838 16904 7894 16960
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 4618 15952 4674 16008
rect 4342 15816 4398 15872
rect 4066 14456 4122 14512
rect 3790 12552 3846 12608
rect 3974 12552 4030 12608
rect 3790 12416 3846 12472
rect 3882 8880 3938 8936
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5078 12824 5134 12880
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 6734 12008 6790 12064
rect 7194 12280 7250 12336
rect 7654 12008 7710 12064
rect 4434 10784 4490 10840
rect 4802 10648 4858 10704
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 4250 10104 4306 10160
rect 4066 8880 4122 8936
rect 4250 6840 4306 6896
rect 3790 6332 3792 6352
rect 3792 6332 3844 6352
rect 3844 6332 3846 6352
rect 3790 6296 3846 6332
rect 4250 5480 4306 5536
rect 4342 4664 4398 4720
rect 4526 10376 4582 10432
rect 4434 4528 4490 4584
rect 7562 10784 7618 10840
rect 7562 10512 7618 10568
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 4618 8200 4674 8256
rect 4618 6332 4620 6352
rect 4620 6332 4672 6352
rect 4672 6332 4674 6352
rect 4618 6296 4674 6332
rect 4434 3576 4490 3632
rect 2962 2080 3018 2136
rect 2778 1400 2834 1456
rect 7838 9832 7894 9888
rect 7470 9696 7526 9752
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 4986 5772 5042 5808
rect 4986 5752 4988 5772
rect 4988 5752 5040 5772
rect 5040 5752 5042 5772
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 5262 3440 5318 3496
rect 5538 2760 5594 2816
rect 4618 1536 4674 1592
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 7930 8628 7986 8664
rect 7930 8608 7932 8628
rect 7932 8608 7984 8628
rect 7984 8608 7986 8628
rect 7194 6196 7196 6216
rect 7196 6196 7248 6216
rect 7248 6196 7250 6216
rect 7194 6160 7250 6196
rect 8482 4020 8484 4040
rect 8484 4020 8536 4040
rect 8536 4020 8538 4040
rect 8482 3984 8538 4020
rect 9218 18808 9274 18864
rect 9034 11620 9090 11656
rect 9034 11600 9036 11620
rect 9036 11600 9088 11620
rect 9088 11600 9090 11620
rect 9494 16496 9550 16552
rect 9402 12144 9458 12200
rect 9034 7792 9090 7848
rect 9218 7384 9274 7440
rect 8666 7248 8722 7304
rect 8574 3848 8630 3904
rect 8574 3032 8630 3088
rect 6274 2896 6330 2952
rect 8482 2896 8538 2952
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 6642 1536 6698 1592
rect 10046 9696 10102 9752
rect 9954 8608 10010 8664
rect 9770 8064 9826 8120
rect 9770 6160 9826 6216
rect 9310 6060 9312 6080
rect 9312 6060 9364 6080
rect 9364 6060 9366 6080
rect 9310 6024 9366 6060
rect 10138 5888 10194 5944
rect 9310 5616 9366 5672
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 12070 18808 12126 18864
rect 11978 17992 12034 18048
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 11794 14492 11796 14512
rect 11796 14492 11848 14512
rect 11848 14492 11850 14512
rect 11794 14456 11850 14492
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 11794 13232 11850 13288
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 11702 11056 11758 11112
rect 11978 10920 12034 10976
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 11150 9460 11152 9480
rect 11152 9460 11204 9480
rect 11204 9460 11206 9480
rect 11150 9424 11206 9460
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 10782 7928 10838 7984
rect 10690 6976 10746 7032
rect 12714 19352 12770 19408
rect 12530 18128 12586 18184
rect 12898 13388 12954 13424
rect 12898 13368 12900 13388
rect 12900 13368 12952 13388
rect 12952 13368 12954 13388
rect 12346 11772 12348 11792
rect 12348 11772 12400 11792
rect 12400 11772 12402 11792
rect 12346 11736 12402 11772
rect 13450 17720 13506 17776
rect 14002 14320 14058 14376
rect 13542 11872 13598 11928
rect 13542 11620 13598 11656
rect 13542 11600 13544 11620
rect 13544 11600 13596 11620
rect 13596 11600 13598 11620
rect 13266 11056 13322 11112
rect 13542 10804 13598 10840
rect 13542 10784 13544 10804
rect 13544 10784 13596 10804
rect 13596 10784 13598 10804
rect 13174 9016 13230 9072
rect 13542 9016 13598 9072
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 11702 7268 11758 7304
rect 11702 7248 11704 7268
rect 11704 7248 11756 7268
rect 11756 7248 11758 7268
rect 10874 6296 10930 6352
rect 11334 6024 11390 6080
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 10230 5208 10286 5264
rect 10230 4936 10286 4992
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 9770 3848 9826 3904
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 11886 4936 11942 4992
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 12622 7812 12678 7848
rect 12622 7792 12624 7812
rect 12624 7792 12676 7812
rect 12676 7792 12678 7812
rect 12806 6976 12862 7032
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 16486 20304 16542 20360
rect 18234 20304 18290 20360
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 18602 19896 18658 19952
rect 17498 19780 17554 19816
rect 17498 19760 17500 19780
rect 17500 19760 17552 19780
rect 17552 19760 17554 19780
rect 14186 7656 14242 7712
rect 14278 5908 14334 5944
rect 14278 5888 14280 5908
rect 14280 5888 14332 5908
rect 14332 5888 14334 5908
rect 12346 3984 12402 4040
rect 13082 4276 13138 4312
rect 13082 4256 13084 4276
rect 13084 4256 13136 4276
rect 13136 4256 13138 4276
rect 12254 3440 12310 3496
rect 11610 2760 11666 2816
rect 14370 4528 14426 4584
rect 12070 2896 12126 2952
rect 13818 2896 13874 2952
rect 13910 2760 13966 2816
rect 14278 3032 14334 3088
rect 14370 2896 14426 2952
rect 14462 2760 14518 2816
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 15750 17040 15806 17096
rect 15290 5480 15346 5536
rect 15290 4256 15346 4312
rect 14554 2488 14610 2544
rect 15658 9832 15714 9888
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 17682 13096 17738 13152
rect 16394 11736 16450 11792
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 16486 9696 16542 9752
rect 16394 9560 16450 9616
rect 16210 9152 16266 9208
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 15750 6704 15806 6760
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 16486 6316 16542 6352
rect 16486 6296 16488 6316
rect 16488 6296 16540 6316
rect 16540 6296 16542 6316
rect 16302 5616 16358 5672
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 16486 5480 16542 5536
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 16762 5208 16818 5264
rect 16854 4528 16910 4584
rect 17314 10004 17316 10024
rect 17316 10004 17368 10024
rect 17368 10004 17370 10024
rect 17314 9968 17370 10004
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 19430 20596 19486 20632
rect 19430 20576 19432 20596
rect 19432 20576 19484 20596
rect 19484 20576 19486 20596
rect 18786 19352 18842 19408
rect 18694 12416 18750 12472
rect 18418 12280 18474 12336
rect 17774 10668 17830 10704
rect 17774 10648 17776 10668
rect 17776 10648 17828 10668
rect 17828 10648 17830 10668
rect 17958 10648 18014 10704
rect 18050 9152 18106 9208
rect 18418 10412 18420 10432
rect 18420 10412 18472 10432
rect 18472 10412 18474 10432
rect 18418 10376 18474 10412
rect 18418 9696 18474 9752
rect 18510 9580 18566 9616
rect 18510 9560 18512 9580
rect 18512 9560 18564 9580
rect 18564 9560 18566 9580
rect 17314 5344 17370 5400
rect 17682 6432 17738 6488
rect 17498 6024 17554 6080
rect 17406 5072 17462 5128
rect 17314 4800 17370 4856
rect 17130 4664 17186 4720
rect 16946 3576 17002 3632
rect 15474 2624 15530 2680
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 17866 5888 17922 5944
rect 17774 4972 17776 4992
rect 17776 4972 17828 4992
rect 17828 4972 17830 4992
rect 17774 4936 17830 4972
rect 17498 3032 17554 3088
rect 18326 8492 18382 8528
rect 18326 8472 18328 8492
rect 18328 8472 18380 8492
rect 18380 8472 18382 8492
rect 18418 7928 18474 7984
rect 18050 5480 18106 5536
rect 18510 4392 18566 4448
rect 18970 15000 19026 15056
rect 19062 12416 19118 12472
rect 18878 7384 18934 7440
rect 18786 4120 18842 4176
rect 16946 2760 17002 2816
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 19706 19780 19762 19816
rect 19706 19760 19708 19780
rect 19708 19760 19760 19780
rect 19760 19760 19762 19780
rect 19338 15988 19340 16008
rect 19340 15988 19392 16008
rect 19392 15988 19394 16008
rect 19338 15952 19394 15988
rect 19338 12416 19394 12472
rect 19246 9696 19302 9752
rect 19154 9560 19210 9616
rect 20626 20476 20628 20496
rect 20628 20476 20680 20496
rect 20680 20476 20682 20496
rect 20626 20440 20682 20476
rect 23202 20576 23258 20632
rect 23846 20476 23848 20496
rect 23848 20476 23900 20496
rect 23900 20476 23902 20496
rect 23846 20440 23902 20476
rect 21730 20304 21786 20360
rect 22006 20304 22062 20360
rect 23662 20340 23664 20360
rect 23664 20340 23716 20360
rect 23716 20340 23718 20360
rect 21914 20204 21916 20224
rect 21916 20204 21968 20224
rect 21968 20204 21970 20224
rect 21914 20168 21970 20204
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 21546 19896 21602 19952
rect 20074 12416 20130 12472
rect 19246 6296 19302 6352
rect 19154 3984 19210 4040
rect 18418 3576 18474 3632
rect 19062 3576 19118 3632
rect 1674 312 1730 368
rect 19430 2624 19486 2680
rect 19154 2352 19210 2408
rect 18510 1400 18566 1456
rect 19614 8608 19670 8664
rect 19890 8336 19946 8392
rect 19614 3440 19670 3496
rect 20166 2352 20222 2408
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 21362 15816 21418 15872
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 21362 14592 21418 14648
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 23662 20304 23718 20340
rect 24858 22344 24914 22400
rect 24674 19760 24730 19816
rect 25042 19352 25098 19408
rect 25042 14864 25098 14920
rect 25042 13912 25098 13968
rect 25410 20032 25466 20088
rect 25410 14320 25466 14376
rect 25318 12960 25374 13016
rect 25318 12824 25374 12880
rect 25042 7928 25098 7984
rect 23018 2760 23074 2816
rect 22834 2508 22890 2544
rect 22834 2488 22836 2508
rect 22836 2488 22888 2508
rect 22888 2488 22890 2508
rect 25686 23024 25742 23080
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25686 21528 25742 21584
rect 25778 21256 25834 21312
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 25594 20304 25650 20360
rect 25502 11600 25558 11656
rect 29182 20440 29238 20496
rect 27710 20168 27766 20224
rect 26330 19896 26386 19952
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25778 17040 25834 17096
rect 25686 16088 25742 16144
rect 25686 13368 25742 13424
rect 25594 9696 25650 9752
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25870 15408 25926 15464
rect 25778 8608 25834 8664
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 27526 14456 27582 14512
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 26146 12688 26202 12744
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 26606 11600 26662 11656
rect 26422 11056 26478 11112
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 26698 11076 26754 11112
rect 26698 11056 26700 11076
rect 26700 11056 26752 11076
rect 26752 11056 26754 11076
rect 26330 10648 26386 10704
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 25318 6432 25374 6488
rect 24398 5344 24454 5400
rect 25870 6704 25926 6760
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 25778 5208 25834 5264
rect 24398 4936 24454 4992
rect 25686 4392 25742 4448
rect 24214 4120 24270 4176
rect 25318 3984 25374 4040
rect 25134 3576 25190 3632
rect 25502 3032 25558 3088
rect 25042 2896 25098 2952
rect 25226 2760 25282 2816
rect 25502 2796 25504 2816
rect 25504 2796 25556 2816
rect 25556 2796 25558 2816
rect 25502 2760 25558 2796
rect 24582 2352 24638 2408
rect 24766 1672 24822 1728
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 26698 10376 26754 10432
rect 26698 9832 26754 9888
rect 26514 9460 26516 9480
rect 26516 9460 26568 9480
rect 26568 9460 26570 9480
rect 26514 9424 26570 9460
rect 26606 9288 26662 9344
rect 26422 9016 26478 9072
rect 26514 8880 26570 8936
rect 26698 8608 26754 8664
rect 26514 8336 26570 8392
rect 27710 8336 27766 8392
rect 26698 7384 26754 7440
rect 26606 6976 26662 7032
rect 26698 6296 26754 6352
rect 26514 6196 26516 6216
rect 26516 6196 26568 6216
rect 26568 6196 26570 6216
rect 26514 6160 26570 6196
rect 26514 5772 26570 5808
rect 26514 5752 26516 5772
rect 26516 5752 26568 5772
rect 26568 5752 26570 5772
rect 26606 5616 26662 5672
rect 26698 5072 26754 5128
rect 26790 4936 26846 4992
rect 26514 4684 26570 4720
rect 26514 4664 26516 4684
rect 26516 4664 26568 4684
rect 26568 4664 26570 4684
rect 26422 4528 26478 4584
rect 26330 3440 26386 3496
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 25870 1944 25926 2000
rect 26606 4392 26662 4448
rect 26698 3848 26754 3904
rect 26606 3304 26662 3360
rect 27342 3032 27398 3088
rect 27066 2644 27122 2680
rect 27066 2624 27068 2644
rect 27068 2624 27120 2644
rect 27120 2624 27122 2644
rect 27526 2932 27528 2952
rect 27528 2932 27580 2952
rect 27580 2932 27582 2952
rect 27526 2896 27582 2932
rect 28354 2760 28410 2816
rect 27710 856 27766 912
rect 29366 1672 29422 1728
rect 18326 312 18382 368
<< metal3 >>
rect 0 23626 480 23656
rect 2957 23626 3023 23629
rect 0 23624 3023 23626
rect 0 23568 2962 23624
rect 3018 23568 3023 23624
rect 0 23566 3023 23568
rect 0 23536 480 23566
rect 2957 23563 3023 23566
rect 25497 23626 25563 23629
rect 29520 23626 30000 23656
rect 25497 23624 30000 23626
rect 25497 23568 25502 23624
rect 25558 23568 30000 23624
rect 25497 23566 30000 23568
rect 25497 23563 25563 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 2773 23082 2839 23085
rect 0 23080 2839 23082
rect 0 23024 2778 23080
rect 2834 23024 2839 23080
rect 0 23022 2839 23024
rect 0 22992 480 23022
rect 2773 23019 2839 23022
rect 25681 23082 25747 23085
rect 29520 23082 30000 23112
rect 25681 23080 30000 23082
rect 25681 23024 25686 23080
rect 25742 23024 30000 23080
rect 25681 23022 30000 23024
rect 25681 23019 25747 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 4061 22402 4127 22405
rect 0 22400 4127 22402
rect 0 22344 4066 22400
rect 4122 22344 4127 22400
rect 0 22342 4127 22344
rect 0 22312 480 22342
rect 4061 22339 4127 22342
rect 24853 22402 24919 22405
rect 29520 22402 30000 22432
rect 24853 22400 30000 22402
rect 24853 22344 24858 22400
rect 24914 22344 30000 22400
rect 24853 22342 30000 22344
rect 24853 22339 24919 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 3969 21858 4035 21861
rect 29520 21858 30000 21888
rect 0 21856 4035 21858
rect 0 21800 3974 21856
rect 4030 21800 4035 21856
rect 0 21798 4035 21800
rect 0 21768 480 21798
rect 3969 21795 4035 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 25681 21586 25747 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 25681 21584 26434 21586
rect 25681 21528 25686 21584
rect 25742 21528 26434 21584
rect 25681 21526 26434 21528
rect 25681 21523 25747 21526
rect 0 21314 480 21344
rect 3877 21314 3943 21317
rect 0 21312 3943 21314
rect 0 21256 3882 21312
rect 3938 21256 3943 21312
rect 0 21254 3943 21256
rect 0 21224 480 21254
rect 3877 21251 3943 21254
rect 25773 21314 25839 21317
rect 29520 21314 30000 21344
rect 25773 21312 30000 21314
rect 25773 21256 25778 21312
rect 25834 21256 30000 21312
rect 25773 21254 30000 21256
rect 25773 21251 25839 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 3877 20634 3943 20637
rect 0 20632 3943 20634
rect 0 20576 3882 20632
rect 3938 20576 3943 20632
rect 0 20574 3943 20576
rect 0 20544 480 20574
rect 3877 20571 3943 20574
rect 19425 20634 19491 20637
rect 23197 20634 23263 20637
rect 29520 20634 30000 20664
rect 19425 20632 23263 20634
rect 19425 20576 19430 20632
rect 19486 20576 23202 20632
rect 23258 20576 23263 20632
rect 19425 20574 23263 20576
rect 19425 20571 19491 20574
rect 23197 20571 23263 20574
rect 29318 20574 30000 20634
rect 6729 20498 6795 20501
rect 20621 20498 20687 20501
rect 6729 20496 20687 20498
rect 6729 20440 6734 20496
rect 6790 20440 20626 20496
rect 20682 20440 20687 20496
rect 6729 20438 20687 20440
rect 6729 20435 6795 20438
rect 20621 20435 20687 20438
rect 23841 20498 23907 20501
rect 29177 20498 29243 20501
rect 23841 20496 29243 20498
rect 23841 20440 23846 20496
rect 23902 20440 29182 20496
rect 29238 20440 29243 20496
rect 23841 20438 29243 20440
rect 23841 20435 23907 20438
rect 29177 20435 29243 20438
rect 749 20362 815 20365
rect 16481 20362 16547 20365
rect 749 20360 16547 20362
rect 749 20304 754 20360
rect 810 20304 16486 20360
rect 16542 20304 16547 20360
rect 749 20302 16547 20304
rect 749 20299 815 20302
rect 16481 20299 16547 20302
rect 18229 20362 18295 20365
rect 21725 20362 21791 20365
rect 18229 20360 21791 20362
rect 18229 20304 18234 20360
rect 18290 20304 21730 20360
rect 21786 20304 21791 20360
rect 18229 20302 21791 20304
rect 18229 20299 18295 20302
rect 21725 20299 21791 20302
rect 22001 20362 22067 20365
rect 23657 20362 23723 20365
rect 22001 20360 23723 20362
rect 22001 20304 22006 20360
rect 22062 20304 23662 20360
rect 23718 20304 23723 20360
rect 22001 20302 23723 20304
rect 22001 20299 22067 20302
rect 23657 20299 23723 20302
rect 25589 20362 25655 20365
rect 29318 20362 29378 20574
rect 29520 20544 30000 20574
rect 25589 20360 29378 20362
rect 25589 20304 25594 20360
rect 25650 20304 29378 20360
rect 25589 20302 29378 20304
rect 25589 20299 25655 20302
rect 21909 20226 21975 20229
rect 27705 20226 27771 20229
rect 21909 20224 27771 20226
rect 21909 20168 21914 20224
rect 21970 20168 27710 20224
rect 27766 20168 27771 20224
rect 21909 20166 27771 20168
rect 21909 20163 21975 20166
rect 27705 20163 27771 20166
rect 10944 20160 11264 20161
rect 0 20090 480 20120
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 4061 20090 4127 20093
rect 0 20088 4127 20090
rect 0 20032 4066 20088
rect 4122 20032 4127 20088
rect 0 20030 4127 20032
rect 0 20000 480 20030
rect 4061 20027 4127 20030
rect 25405 20090 25471 20093
rect 29520 20090 30000 20120
rect 25405 20088 30000 20090
rect 25405 20032 25410 20088
rect 25466 20032 30000 20088
rect 25405 20030 30000 20032
rect 25405 20027 25471 20030
rect 29520 20000 30000 20030
rect 3693 19954 3759 19957
rect 18597 19954 18663 19957
rect 3693 19952 18663 19954
rect 3693 19896 3698 19952
rect 3754 19896 18602 19952
rect 18658 19896 18663 19952
rect 3693 19894 18663 19896
rect 3693 19891 3759 19894
rect 18597 19891 18663 19894
rect 21541 19954 21607 19957
rect 26325 19954 26391 19957
rect 21541 19952 26391 19954
rect 21541 19896 21546 19952
rect 21602 19896 26330 19952
rect 26386 19896 26391 19952
rect 21541 19894 26391 19896
rect 21541 19891 21607 19894
rect 26325 19891 26391 19894
rect 2221 19818 2287 19821
rect 17493 19818 17559 19821
rect 2221 19816 17559 19818
rect 2221 19760 2226 19816
rect 2282 19760 17498 19816
rect 17554 19760 17559 19816
rect 2221 19758 17559 19760
rect 2221 19755 2287 19758
rect 17493 19755 17559 19758
rect 19701 19818 19767 19821
rect 24669 19818 24735 19821
rect 19701 19816 24735 19818
rect 19701 19760 19706 19816
rect 19762 19760 24674 19816
rect 24730 19760 24735 19816
rect 19701 19758 24735 19760
rect 19701 19755 19767 19758
rect 24669 19755 24735 19758
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 0 19410 480 19440
rect 2773 19410 2839 19413
rect 0 19408 2839 19410
rect 0 19352 2778 19408
rect 2834 19352 2839 19408
rect 0 19350 2839 19352
rect 0 19320 480 19350
rect 2773 19347 2839 19350
rect 12709 19410 12775 19413
rect 18781 19410 18847 19413
rect 12709 19408 18847 19410
rect 12709 19352 12714 19408
rect 12770 19352 18786 19408
rect 18842 19352 18847 19408
rect 12709 19350 18847 19352
rect 12709 19347 12775 19350
rect 18781 19347 18847 19350
rect 25037 19410 25103 19413
rect 29520 19410 30000 19440
rect 25037 19408 30000 19410
rect 25037 19352 25042 19408
rect 25098 19352 30000 19408
rect 25037 19350 30000 19352
rect 25037 19347 25103 19350
rect 29520 19320 30000 19350
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 0 18866 480 18896
rect 9213 18866 9279 18869
rect 0 18864 9279 18866
rect 0 18808 9218 18864
rect 9274 18808 9279 18864
rect 0 18806 9279 18808
rect 0 18776 480 18806
rect 9213 18803 9279 18806
rect 12065 18866 12131 18869
rect 29520 18866 30000 18896
rect 12065 18864 30000 18866
rect 12065 18808 12070 18864
rect 12126 18808 30000 18864
rect 12065 18806 30000 18808
rect 12065 18803 12131 18806
rect 29520 18776 30000 18806
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 0 18322 480 18352
rect 3417 18322 3483 18325
rect 0 18320 3483 18322
rect 0 18264 3422 18320
rect 3478 18264 3483 18320
rect 0 18262 3483 18264
rect 0 18232 480 18262
rect 3417 18259 3483 18262
rect 3693 18322 3759 18325
rect 29520 18322 30000 18352
rect 3693 18320 30000 18322
rect 3693 18264 3698 18320
rect 3754 18264 30000 18320
rect 3693 18262 30000 18264
rect 3693 18259 3759 18262
rect 29520 18232 30000 18262
rect 12525 18186 12591 18189
rect 11838 18184 12591 18186
rect 11838 18128 12530 18184
rect 12586 18128 12591 18184
rect 11838 18126 12591 18128
rect 11838 18050 11898 18126
rect 12525 18123 12591 18126
rect 11973 18050 12039 18053
rect 11838 18048 12039 18050
rect 11838 17992 11978 18048
rect 12034 17992 12039 18048
rect 11838 17990 12039 17992
rect 11973 17987 12039 17990
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 13445 17778 13511 17781
rect 13445 17776 29378 17778
rect 13445 17720 13450 17776
rect 13506 17720 29378 17776
rect 13445 17718 29378 17720
rect 13445 17715 13511 17718
rect 0 17642 480 17672
rect 29318 17642 29378 17718
rect 29520 17642 30000 17672
rect 0 17582 674 17642
rect 29318 17582 30000 17642
rect 0 17552 480 17582
rect 614 17506 674 17582
rect 29520 17552 30000 17582
rect 614 17446 5826 17506
rect 0 17098 480 17128
rect 5766 17098 5826 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 15745 17098 15811 17101
rect 0 17038 4170 17098
rect 5766 17096 15811 17098
rect 5766 17040 15750 17096
rect 15806 17040 15811 17096
rect 5766 17038 15811 17040
rect 0 17008 480 17038
rect 4110 16962 4170 17038
rect 15745 17035 15811 17038
rect 25773 17098 25839 17101
rect 29520 17098 30000 17128
rect 25773 17096 30000 17098
rect 25773 17040 25778 17096
rect 25834 17040 30000 17096
rect 25773 17038 30000 17040
rect 25773 17035 25839 17038
rect 29520 17008 30000 17038
rect 7833 16962 7899 16965
rect 4110 16960 7899 16962
rect 4110 16904 7838 16960
rect 7894 16904 7899 16960
rect 4110 16902 7899 16904
rect 7833 16899 7899 16902
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 9489 16554 9555 16557
rect 4110 16552 9555 16554
rect 4110 16496 9494 16552
rect 9550 16496 9555 16552
rect 4110 16494 9555 16496
rect 0 16418 480 16448
rect 4110 16418 4170 16494
rect 9489 16491 9555 16494
rect 29520 16418 30000 16448
rect 0 16358 4170 16418
rect 26374 16358 30000 16418
rect 0 16328 480 16358
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 25681 16146 25747 16149
rect 26374 16146 26434 16358
rect 29520 16328 30000 16358
rect 25681 16144 26434 16146
rect 25681 16088 25686 16144
rect 25742 16088 26434 16144
rect 25681 16086 26434 16088
rect 25681 16083 25747 16086
rect 4613 16010 4679 16013
rect 19333 16010 19399 16013
rect 4613 16008 19399 16010
rect 4613 15952 4618 16008
rect 4674 15952 19338 16008
rect 19394 15952 19399 16008
rect 4613 15950 19399 15952
rect 4613 15947 4679 15950
rect 19333 15947 19399 15950
rect 0 15874 480 15904
rect 4337 15874 4403 15877
rect 0 15872 4403 15874
rect 0 15816 4342 15872
rect 4398 15816 4403 15872
rect 0 15814 4403 15816
rect 0 15784 480 15814
rect 4337 15811 4403 15814
rect 21357 15874 21423 15877
rect 29520 15874 30000 15904
rect 21357 15872 30000 15874
rect 21357 15816 21362 15872
rect 21418 15816 30000 15872
rect 21357 15814 30000 15816
rect 21357 15811 21423 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 25865 15466 25931 15469
rect 25865 15464 26434 15466
rect 25865 15408 25870 15464
rect 25926 15408 26434 15464
rect 25865 15406 26434 15408
rect 25865 15403 25931 15406
rect 0 15330 480 15360
rect 2957 15330 3023 15333
rect 0 15328 3023 15330
rect 0 15272 2962 15328
rect 3018 15272 3023 15328
rect 0 15270 3023 15272
rect 26374 15330 26434 15406
rect 29520 15330 30000 15360
rect 26374 15270 30000 15330
rect 0 15240 480 15270
rect 2957 15267 3023 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 3877 15058 3943 15061
rect 18965 15058 19031 15061
rect 3877 15056 19031 15058
rect 3877 15000 3882 15056
rect 3938 15000 18970 15056
rect 19026 15000 19031 15056
rect 3877 14998 19031 15000
rect 3877 14995 3943 14998
rect 18965 14995 19031 14998
rect 3509 14922 3575 14925
rect 25037 14922 25103 14925
rect 3509 14920 25103 14922
rect 3509 14864 3514 14920
rect 3570 14864 25042 14920
rect 25098 14864 25103 14920
rect 3509 14862 25103 14864
rect 3509 14859 3575 14862
rect 25037 14859 25103 14862
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 2313 14650 2379 14653
rect 0 14648 2379 14650
rect 0 14592 2318 14648
rect 2374 14592 2379 14648
rect 0 14590 2379 14592
rect 0 14560 480 14590
rect 2313 14587 2379 14590
rect 21357 14650 21423 14653
rect 29520 14650 30000 14680
rect 21357 14648 30000 14650
rect 21357 14592 21362 14648
rect 21418 14592 30000 14648
rect 21357 14590 30000 14592
rect 21357 14587 21423 14590
rect 29520 14560 30000 14590
rect 4061 14514 4127 14517
rect 11789 14514 11855 14517
rect 27521 14514 27587 14517
rect 4061 14512 27587 14514
rect 4061 14456 4066 14512
rect 4122 14456 11794 14512
rect 11850 14456 27526 14512
rect 27582 14456 27587 14512
rect 4061 14454 27587 14456
rect 4061 14451 4127 14454
rect 11789 14451 11855 14454
rect 27521 14451 27587 14454
rect 13997 14378 14063 14381
rect 25405 14378 25471 14381
rect 13997 14376 25471 14378
rect 13997 14320 14002 14376
rect 14058 14320 25410 14376
rect 25466 14320 25471 14376
rect 13997 14318 25471 14320
rect 13997 14315 14063 14318
rect 25405 14315 25471 14318
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 3233 14106 3299 14109
rect 29520 14106 30000 14136
rect 0 14104 3299 14106
rect 0 14048 3238 14104
rect 3294 14048 3299 14104
rect 0 14046 3299 14048
rect 0 14016 480 14046
rect 3233 14043 3299 14046
rect 26374 14046 30000 14106
rect 25037 13970 25103 13973
rect 26374 13970 26434 14046
rect 29520 14016 30000 14046
rect 25037 13968 26434 13970
rect 25037 13912 25042 13968
rect 25098 13912 26434 13968
rect 25037 13910 26434 13912
rect 25037 13907 25103 13910
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 0 13426 480 13456
rect 3693 13426 3759 13429
rect 0 13424 3759 13426
rect 0 13368 3698 13424
rect 3754 13368 3759 13424
rect 0 13366 3759 13368
rect 0 13336 480 13366
rect 3693 13363 3759 13366
rect 12893 13426 12959 13429
rect 25681 13426 25747 13429
rect 29520 13426 30000 13456
rect 12893 13424 25747 13426
rect 12893 13368 12898 13424
rect 12954 13368 25686 13424
rect 25742 13368 25747 13424
rect 12893 13366 25747 13368
rect 12893 13363 12959 13366
rect 25681 13363 25747 13366
rect 25822 13366 30000 13426
rect 1485 13290 1551 13293
rect 11789 13290 11855 13293
rect 1485 13288 11855 13290
rect 1485 13232 1490 13288
rect 1546 13232 11794 13288
rect 11850 13232 11855 13288
rect 1485 13230 11855 13232
rect 1485 13227 1551 13230
rect 11789 13227 11855 13230
rect 17677 13154 17743 13157
rect 25822 13154 25882 13366
rect 29520 13336 30000 13366
rect 17677 13152 25882 13154
rect 17677 13096 17682 13152
rect 17738 13096 25882 13152
rect 17677 13094 25882 13096
rect 17677 13091 17743 13094
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 25313 13018 25379 13021
rect 17174 13016 25379 13018
rect 17174 12960 25318 13016
rect 25374 12960 25379 13016
rect 17174 12958 25379 12960
rect 0 12882 480 12912
rect 3509 12882 3575 12885
rect 0 12880 3575 12882
rect 0 12824 3514 12880
rect 3570 12824 3575 12880
rect 0 12822 3575 12824
rect 0 12792 480 12822
rect 3509 12819 3575 12822
rect 5073 12882 5139 12885
rect 17174 12882 17234 12958
rect 25313 12955 25379 12958
rect 5073 12880 17234 12882
rect 5073 12824 5078 12880
rect 5134 12824 17234 12880
rect 5073 12822 17234 12824
rect 25313 12882 25379 12885
rect 29520 12882 30000 12912
rect 25313 12880 30000 12882
rect 25313 12824 25318 12880
rect 25374 12824 30000 12880
rect 25313 12822 30000 12824
rect 5073 12819 5139 12822
rect 25313 12819 25379 12822
rect 29520 12792 30000 12822
rect 3325 12746 3391 12749
rect 26141 12746 26207 12749
rect 3325 12744 26207 12746
rect 3325 12688 3330 12744
rect 3386 12688 26146 12744
rect 26202 12688 26207 12744
rect 3325 12686 26207 12688
rect 3325 12683 3391 12686
rect 26141 12683 26207 12686
rect 3785 12610 3851 12613
rect 3969 12610 4035 12613
rect 3785 12608 4035 12610
rect 3785 12552 3790 12608
rect 3846 12552 3974 12608
rect 4030 12552 4035 12608
rect 3785 12550 4035 12552
rect 3785 12547 3851 12550
rect 3969 12547 4035 12550
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 3325 12474 3391 12477
rect 3785 12474 3851 12477
rect 3325 12472 3851 12474
rect 3325 12416 3330 12472
rect 3386 12416 3790 12472
rect 3846 12416 3851 12472
rect 3325 12414 3851 12416
rect 3325 12411 3391 12414
rect 3785 12411 3851 12414
rect 18689 12474 18755 12477
rect 19057 12474 19123 12477
rect 18689 12472 19123 12474
rect 18689 12416 18694 12472
rect 18750 12416 19062 12472
rect 19118 12416 19123 12472
rect 18689 12414 19123 12416
rect 18689 12411 18755 12414
rect 19057 12411 19123 12414
rect 19333 12474 19399 12477
rect 20069 12474 20135 12477
rect 19333 12472 20135 12474
rect 19333 12416 19338 12472
rect 19394 12416 20074 12472
rect 20130 12416 20135 12472
rect 19333 12414 20135 12416
rect 19333 12411 19399 12414
rect 20069 12411 20135 12414
rect 0 12338 480 12368
rect 2037 12338 2103 12341
rect 7189 12338 7255 12341
rect 0 12278 1226 12338
rect 0 12248 480 12278
rect 1166 12066 1226 12278
rect 2037 12336 7255 12338
rect 2037 12280 2042 12336
rect 2098 12280 7194 12336
rect 7250 12280 7255 12336
rect 2037 12278 7255 12280
rect 2037 12275 2103 12278
rect 7189 12275 7255 12278
rect 18413 12338 18479 12341
rect 29520 12338 30000 12368
rect 18413 12336 30000 12338
rect 18413 12280 18418 12336
rect 18474 12280 30000 12336
rect 18413 12278 30000 12280
rect 18413 12275 18479 12278
rect 29520 12248 30000 12278
rect 3509 12202 3575 12205
rect 9397 12202 9463 12205
rect 3509 12200 9463 12202
rect 3509 12144 3514 12200
rect 3570 12144 9402 12200
rect 9458 12144 9463 12200
rect 3509 12142 9463 12144
rect 3509 12139 3575 12142
rect 9397 12139 9463 12142
rect 3049 12066 3115 12069
rect 1166 12064 3115 12066
rect 1166 12008 3054 12064
rect 3110 12008 3115 12064
rect 1166 12006 3115 12008
rect 3049 12003 3115 12006
rect 6729 12066 6795 12069
rect 7649 12066 7715 12069
rect 6729 12064 7715 12066
rect 6729 12008 6734 12064
rect 6790 12008 7654 12064
rect 7710 12008 7715 12064
rect 6729 12006 7715 12008
rect 6729 12003 6795 12006
rect 7649 12003 7715 12006
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 13537 11930 13603 11933
rect 7606 11928 13603 11930
rect 7606 11872 13542 11928
rect 13598 11872 13603 11928
rect 7606 11870 13603 11872
rect 2681 11794 2747 11797
rect 7606 11794 7666 11870
rect 13537 11867 13603 11870
rect 2681 11792 7666 11794
rect 2681 11736 2686 11792
rect 2742 11736 7666 11792
rect 2681 11734 7666 11736
rect 12341 11794 12407 11797
rect 16389 11794 16455 11797
rect 12341 11792 16455 11794
rect 12341 11736 12346 11792
rect 12402 11736 16394 11792
rect 16450 11736 16455 11792
rect 12341 11734 16455 11736
rect 2681 11731 2747 11734
rect 12341 11731 12407 11734
rect 16389 11731 16455 11734
rect 0 11658 480 11688
rect 1577 11658 1643 11661
rect 0 11656 1643 11658
rect 0 11600 1582 11656
rect 1638 11600 1643 11656
rect 0 11598 1643 11600
rect 0 11568 480 11598
rect 1577 11595 1643 11598
rect 3233 11658 3299 11661
rect 9029 11658 9095 11661
rect 3233 11656 9095 11658
rect 3233 11600 3238 11656
rect 3294 11600 9034 11656
rect 9090 11600 9095 11656
rect 3233 11598 9095 11600
rect 3233 11595 3299 11598
rect 9029 11595 9095 11598
rect 13537 11658 13603 11661
rect 25497 11658 25563 11661
rect 13537 11656 25563 11658
rect 13537 11600 13542 11656
rect 13598 11600 25502 11656
rect 25558 11600 25563 11656
rect 13537 11598 25563 11600
rect 13537 11595 13603 11598
rect 25497 11595 25563 11598
rect 26601 11658 26667 11661
rect 29520 11658 30000 11688
rect 26601 11656 30000 11658
rect 26601 11600 26606 11656
rect 26662 11600 30000 11656
rect 26601 11598 30000 11600
rect 26601 11595 26667 11598
rect 29520 11568 30000 11598
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 0 11114 480 11144
rect 1577 11114 1643 11117
rect 0 11112 1643 11114
rect 0 11056 1582 11112
rect 1638 11056 1643 11112
rect 0 11054 1643 11056
rect 0 11024 480 11054
rect 1577 11051 1643 11054
rect 3233 11114 3299 11117
rect 11697 11114 11763 11117
rect 3233 11112 11763 11114
rect 3233 11056 3238 11112
rect 3294 11056 11702 11112
rect 11758 11056 11763 11112
rect 3233 11054 11763 11056
rect 3233 11051 3299 11054
rect 11697 11051 11763 11054
rect 13261 11114 13327 11117
rect 26417 11114 26483 11117
rect 13261 11112 26483 11114
rect 13261 11056 13266 11112
rect 13322 11056 26422 11112
rect 26478 11056 26483 11112
rect 13261 11054 26483 11056
rect 13261 11051 13327 11054
rect 26417 11051 26483 11054
rect 26693 11114 26759 11117
rect 29520 11114 30000 11144
rect 26693 11112 30000 11114
rect 26693 11056 26698 11112
rect 26754 11056 30000 11112
rect 26693 11054 30000 11056
rect 26693 11051 26759 11054
rect 29520 11024 30000 11054
rect 9622 10916 9628 10980
rect 9692 10978 9698 10980
rect 11973 10978 12039 10981
rect 9692 10976 12039 10978
rect 9692 10920 11978 10976
rect 12034 10920 12039 10976
rect 9692 10918 12039 10920
rect 9692 10916 9698 10918
rect 11973 10915 12039 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 2037 10842 2103 10845
rect 4429 10842 4495 10845
rect 2037 10840 4495 10842
rect 2037 10784 2042 10840
rect 2098 10784 4434 10840
rect 4490 10784 4495 10840
rect 2037 10782 4495 10784
rect 2037 10779 2103 10782
rect 4429 10779 4495 10782
rect 7557 10842 7623 10845
rect 13537 10842 13603 10845
rect 7557 10840 13603 10842
rect 7557 10784 7562 10840
rect 7618 10784 13542 10840
rect 13598 10784 13603 10840
rect 7557 10782 13603 10784
rect 7557 10779 7623 10782
rect 13537 10779 13603 10782
rect 3049 10706 3115 10709
rect 4797 10706 4863 10709
rect 17769 10706 17835 10709
rect 3049 10704 17835 10706
rect 3049 10648 3054 10704
rect 3110 10648 4802 10704
rect 4858 10648 17774 10704
rect 17830 10648 17835 10704
rect 3049 10646 17835 10648
rect 3049 10643 3115 10646
rect 4797 10643 4863 10646
rect 17769 10643 17835 10646
rect 17953 10706 18019 10709
rect 26325 10706 26391 10709
rect 17953 10704 26391 10706
rect 17953 10648 17958 10704
rect 18014 10648 26330 10704
rect 26386 10648 26391 10704
rect 17953 10646 26391 10648
rect 17953 10643 18019 10646
rect 26325 10643 26391 10646
rect 2497 10570 2563 10573
rect 7557 10570 7623 10573
rect 2497 10568 7623 10570
rect 2497 10512 2502 10568
rect 2558 10512 7562 10568
rect 7618 10512 7623 10568
rect 2497 10510 7623 10512
rect 2497 10507 2563 10510
rect 7557 10507 7623 10510
rect 7790 10510 12312 10570
rect 0 10434 480 10464
rect 1577 10434 1643 10437
rect 0 10432 1643 10434
rect 0 10376 1582 10432
rect 1638 10376 1643 10432
rect 0 10374 1643 10376
rect 0 10344 480 10374
rect 1577 10371 1643 10374
rect 4521 10434 4587 10437
rect 7790 10434 7850 10510
rect 4521 10432 7850 10434
rect 4521 10376 4526 10432
rect 4582 10376 7850 10432
rect 4521 10374 7850 10376
rect 12252 10434 12312 10510
rect 18413 10434 18479 10437
rect 12252 10432 18479 10434
rect 12252 10376 18418 10432
rect 18474 10376 18479 10432
rect 12252 10374 18479 10376
rect 4521 10371 4587 10374
rect 18413 10371 18479 10374
rect 26693 10434 26759 10437
rect 29520 10434 30000 10464
rect 26693 10432 30000 10434
rect 26693 10376 26698 10432
rect 26754 10376 30000 10432
rect 26693 10374 30000 10376
rect 26693 10371 26759 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 3417 10298 3483 10301
rect 8150 10298 8156 10300
rect 3417 10296 8156 10298
rect 3417 10240 3422 10296
rect 3478 10240 8156 10296
rect 3417 10238 8156 10240
rect 3417 10235 3483 10238
rect 8150 10236 8156 10238
rect 8220 10236 8226 10300
rect 4245 10162 4311 10165
rect 9622 10162 9628 10164
rect 4245 10160 9628 10162
rect 4245 10104 4250 10160
rect 4306 10104 9628 10160
rect 4245 10102 9628 10104
rect 4245 10099 4311 10102
rect 9622 10100 9628 10102
rect 9692 10100 9698 10164
rect 8150 9964 8156 10028
rect 8220 10026 8226 10028
rect 17309 10026 17375 10029
rect 8220 10024 17375 10026
rect 8220 9968 17314 10024
rect 17370 9968 17375 10024
rect 8220 9966 17375 9968
rect 8220 9964 8226 9966
rect 17309 9963 17375 9966
rect 0 9890 480 9920
rect 1577 9890 1643 9893
rect 0 9888 1643 9890
rect 0 9832 1582 9888
rect 1638 9832 1643 9888
rect 0 9830 1643 9832
rect 0 9800 480 9830
rect 1577 9827 1643 9830
rect 7833 9890 7899 9893
rect 15653 9890 15719 9893
rect 7833 9888 15719 9890
rect 7833 9832 7838 9888
rect 7894 9832 15658 9888
rect 15714 9832 15719 9888
rect 7833 9830 15719 9832
rect 7833 9827 7899 9830
rect 15653 9827 15719 9830
rect 26693 9890 26759 9893
rect 29520 9890 30000 9920
rect 26693 9888 30000 9890
rect 26693 9832 26698 9888
rect 26754 9832 30000 9888
rect 26693 9830 30000 9832
rect 26693 9827 26759 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 7465 9754 7531 9757
rect 10041 9754 10107 9757
rect 7465 9752 10107 9754
rect 7465 9696 7470 9752
rect 7526 9696 10046 9752
rect 10102 9696 10107 9752
rect 7465 9694 10107 9696
rect 7465 9691 7531 9694
rect 10041 9691 10107 9694
rect 16481 9754 16547 9757
rect 18413 9754 18479 9757
rect 16481 9752 18479 9754
rect 16481 9696 16486 9752
rect 16542 9696 18418 9752
rect 18474 9696 18479 9752
rect 16481 9694 18479 9696
rect 16481 9691 16547 9694
rect 18413 9691 18479 9694
rect 19241 9754 19307 9757
rect 25589 9754 25655 9757
rect 19241 9752 25655 9754
rect 19241 9696 19246 9752
rect 19302 9696 25594 9752
rect 25650 9696 25655 9752
rect 19241 9694 25655 9696
rect 19241 9691 19307 9694
rect 25589 9691 25655 9694
rect 16389 9618 16455 9621
rect 18505 9618 18571 9621
rect 16389 9616 18571 9618
rect 16389 9560 16394 9616
rect 16450 9560 18510 9616
rect 18566 9560 18571 9616
rect 16389 9558 18571 9560
rect 16389 9555 16455 9558
rect 18505 9555 18571 9558
rect 19149 9620 19215 9621
rect 19149 9616 19196 9620
rect 19260 9618 19266 9620
rect 19149 9560 19154 9616
rect 19149 9556 19196 9560
rect 19260 9558 19306 9618
rect 19260 9556 19266 9558
rect 19149 9555 19215 9556
rect 11145 9482 11211 9485
rect 26509 9482 26575 9485
rect 11145 9480 26575 9482
rect 11145 9424 11150 9480
rect 11206 9424 26514 9480
rect 26570 9424 26575 9480
rect 11145 9422 26575 9424
rect 11145 9419 11211 9422
rect 26509 9419 26575 9422
rect 0 9346 480 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 480 9286
rect 1577 9283 1643 9286
rect 26601 9346 26667 9349
rect 29520 9346 30000 9376
rect 26601 9344 30000 9346
rect 26601 9288 26606 9344
rect 26662 9288 30000 9344
rect 26601 9286 30000 9288
rect 26601 9283 26667 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 16205 9210 16271 9213
rect 18045 9210 18111 9213
rect 16205 9208 18111 9210
rect 16205 9152 16210 9208
rect 16266 9152 18050 9208
rect 18106 9152 18111 9208
rect 16205 9150 18111 9152
rect 16205 9147 16271 9150
rect 18045 9147 18111 9150
rect 13169 9074 13235 9077
rect 13537 9074 13603 9077
rect 26417 9074 26483 9077
rect 13169 9072 26483 9074
rect 13169 9016 13174 9072
rect 13230 9016 13542 9072
rect 13598 9016 26422 9072
rect 26478 9016 26483 9072
rect 13169 9014 26483 9016
rect 13169 9011 13235 9014
rect 13537 9011 13603 9014
rect 26417 9011 26483 9014
rect 3877 8938 3943 8941
rect 4061 8938 4127 8941
rect 26509 8938 26575 8941
rect 3877 8936 26575 8938
rect 3877 8880 3882 8936
rect 3938 8880 4066 8936
rect 4122 8880 26514 8936
rect 26570 8880 26575 8936
rect 3877 8878 26575 8880
rect 3877 8875 3943 8878
rect 4061 8875 4127 8878
rect 26509 8875 26575 8878
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 1577 8666 1643 8669
rect 0 8664 1643 8666
rect 0 8608 1582 8664
rect 1638 8608 1643 8664
rect 0 8606 1643 8608
rect 0 8576 480 8606
rect 1577 8603 1643 8606
rect 7925 8666 7991 8669
rect 9949 8666 10015 8669
rect 7925 8664 10015 8666
rect 7925 8608 7930 8664
rect 7986 8608 9954 8664
rect 10010 8608 10015 8664
rect 7925 8606 10015 8608
rect 7925 8603 7991 8606
rect 9949 8603 10015 8606
rect 19609 8666 19675 8669
rect 25773 8666 25839 8669
rect 19609 8664 25839 8666
rect 19609 8608 19614 8664
rect 19670 8608 25778 8664
rect 25834 8608 25839 8664
rect 19609 8606 25839 8608
rect 19609 8603 19675 8606
rect 25773 8603 25839 8606
rect 26693 8666 26759 8669
rect 29520 8666 30000 8696
rect 26693 8664 30000 8666
rect 26693 8608 26698 8664
rect 26754 8608 30000 8664
rect 26693 8606 30000 8608
rect 26693 8603 26759 8606
rect 29520 8576 30000 8606
rect 2037 8530 2103 8533
rect 18321 8530 18387 8533
rect 2037 8528 18387 8530
rect 2037 8472 2042 8528
rect 2098 8472 18326 8528
rect 18382 8472 18387 8528
rect 2037 8470 18387 8472
rect 2037 8467 2103 8470
rect 18321 8467 18387 8470
rect 19885 8394 19951 8397
rect 26509 8394 26575 8397
rect 19885 8392 26575 8394
rect 19885 8336 19890 8392
rect 19946 8336 26514 8392
rect 26570 8336 26575 8392
rect 19885 8334 26575 8336
rect 19885 8331 19951 8334
rect 26509 8331 26575 8334
rect 27705 8394 27771 8397
rect 27705 8392 28642 8394
rect 27705 8336 27710 8392
rect 27766 8336 28642 8392
rect 27705 8334 28642 8336
rect 27705 8331 27771 8334
rect 1945 8258 2011 8261
rect 4613 8258 4679 8261
rect 1945 8256 4679 8258
rect 1945 8200 1950 8256
rect 2006 8200 4618 8256
rect 4674 8200 4679 8256
rect 1945 8198 4679 8200
rect 1945 8195 2011 8198
rect 4613 8195 4679 8198
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 2681 8122 2747 8125
rect 0 8120 2747 8122
rect 0 8064 2686 8120
rect 2742 8064 2747 8120
rect 0 8062 2747 8064
rect 0 8032 480 8062
rect 2681 8059 2747 8062
rect 3325 8122 3391 8125
rect 9765 8122 9831 8125
rect 3325 8120 9831 8122
rect 3325 8064 3330 8120
rect 3386 8064 9770 8120
rect 9826 8064 9831 8120
rect 3325 8062 9831 8064
rect 28582 8122 28642 8334
rect 29520 8122 30000 8152
rect 28582 8062 30000 8122
rect 3325 8059 3391 8062
rect 9765 8059 9831 8062
rect 29520 8032 30000 8062
rect 10777 7986 10843 7989
rect 18413 7986 18479 7989
rect 25037 7986 25103 7989
rect 10777 7984 25103 7986
rect 10777 7928 10782 7984
rect 10838 7928 18418 7984
rect 18474 7928 25042 7984
rect 25098 7928 25103 7984
rect 10777 7926 25103 7928
rect 10777 7923 10843 7926
rect 18413 7923 18479 7926
rect 25037 7923 25103 7926
rect 2681 7850 2747 7853
rect 9029 7850 9095 7853
rect 12617 7850 12683 7853
rect 2681 7848 7666 7850
rect 2681 7792 2686 7848
rect 2742 7792 7666 7848
rect 2681 7790 7666 7792
rect 2681 7787 2747 7790
rect 7606 7714 7666 7790
rect 9029 7848 12683 7850
rect 9029 7792 9034 7848
rect 9090 7792 12622 7848
rect 12678 7792 12683 7848
rect 9029 7790 12683 7792
rect 9029 7787 9095 7790
rect 12617 7787 12683 7790
rect 14181 7714 14247 7717
rect 7606 7712 14247 7714
rect 7606 7656 14186 7712
rect 14242 7656 14247 7712
rect 7606 7654 14247 7656
rect 14181 7651 14247 7654
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 0 7442 480 7472
rect 2589 7442 2655 7445
rect 0 7440 2655 7442
rect 0 7384 2594 7440
rect 2650 7384 2655 7440
rect 0 7382 2655 7384
rect 0 7352 480 7382
rect 2589 7379 2655 7382
rect 9213 7442 9279 7445
rect 18873 7442 18939 7445
rect 9213 7440 18939 7442
rect 9213 7384 9218 7440
rect 9274 7384 18878 7440
rect 18934 7384 18939 7440
rect 9213 7382 18939 7384
rect 9213 7379 9279 7382
rect 18873 7379 18939 7382
rect 26693 7442 26759 7445
rect 29520 7442 30000 7472
rect 26693 7440 30000 7442
rect 26693 7384 26698 7440
rect 26754 7384 30000 7440
rect 26693 7382 30000 7384
rect 26693 7379 26759 7382
rect 29520 7352 30000 7382
rect 8661 7306 8727 7309
rect 11697 7306 11763 7309
rect 8661 7304 11763 7306
rect 8661 7248 8666 7304
rect 8722 7248 11702 7304
rect 11758 7248 11763 7304
rect 8661 7246 11763 7248
rect 8661 7243 8727 7246
rect 11697 7243 11763 7246
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 3325 7034 3391 7037
rect 10685 7034 10751 7037
rect 12801 7034 12867 7037
rect 3325 7032 10751 7034
rect 3325 6976 3330 7032
rect 3386 6976 10690 7032
rect 10746 6976 10751 7032
rect 3325 6974 10751 6976
rect 3325 6971 3391 6974
rect 10685 6971 10751 6974
rect 11470 7032 12867 7034
rect 11470 6976 12806 7032
rect 12862 6976 12867 7032
rect 11470 6974 12867 6976
rect 0 6898 480 6928
rect 4245 6898 4311 6901
rect 11470 6898 11530 6974
rect 12801 6971 12867 6974
rect 26601 7034 26667 7037
rect 26601 7032 26802 7034
rect 26601 6976 26606 7032
rect 26662 6976 26802 7032
rect 26601 6974 26802 6976
rect 26601 6971 26667 6974
rect 0 6896 4311 6898
rect 0 6840 4250 6896
rect 4306 6840 4311 6896
rect 0 6838 4311 6840
rect 0 6808 480 6838
rect 4245 6835 4311 6838
rect 5766 6838 11530 6898
rect 26742 6898 26802 6974
rect 29520 6898 30000 6928
rect 26742 6838 30000 6898
rect 1669 6626 1735 6629
rect 5766 6626 5826 6838
rect 29520 6808 30000 6838
rect 15745 6762 15811 6765
rect 25865 6762 25931 6765
rect 15745 6760 25931 6762
rect 15745 6704 15750 6760
rect 15806 6704 25870 6760
rect 25926 6704 25931 6760
rect 15745 6702 25931 6704
rect 15745 6699 15811 6702
rect 25865 6699 25931 6702
rect 1669 6624 5826 6626
rect 1669 6568 1674 6624
rect 1730 6568 5826 6624
rect 1669 6566 5826 6568
rect 1669 6563 1735 6566
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 17677 6490 17743 6493
rect 25313 6490 25379 6493
rect 17677 6488 25379 6490
rect 17677 6432 17682 6488
rect 17738 6432 25318 6488
rect 25374 6432 25379 6488
rect 17677 6430 25379 6432
rect 17677 6427 17743 6430
rect 25313 6427 25379 6430
rect 0 6354 480 6384
rect 3785 6354 3851 6357
rect 0 6352 3851 6354
rect 0 6296 3790 6352
rect 3846 6296 3851 6352
rect 0 6294 3851 6296
rect 0 6264 480 6294
rect 3785 6291 3851 6294
rect 4613 6354 4679 6357
rect 10869 6354 10935 6357
rect 4613 6352 10935 6354
rect 4613 6296 4618 6352
rect 4674 6296 10874 6352
rect 10930 6296 10935 6352
rect 4613 6294 10935 6296
rect 4613 6291 4679 6294
rect 10869 6291 10935 6294
rect 16481 6354 16547 6357
rect 19241 6354 19307 6357
rect 16481 6352 19307 6354
rect 16481 6296 16486 6352
rect 16542 6296 19246 6352
rect 19302 6296 19307 6352
rect 16481 6294 19307 6296
rect 16481 6291 16547 6294
rect 19241 6291 19307 6294
rect 26693 6354 26759 6357
rect 29520 6354 30000 6384
rect 26693 6352 30000 6354
rect 26693 6296 26698 6352
rect 26754 6296 30000 6352
rect 26693 6294 30000 6296
rect 26693 6291 26759 6294
rect 29520 6264 30000 6294
rect 2129 6218 2195 6221
rect 7189 6218 7255 6221
rect 2129 6216 7255 6218
rect 2129 6160 2134 6216
rect 2190 6160 7194 6216
rect 7250 6160 7255 6216
rect 2129 6158 7255 6160
rect 2129 6155 2195 6158
rect 7189 6155 7255 6158
rect 9765 6218 9831 6221
rect 26509 6218 26575 6221
rect 9765 6216 26575 6218
rect 9765 6160 9770 6216
rect 9826 6160 26514 6216
rect 26570 6160 26575 6216
rect 9765 6158 26575 6160
rect 9765 6155 9831 6158
rect 26509 6155 26575 6158
rect 3141 6082 3207 6085
rect 9305 6082 9371 6085
rect 3141 6080 9371 6082
rect 3141 6024 3146 6080
rect 3202 6024 9310 6080
rect 9366 6024 9371 6080
rect 3141 6022 9371 6024
rect 3141 6019 3207 6022
rect 9305 6019 9371 6022
rect 11329 6082 11395 6085
rect 17493 6082 17559 6085
rect 11329 6080 17559 6082
rect 11329 6024 11334 6080
rect 11390 6024 17498 6080
rect 17554 6024 17559 6080
rect 11329 6022 17559 6024
rect 11329 6019 11395 6022
rect 17493 6019 17559 6022
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 2037 5946 2103 5949
rect 10133 5946 10199 5949
rect 2037 5944 10199 5946
rect 2037 5888 2042 5944
rect 2098 5888 10138 5944
rect 10194 5888 10199 5944
rect 2037 5886 10199 5888
rect 2037 5883 2103 5886
rect 10133 5883 10199 5886
rect 14273 5946 14339 5949
rect 17861 5946 17927 5949
rect 14273 5944 17927 5946
rect 14273 5888 14278 5944
rect 14334 5888 17866 5944
rect 17922 5888 17927 5944
rect 14273 5886 17927 5888
rect 14273 5883 14339 5886
rect 17861 5883 17927 5886
rect 4981 5810 5047 5813
rect 26509 5810 26575 5813
rect 4981 5808 26575 5810
rect 4981 5752 4986 5808
rect 5042 5752 26514 5808
rect 26570 5752 26575 5808
rect 4981 5750 26575 5752
rect 4981 5747 5047 5750
rect 26509 5747 26575 5750
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 9305 5674 9371 5677
rect 16297 5674 16363 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 5766 5614 6562 5674
rect 4245 5538 4311 5541
rect 5766 5538 5826 5614
rect 4245 5536 5826 5538
rect 4245 5480 4250 5536
rect 4306 5480 5826 5536
rect 4245 5478 5826 5480
rect 6502 5538 6562 5614
rect 9305 5672 16363 5674
rect 9305 5616 9310 5672
rect 9366 5616 16302 5672
rect 16358 5616 16363 5672
rect 9305 5614 16363 5616
rect 9305 5611 9371 5614
rect 16297 5611 16363 5614
rect 26601 5674 26667 5677
rect 29520 5674 30000 5704
rect 26601 5672 30000 5674
rect 26601 5616 26606 5672
rect 26662 5616 30000 5672
rect 26601 5614 30000 5616
rect 26601 5611 26667 5614
rect 29520 5584 30000 5614
rect 15285 5538 15351 5541
rect 6502 5536 15351 5538
rect 6502 5480 15290 5536
rect 15346 5480 15351 5536
rect 6502 5478 15351 5480
rect 4245 5475 4311 5478
rect 15285 5475 15351 5478
rect 16481 5538 16547 5541
rect 18045 5538 18111 5541
rect 16481 5536 18111 5538
rect 16481 5480 16486 5536
rect 16542 5480 18050 5536
rect 18106 5480 18111 5536
rect 16481 5478 18111 5480
rect 16481 5475 16547 5478
rect 18045 5475 18111 5478
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 17309 5402 17375 5405
rect 24393 5402 24459 5405
rect 17309 5400 24459 5402
rect 17309 5344 17314 5400
rect 17370 5344 24398 5400
rect 24454 5344 24459 5400
rect 17309 5342 24459 5344
rect 17309 5339 17375 5342
rect 24393 5339 24459 5342
rect 2497 5266 2563 5269
rect 10225 5266 10291 5269
rect 16757 5266 16823 5269
rect 25773 5266 25839 5269
rect 2497 5264 7666 5266
rect 2497 5208 2502 5264
rect 2558 5208 7666 5264
rect 2497 5206 7666 5208
rect 2497 5203 2563 5206
rect 0 5130 480 5160
rect 2681 5130 2747 5133
rect 0 5128 2747 5130
rect 0 5072 2686 5128
rect 2742 5072 2747 5128
rect 0 5070 2747 5072
rect 7606 5130 7666 5206
rect 10225 5264 25839 5266
rect 10225 5208 10230 5264
rect 10286 5208 16762 5264
rect 16818 5208 25778 5264
rect 25834 5208 25839 5264
rect 10225 5206 25839 5208
rect 10225 5203 10291 5206
rect 16757 5203 16823 5206
rect 25773 5203 25839 5206
rect 17401 5130 17467 5133
rect 7606 5128 17467 5130
rect 7606 5072 17406 5128
rect 17462 5072 17467 5128
rect 7606 5070 17467 5072
rect 0 5040 480 5070
rect 2681 5067 2747 5070
rect 17401 5067 17467 5070
rect 26693 5130 26759 5133
rect 29520 5130 30000 5160
rect 26693 5128 30000 5130
rect 26693 5072 26698 5128
rect 26754 5072 30000 5128
rect 26693 5070 30000 5072
rect 26693 5067 26759 5070
rect 29520 5040 30000 5070
rect 2221 4994 2287 4997
rect 10225 4994 10291 4997
rect 2221 4992 10291 4994
rect 2221 4936 2226 4992
rect 2282 4936 10230 4992
rect 10286 4936 10291 4992
rect 2221 4934 10291 4936
rect 2221 4931 2287 4934
rect 10225 4931 10291 4934
rect 11881 4994 11947 4997
rect 17769 4994 17835 4997
rect 11881 4992 17835 4994
rect 11881 4936 11886 4992
rect 11942 4936 17774 4992
rect 17830 4936 17835 4992
rect 11881 4934 17835 4936
rect 11881 4931 11947 4934
rect 17769 4931 17835 4934
rect 24393 4994 24459 4997
rect 26785 4994 26851 4997
rect 24393 4992 26851 4994
rect 24393 4936 24398 4992
rect 24454 4936 26790 4992
rect 26846 4936 26851 4992
rect 24393 4934 26851 4936
rect 24393 4931 24459 4934
rect 26785 4931 26851 4934
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 17309 4858 17375 4861
rect 11470 4856 17375 4858
rect 11470 4800 17314 4856
rect 17370 4800 17375 4856
rect 11470 4798 17375 4800
rect 4337 4722 4403 4725
rect 11470 4722 11530 4798
rect 17309 4795 17375 4798
rect 4337 4720 11530 4722
rect 4337 4664 4342 4720
rect 4398 4664 11530 4720
rect 4337 4662 11530 4664
rect 17125 4722 17191 4725
rect 26509 4722 26575 4725
rect 17125 4720 26575 4722
rect 17125 4664 17130 4720
rect 17186 4664 26514 4720
rect 26570 4664 26575 4720
rect 17125 4662 26575 4664
rect 4337 4659 4403 4662
rect 17125 4659 17191 4662
rect 26509 4659 26575 4662
rect 4429 4586 4495 4589
rect 14365 4586 14431 4589
rect 4429 4584 14431 4586
rect 4429 4528 4434 4584
rect 4490 4528 14370 4584
rect 14426 4528 14431 4584
rect 4429 4526 14431 4528
rect 4429 4523 4495 4526
rect 14365 4523 14431 4526
rect 16849 4586 16915 4589
rect 26417 4586 26483 4589
rect 16849 4584 26483 4586
rect 16849 4528 16854 4584
rect 16910 4528 26422 4584
rect 26478 4528 26483 4584
rect 16849 4526 26483 4528
rect 16849 4523 16915 4526
rect 26417 4523 26483 4526
rect 0 4450 480 4480
rect 1577 4450 1643 4453
rect 0 4448 1643 4450
rect 0 4392 1582 4448
rect 1638 4392 1643 4448
rect 0 4390 1643 4392
rect 0 4360 480 4390
rect 1577 4387 1643 4390
rect 18505 4450 18571 4453
rect 25681 4450 25747 4453
rect 18505 4448 25747 4450
rect 18505 4392 18510 4448
rect 18566 4392 25686 4448
rect 25742 4392 25747 4448
rect 18505 4390 25747 4392
rect 18505 4387 18571 4390
rect 25681 4387 25747 4390
rect 26601 4450 26667 4453
rect 29520 4450 30000 4480
rect 26601 4448 30000 4450
rect 26601 4392 26606 4448
rect 26662 4392 30000 4448
rect 26601 4390 30000 4392
rect 26601 4387 26667 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 13077 4314 13143 4317
rect 15285 4314 15351 4317
rect 13077 4312 15351 4314
rect 13077 4256 13082 4312
rect 13138 4256 15290 4312
rect 15346 4256 15351 4312
rect 13077 4254 15351 4256
rect 13077 4251 13143 4254
rect 15285 4251 15351 4254
rect 18781 4178 18847 4181
rect 24209 4178 24275 4181
rect 18781 4176 24275 4178
rect 18781 4120 18786 4176
rect 18842 4120 24214 4176
rect 24270 4120 24275 4176
rect 18781 4118 24275 4120
rect 18781 4115 18847 4118
rect 24209 4115 24275 4118
rect 8477 4042 8543 4045
rect 12341 4042 12407 4045
rect 8477 4040 12407 4042
rect 8477 3984 8482 4040
rect 8538 3984 12346 4040
rect 12402 3984 12407 4040
rect 8477 3982 12407 3984
rect 8477 3979 8543 3982
rect 12341 3979 12407 3982
rect 19149 4042 19215 4045
rect 25313 4042 25379 4045
rect 19149 4040 25379 4042
rect 19149 3984 19154 4040
rect 19210 3984 25318 4040
rect 25374 3984 25379 4040
rect 19149 3982 25379 3984
rect 19149 3979 19215 3982
rect 25313 3979 25379 3982
rect 0 3906 480 3936
rect 1577 3906 1643 3909
rect 0 3904 1643 3906
rect 0 3848 1582 3904
rect 1638 3848 1643 3904
rect 0 3846 1643 3848
rect 0 3816 480 3846
rect 1577 3843 1643 3846
rect 8569 3906 8635 3909
rect 9765 3906 9831 3909
rect 8569 3904 9831 3906
rect 8569 3848 8574 3904
rect 8630 3848 9770 3904
rect 9826 3848 9831 3904
rect 8569 3846 9831 3848
rect 8569 3843 8635 3846
rect 9765 3843 9831 3846
rect 26693 3906 26759 3909
rect 29520 3906 30000 3936
rect 26693 3904 30000 3906
rect 26693 3848 26698 3904
rect 26754 3848 30000 3904
rect 26693 3846 30000 3848
rect 26693 3843 26759 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 4429 3634 4495 3637
rect 16941 3634 17007 3637
rect 18413 3634 18479 3637
rect 4429 3632 18479 3634
rect 4429 3576 4434 3632
rect 4490 3576 16946 3632
rect 17002 3576 18418 3632
rect 18474 3576 18479 3632
rect 4429 3574 18479 3576
rect 4429 3571 4495 3574
rect 16941 3571 17007 3574
rect 18413 3571 18479 3574
rect 19057 3634 19123 3637
rect 25129 3634 25195 3637
rect 19057 3632 25195 3634
rect 19057 3576 19062 3632
rect 19118 3576 25134 3632
rect 25190 3576 25195 3632
rect 19057 3574 25195 3576
rect 19057 3571 19123 3574
rect 25129 3571 25195 3574
rect 5257 3498 5323 3501
rect 12249 3498 12315 3501
rect 5257 3496 12315 3498
rect 5257 3440 5262 3496
rect 5318 3440 12254 3496
rect 12310 3440 12315 3496
rect 5257 3438 12315 3440
rect 5257 3435 5323 3438
rect 12249 3435 12315 3438
rect 19609 3498 19675 3501
rect 26325 3498 26391 3501
rect 19609 3496 26391 3498
rect 19609 3440 19614 3496
rect 19670 3440 26330 3496
rect 26386 3440 26391 3496
rect 19609 3438 26391 3440
rect 19609 3435 19675 3438
rect 26325 3435 26391 3438
rect 0 3362 480 3392
rect 1577 3362 1643 3365
rect 0 3360 1643 3362
rect 0 3304 1582 3360
rect 1638 3304 1643 3360
rect 0 3302 1643 3304
rect 0 3272 480 3302
rect 1577 3299 1643 3302
rect 26601 3362 26667 3365
rect 29520 3362 30000 3392
rect 26601 3360 30000 3362
rect 26601 3304 26606 3360
rect 26662 3304 30000 3360
rect 26601 3302 30000 3304
rect 26601 3299 26667 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 8569 3090 8635 3093
rect 14273 3090 14339 3093
rect 8569 3088 14339 3090
rect 8569 3032 8574 3088
rect 8630 3032 14278 3088
rect 14334 3032 14339 3088
rect 8569 3030 14339 3032
rect 8569 3027 8635 3030
rect 14273 3027 14339 3030
rect 17493 3090 17559 3093
rect 25497 3090 25563 3093
rect 27337 3090 27403 3093
rect 17493 3088 25330 3090
rect 17493 3032 17498 3088
rect 17554 3032 25330 3088
rect 17493 3030 25330 3032
rect 17493 3027 17559 3030
rect 6269 2954 6335 2957
rect 8477 2954 8543 2957
rect 6269 2952 8543 2954
rect 6269 2896 6274 2952
rect 6330 2896 8482 2952
rect 8538 2896 8543 2952
rect 6269 2894 8543 2896
rect 6269 2891 6335 2894
rect 8477 2891 8543 2894
rect 12065 2954 12131 2957
rect 13813 2954 13879 2957
rect 12065 2952 13879 2954
rect 12065 2896 12070 2952
rect 12126 2896 13818 2952
rect 13874 2896 13879 2952
rect 12065 2894 13879 2896
rect 12065 2891 12131 2894
rect 13813 2891 13879 2894
rect 14365 2954 14431 2957
rect 25037 2954 25103 2957
rect 14365 2952 25103 2954
rect 14365 2896 14370 2952
rect 14426 2896 25042 2952
rect 25098 2896 25103 2952
rect 14365 2894 25103 2896
rect 25270 2954 25330 3030
rect 25497 3088 27403 3090
rect 25497 3032 25502 3088
rect 25558 3032 27342 3088
rect 27398 3032 27403 3088
rect 25497 3030 27403 3032
rect 25497 3027 25563 3030
rect 27337 3027 27403 3030
rect 27521 2954 27587 2957
rect 25270 2952 27587 2954
rect 25270 2896 27526 2952
rect 27582 2896 27587 2952
rect 25270 2894 27587 2896
rect 14365 2891 14431 2894
rect 25037 2891 25103 2894
rect 27521 2891 27587 2894
rect 1485 2818 1551 2821
rect 5533 2818 5599 2821
rect 1485 2816 5599 2818
rect 1485 2760 1490 2816
rect 1546 2760 5538 2816
rect 5594 2760 5599 2816
rect 1485 2758 5599 2760
rect 1485 2755 1551 2758
rect 5533 2755 5599 2758
rect 11605 2818 11671 2821
rect 13905 2818 13971 2821
rect 11605 2816 13971 2818
rect 11605 2760 11610 2816
rect 11666 2760 13910 2816
rect 13966 2760 13971 2816
rect 11605 2758 13971 2760
rect 11605 2755 11671 2758
rect 13905 2755 13971 2758
rect 14457 2818 14523 2821
rect 16941 2818 17007 2821
rect 14457 2816 17007 2818
rect 14457 2760 14462 2816
rect 14518 2760 16946 2816
rect 17002 2760 17007 2816
rect 14457 2758 17007 2760
rect 14457 2755 14523 2758
rect 16941 2755 17007 2758
rect 23013 2818 23079 2821
rect 25221 2818 25287 2821
rect 23013 2816 25287 2818
rect 23013 2760 23018 2816
rect 23074 2760 25226 2816
rect 25282 2760 25287 2816
rect 23013 2758 25287 2760
rect 23013 2755 23079 2758
rect 25221 2755 25287 2758
rect 25497 2818 25563 2821
rect 28349 2818 28415 2821
rect 25497 2816 28415 2818
rect 25497 2760 25502 2816
rect 25558 2760 28354 2816
rect 28410 2760 28415 2816
rect 25497 2758 28415 2760
rect 25497 2755 25563 2758
rect 28349 2755 28415 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 2681 2682 2747 2685
rect 0 2680 2747 2682
rect 0 2624 2686 2680
rect 2742 2624 2747 2680
rect 0 2622 2747 2624
rect 0 2592 480 2622
rect 2681 2619 2747 2622
rect 15469 2682 15535 2685
rect 19425 2682 19491 2685
rect 15469 2680 19491 2682
rect 15469 2624 15474 2680
rect 15530 2624 19430 2680
rect 19486 2624 19491 2680
rect 15469 2622 19491 2624
rect 15469 2619 15535 2622
rect 19425 2619 19491 2622
rect 27061 2682 27127 2685
rect 29520 2682 30000 2712
rect 27061 2680 30000 2682
rect 27061 2624 27066 2680
rect 27122 2624 30000 2680
rect 27061 2622 30000 2624
rect 27061 2619 27127 2622
rect 29520 2592 30000 2622
rect 14549 2546 14615 2549
rect 22829 2546 22895 2549
rect 14549 2544 22895 2546
rect 14549 2488 14554 2544
rect 14610 2488 22834 2544
rect 22890 2488 22895 2544
rect 14549 2486 22895 2488
rect 14549 2483 14615 2486
rect 22829 2483 22895 2486
rect 19149 2412 19215 2413
rect 19149 2410 19196 2412
rect 19104 2408 19196 2410
rect 19104 2352 19154 2408
rect 19104 2350 19196 2352
rect 19149 2348 19196 2350
rect 19260 2348 19266 2412
rect 20161 2410 20227 2413
rect 24577 2410 24643 2413
rect 20161 2408 24643 2410
rect 20161 2352 20166 2408
rect 20222 2352 24582 2408
rect 24638 2352 24643 2408
rect 20161 2350 24643 2352
rect 19149 2347 19215 2348
rect 20161 2347 20227 2350
rect 24577 2347 24643 2350
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 2957 2138 3023 2141
rect 29520 2138 30000 2168
rect 0 2136 3023 2138
rect 0 2080 2962 2136
rect 3018 2080 3023 2136
rect 0 2078 3023 2080
rect 0 2048 480 2078
rect 2957 2075 3023 2078
rect 27478 2078 30000 2138
rect 25865 2002 25931 2005
rect 27478 2002 27538 2078
rect 29520 2048 30000 2078
rect 25865 2000 27538 2002
rect 25865 1944 25870 2000
rect 25926 1944 27538 2000
rect 25865 1942 27538 1944
rect 25865 1939 25931 1942
rect 24761 1730 24827 1733
rect 29361 1730 29427 1733
rect 24761 1728 29427 1730
rect 24761 1672 24766 1728
rect 24822 1672 29366 1728
rect 29422 1672 29427 1728
rect 24761 1670 29427 1672
rect 24761 1667 24827 1670
rect 29361 1667 29427 1670
rect 4613 1594 4679 1597
rect 6637 1594 6703 1597
rect 4613 1592 6703 1594
rect 4613 1536 4618 1592
rect 4674 1536 6642 1592
rect 6698 1536 6703 1592
rect 4613 1534 6703 1536
rect 4613 1531 4679 1534
rect 6637 1531 6703 1534
rect 0 1458 480 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 480 1398
rect 2773 1395 2839 1398
rect 18505 1458 18571 1461
rect 29520 1458 30000 1488
rect 18505 1456 30000 1458
rect 18505 1400 18510 1456
rect 18566 1400 30000 1456
rect 18505 1398 30000 1400
rect 18505 1395 18571 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 1393 914 1459 917
rect 0 912 1459 914
rect 0 856 1398 912
rect 1454 856 1459 912
rect 0 854 1459 856
rect 0 824 480 854
rect 1393 851 1459 854
rect 27705 914 27771 917
rect 29520 914 30000 944
rect 27705 912 30000 914
rect 27705 856 27710 912
rect 27766 856 30000 912
rect 27705 854 30000 856
rect 27705 851 27771 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 1669 370 1735 373
rect 0 368 1735 370
rect 0 312 1674 368
rect 1730 312 1735 368
rect 0 310 1735 312
rect 0 280 480 310
rect 1669 307 1735 310
rect 18321 370 18387 373
rect 29520 370 30000 400
rect 18321 368 30000 370
rect 18321 312 18326 368
rect 18382 312 30000 368
rect 18321 310 30000 312
rect 18321 307 18387 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 9628 10916 9692 10980
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 8156 10236 8220 10300
rect 9628 10100 9692 10164
rect 8156 9964 8220 10028
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 19196 9616 19260 9620
rect 19196 9560 19210 9616
rect 19210 9560 19260 9616
rect 19196 9556 19260 9560
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 19196 2408 19260 2412
rect 19196 2352 19210 2408
rect 19210 2352 19260 2408
rect 19196 2348 19260 2352
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 9627 10980 9693 10981
rect 9627 10916 9628 10980
rect 9692 10916 9693 10980
rect 9627 10915 9693 10916
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 8155 10300 8221 10301
rect 8155 10236 8156 10300
rect 8220 10236 8221 10300
rect 8155 10235 8221 10236
rect 8158 10029 8218 10235
rect 9630 10165 9690 10915
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 9627 10164 9693 10165
rect 9627 10100 9628 10164
rect 9692 10100 9693 10164
rect 9627 10099 9693 10100
rect 8155 10028 8221 10029
rect 8155 9964 8156 10028
rect 8220 9964 8221 10028
rect 8155 9963 8221 9964
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 19195 9620 19261 9621
rect 19195 9556 19196 9620
rect 19260 9556 19261 9620
rect 19195 9555 19261 9556
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 19198 2413 19258 9555
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 19195 2412 19261 2413
rect 19195 2348 19196 2412
rect 19260 2348 19261 2412
rect 19195 2347 19261 2348
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 2128 21264 2688
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
use sky130_fd_sc_hd__fill_1  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1472 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10
timestamp 1604681595
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_17
timestamp 1604681595
transform 1 0 2668 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14
timestamp 1604681595
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2760 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _16_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_28
timestamp 1604681595
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_24
timestamp 1604681595
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26
timestamp 1604681595
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22
timestamp 1604681595
transform 1 0 3128 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1604681595
transform 1 0 3312 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_38
timestamp 1604681595
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_52
timestamp 1604681595
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1604681595
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5336 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1604681595
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__5.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__5.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8556 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__5.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1604681595
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98
timestamp 1604681595
transform 1 0 10120 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_104
timestamp 1604681595
transform 1 0 10672 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__1.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__1.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__2.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__2.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1604681595
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__2.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_139
timestamp 1604681595
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1604681595
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1604681595
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__4.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__3.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__4.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__4.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__3.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1604681595
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 18124 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1604681595
transform 1 0 17204 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_183
timestamp 1604681595
transform 1 0 17940 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1604681595
transform 1 0 16652 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_189
timestamp 1604681595
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_195
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1604681595
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_207
timestamp 1604681595
transform 1 0 20148 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 19964 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1604681595
transform 1 0 19964 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_217
timestamp 1604681595
transform 1 0 21068 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_229
timestamp 1604681595
transform 1 0 22172 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_230 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_241
timestamp 1604681595
transform 1 0 23276 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_259
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_263
timestamp 1604681595
transform 1 0 25300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_267
timestamp 1604681595
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_279
timestamp 1604681595
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1604681595
transform 1 0 26036 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1604681595
transform 1 0 26404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_283
timestamp 1604681595
transform 1 0 27140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_288
timestamp 1604681595
transform 1 0 27600 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_284
timestamp 1604681595
transform 1 0 27232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1604681595
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 27416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 27508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_291
timestamp 1604681595
transform 1 0 27876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp 1604681595
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1604681595
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1604681595
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_45
timestamp 1604681595
transform 1 0 5244 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_57
timestamp 1604681595
transform 1 0 6348 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_69
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_83
timestamp 1604681595
transform 1 0 8740 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 9752 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1604681595
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_98
timestamp 1604681595
transform 1 0 10120 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__1.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_2_106
timestamp 1604681595
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_127
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_139
timestamp 1604681595
transform 1 0 13892 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__3.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_147
timestamp 1604681595
transform 1 0 14628 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1604681595
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_158
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_170
timestamp 1604681595
transform 1 0 16744 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_182
timestamp 1604681595
transform 1 0 17848 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_194
timestamp 1604681595
transform 1 0 18952 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_267
timestamp 1604681595
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_280
timestamp 1604681595
transform 1 0 26864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 1604681595
transform 1 0 27968 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1604681595
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1604681595
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_19
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 3956 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_40
timestamp 1604681595
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_48
timestamp 1604681595
transform 1 0 5520 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1604681595
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1604681595
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1604681595
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_70
timestamp 1604681595
transform 1 0 7544 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1604681595
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1604681595
transform 1 0 8556 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1604681595
transform 1 0 10764 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_117
timestamp 1604681595
transform 1 0 11868 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1604681595
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_131
timestamp 1604681595
transform 1 0 13156 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_143
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_149
timestamp 1604681595
transform 1 0 14812 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_152
timestamp 1604681595
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_156
timestamp 1604681595
transform 1 0 15456 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_161
timestamp 1604681595
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_165
timestamp 1604681595
transform 1 0 16284 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_177
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604681595
transform 1 0 26404 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604681595
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1604681595
transform 1 0 27324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_279
timestamp 1604681595
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_283
timestamp 1604681595
transform 1 0 27140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_287
timestamp 1604681595
transform 1 0 27508 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2300 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_19
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp 1604681595
transform 1 0 4876 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5888 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp 1604681595
transform 1 0 5612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_71
timestamp 1604681595
transform 1 0 7636 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_83
timestamp 1604681595
transform 1 0 8740 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1604681595
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12328 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_121
timestamp 1604681595
transform 1 0 12236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_131
timestamp 1604681595
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1604681595
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_163
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_168
timestamp 1604681595
transform 1 0 16560 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_182
timestamp 1604681595
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_186
timestamp 1604681595
transform 1 0 18216 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_198
timestamp 1604681595
transform 1 0 19320 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604681595
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1604681595
transform 1 0 26864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_292
timestamp 1604681595
transform 1 0 27968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1604681595
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_19
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 3864 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_23
timestamp 1604681595
transform 1 0 3220 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_26
timestamp 1604681595
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp 1604681595
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_47
timestamp 1604681595
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 13340 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_152
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1604681595
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1604681595
transform 1 0 19964 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_217
timestamp 1604681595
transform 1 0 21068 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_229
timestamp 1604681595
transform 1 0 22172 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_241
timestamp 1604681595
transform 1 0 23276 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1604681595
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1604681595
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1604681595
transform 1 0 26220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_279
timestamp 1604681595
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_283
timestamp 1604681595
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_295
timestamp 1604681595
transform 1 0 28244 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1604681595
transform 1 0 1932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1604681595
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_12
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2024 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1604681595
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1604681595
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1604681595
transform 1 0 4876 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1604681595
transform 1 0 5980 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_47
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_52
timestamp 1604681595
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_56
timestamp 1604681595
transform 1 0 6256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1604681595
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7360 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_65
timestamp 1604681595
transform 1 0 7084 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_70
timestamp 1604681595
transform 1 0 7544 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_76
timestamp 1604681595
transform 1 0 8096 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_79
timestamp 1604681595
transform 1 0 8372 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604681595
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1604681595
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1604681595
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_108
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_116
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_125
timestamp 1604681595
transform 1 0 12604 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_130
timestamp 1604681595
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp 1604681595
transform 1 0 13064 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1604681595
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_136
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14260 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_153
timestamp 1604681595
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1604681595
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_146
timestamp 1604681595
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1604681595
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15916 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15732 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17296 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_168
timestamp 1604681595
transform 1 0 16560 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_185
timestamp 1604681595
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_170
timestamp 1604681595
transform 1 0 16744 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1604681595
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_189
timestamp 1604681595
transform 1 0 18492 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1604681595
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1604681595
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_192
timestamp 1604681595
transform 1 0 18768 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_204
timestamp 1604681595
transform 1 0 19872 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1604681595
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_216
timestamp 1604681595
transform 1 0 20976 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_228
timestamp 1604681595
transform 1 0 22080 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1604681595
transform 1 0 26496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1604681595
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_275
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_278
timestamp 1604681595
transform 1 0 26680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_290
timestamp 1604681595
transform 1 0 27784 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_292
timestamp 1604681595
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1604681595
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_298
timestamp 1604681595
transform 1 0 28520 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1604681595
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5704 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_8_48
timestamp 1604681595
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 8188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_69
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_86
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1604681595
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11132 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_8_106
timestamp 1604681595
transform 1 0 10856 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_160
timestamp 1604681595
transform 1 0 15824 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_163
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17848 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_8_175
timestamp 1604681595
transform 1 0 17204 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp 1604681595
transform 1 0 17756 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1604681595
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604681595
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604681595
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604681595
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_10
timestamp 1604681595
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4232 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_31
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_70
timestamp 1604681595
transform 1 0 7544 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_76
timestamp 1604681595
transform 1 0 8096 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1604681595
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_96
timestamp 1604681595
transform 1 0 9936 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1604681595
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1604681595
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1604681595
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_128
timestamp 1604681595
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_141
timestamp 1604681595
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 1604681595
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _11_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_152
timestamp 1604681595
transform 1 0 15088 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_164
timestamp 1604681595
transform 1 0 16192 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1604681595
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_173
timestamp 1604681595
transform 1 0 17020 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1604681595
transform 1 0 26404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1604681595
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1604681595
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_279
timestamp 1604681595
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1604681595
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_287
timestamp 1604681595
transform 1 0 27508 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_36
timestamp 1604681595
transform 1 0 4416 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_48
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_72
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1604681595
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1604681595
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_101
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11316 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_10_106
timestamp 1604681595
transform 1 0 10856 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_110
timestamp 1604681595
transform 1 0 11224 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_131
timestamp 1604681595
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_135
timestamp 1604681595
transform 1 0 13524 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1604681595
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1604681595
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 1604681595
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_165
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16468 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_10_186
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1604681595
transform 1 0 18952 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_191
timestamp 1604681595
transform 1 0 18676 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1604681595
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1604681595
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604681595
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604681595
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604681595
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2760 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_17
timestamp 1604681595
transform 1 0 2668 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _06_
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1604681595
transform 1 0 3956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_38
timestamp 1604681595
transform 1 0 4600 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_52
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_56
timestamp 1604681595
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1604681595
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1604681595
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8832 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1604681595
transform 1 0 9660 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_105
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_111
timestamp 1604681595
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1604681595
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1604681595
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 13800 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_141
timestamp 1604681595
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_145
timestamp 1604681595
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 14812 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_168
timestamp 1604681595
transform 1 0 16560 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_174
timestamp 1604681595
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_178
timestamp 1604681595
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 17664 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18492 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_198
timestamp 1604681595
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_202
timestamp 1604681595
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_206
timestamp 1604681595
transform 1 0 20056 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_218
timestamp 1604681595
transform 1 0 21160 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_230
timestamp 1604681595
transform 1 0 22264 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_242
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1604681595
transform 1 0 26404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1604681595
transform 1 0 27508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1604681595
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1604681595
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_279
timestamp 1604681595
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_283
timestamp 1604681595
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_291
timestamp 1604681595
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1604681595
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1604681595
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5704 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_69
timestamp 1604681595
transform 1 0 7452 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_86
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11132 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1604681595
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_118
timestamp 1604681595
transform 1 0 11960 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_130
timestamp 1604681595
transform 1 0 13064 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_142
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15732 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 17296 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_168
timestamp 1604681595
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_172
timestamp 1604681595
transform 1 0 16928 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_185
timestamp 1604681595
transform 1 0 18124 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_191
timestamp 1604681595
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_280
timestamp 1604681595
transform 1 0 26864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_292
timestamp 1604681595
transform 1 0 27968 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1604681595
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_7
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_20
timestamp 1604681595
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_16
timestamp 1604681595
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_13
timestamp 1604681595
transform 1 0 2300 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_25
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_31
timestamp 1604681595
transform 1 0 3956 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_38
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1604681595
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_42
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_54
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_58
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_53
timestamp 1604681595
transform 1 0 5980 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_61
timestamp 1604681595
transform 1 0 6716 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_64
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1604681595
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_77
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1604681595
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_91
timestamp 1604681595
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_95
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _07_
timestamp 1604681595
transform 1 0 12144 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_112
timestamp 1604681595
transform 1 0 11408 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_127
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_130
timestamp 1604681595
transform 1 0 13064 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_142
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_159
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1604681595
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_162
timestamp 1604681595
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_172
timestamp 1604681595
transform 1 0 16928 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_174
timestamp 1604681595
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_169
timestamp 1604681595
transform 1 0 16652 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_178
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1604681595
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_178
timestamp 1604681595
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17664 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1604681595
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_197
timestamp 1604681595
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1604681595
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1604681595
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_201
timestamp 1604681595
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_193
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1604681595
transform 1 0 19964 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_217
timestamp 1604681595
transform 1 0 21068 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_229
timestamp 1604681595
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_241
timestamp 1604681595
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1604681595
transform 1 0 26496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_275
timestamp 1604681595
transform 1 0 26404 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_278
timestamp 1604681595
transform 1 0 26680 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_290
timestamp 1604681595
transform 1 0 27784 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_280
timestamp 1604681595
transform 1 0 26864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1604681595
transform 1 0 28520 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_292
timestamp 1604681595
transform 1 0 27968 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1604681595
transform 1 0 28520 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 3220 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1604681595
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1604681595
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1604681595
transform 1 0 5152 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_56
timestamp 1604681595
transform 1 0 6256 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1604681595
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1604681595
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1604681595
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_82
timestamp 1604681595
transform 1 0 8648 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_106
timestamp 1604681595
transform 1 0 10856 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _09_
timestamp 1604681595
transform 1 0 13064 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_133
timestamp 1604681595
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1604681595
transform 1 0 13708 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_149
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_157
timestamp 1604681595
transform 1 0 15548 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1604681595
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_197
timestamp 1604681595
transform 1 0 19228 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_209
timestamp 1604681595
transform 1 0 20332 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_221
timestamp 1604681595
transform 1 0 21436 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_233
timestamp 1604681595
transform 1 0 22540 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_241
timestamp 1604681595
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_275
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_278
timestamp 1604681595
transform 1 0 26680 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_290
timestamp 1604681595
transform 1 0 27784 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_298
timestamp 1604681595
transform 1 0 28520 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6716 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_101
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_113
timestamp 1604681595
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_117
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1604681595
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_125
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12880 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_137
timestamp 1604681595
transform 1 0 13708 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1604681595
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17296 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_168
timestamp 1604681595
transform 1 0 16560 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_185
timestamp 1604681595
transform 1 0 18124 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_189
timestamp 1604681595
transform 1 0 18492 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1604681595
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_280
timestamp 1604681595
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_292
timestamp 1604681595
transform 1 0 27968 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_298
timestamp 1604681595
transform 1 0 28520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2760 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_31
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_35
timestamp 1604681595
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_47
timestamp 1604681595
transform 1 0 5428 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9568 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1604681595
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1604681595
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_117
timestamp 1604681595
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_156
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_164
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1604681595
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_173
timestamp 1604681595
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18400 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_207
timestamp 1604681595
transform 1 0 20148 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_219
timestamp 1604681595
transform 1 0 21252 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_231
timestamp 1604681595
transform 1 0 22356 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1604681595
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1604681595
transform 1 0 26404 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1604681595
transform 1 0 26956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_279
timestamp 1604681595
transform 1 0 26772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_283
timestamp 1604681595
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1604681595
transform 1 0 28244 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_7
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1604681595
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_39
timestamp 1604681595
transform 1 0 4692 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5796 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_50
timestamp 1604681595
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_70
timestamp 1604681595
transform 1 0 7544 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_82
timestamp 1604681595
transform 1 0 8648 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 11684 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_106
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_114
timestamp 1604681595
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_124
timestamp 1604681595
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1604681595
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1604681595
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_18_186
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1604681595
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_288
timestamp 1604681595
transform 1 0 27600 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1604681595
transform 1 0 28336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_7
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 1604681595
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1604681595
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_12
timestamp 1604681595
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2944 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_29
timestamp 1604681595
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_39
timestamp 1604681595
transform 1 0 4692 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_33
timestamp 1604681595
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4508 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4508 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4968 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_46
timestamp 1604681595
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_50
timestamp 1604681595
transform 1 0 5704 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1604681595
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_61
timestamp 1604681595
transform 1 0 6716 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_68
timestamp 1604681595
transform 1 0 7360 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_69
timestamp 1604681595
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_73
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_90
timestamp 1604681595
transform 1 0 9384 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_95
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1604681595
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_112
timestamp 1604681595
transform 1 0 11408 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1604681595
transform 1 0 11316 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1604681595
transform 1 0 10948 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12144 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_136
timestamp 1604681595
transform 1 0 13616 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_135
timestamp 1604681595
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_138
timestamp 1604681595
transform 1 0 13800 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 14904 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1604681595
transform 1 0 16652 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_232
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1604681595
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_288
timestamp 1604681595
transform 1 0 27600 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1604681595
transform 1 0 28060 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 1604681595
transform 1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_7
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_13
timestamp 1604681595
transform 1 0 2300 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_16
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_20
timestamp 1604681595
transform 1 0 2944 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _08_
timestamp 1604681595
transform 1 0 3036 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_24
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_36
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_48
timestamp 1604681595
transform 1 0 5520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604681595
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_100
timestamp 1604681595
transform 1 0 10304 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_131
timestamp 1604681595
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_155
timestamp 1604681595
transform 1 0 15364 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_167
timestamp 1604681595
transform 1 0 16468 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604681595
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1604681595
transform 1 0 26956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1604681595
transform 1 0 28060 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11408 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1604681595
transform 1 0 11316 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1604681595
transform 1 0 12236 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_133
timestamp 1604681595
transform 1 0 13340 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1604681595
transform 1 0 27600 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1604681595
transform 1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1604681595
transform 1 0 26956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1604681595
transform 1 0 28060 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_288
timestamp 1604681595
transform 1 0 27600 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_296
timestamp 1604681595
transform 1 0 28336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1604681595
transform 1 0 26956 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1604681595
transform 1 0 28060 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1604681595
transform 1 0 27600 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1604681595
transform 1 0 26956 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_296
timestamp 1604681595
transform 1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1604681595
transform 1 0 28060 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1604681595
transform 1 0 27600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1604681595
transform 1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1604681595
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1604681595
transform 1 0 26956 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1604681595
transform 1 0 28060 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1604681595
transform 1 0 27600 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1604681595
transform 1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1604681595
transform 1 0 17480 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1604681595
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_190
timestamp 1604681595
transform 1 0 18584 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_198
timestamp 1604681595
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_202
timestamp 1604681595
transform 1 0 19688 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_214
timestamp 1604681595
transform 1 0 20792 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_217
timestamp 1604681595
transform 1 0 21068 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1604681595
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_241
timestamp 1604681595
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1604681595
transform 1 0 26956 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1604681595
transform 1 0 28060 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 17296 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1604681595
transform 1 0 17112 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_180
timestamp 1604681595
transform 1 0 17664 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 19504 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 18400 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_192
timestamp 1604681595
transform 1 0 18768 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_204
timestamp 1604681595
transform 1 0 19872 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_219
timestamp 1604681595
transform 1 0 21252 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_231
timestamp 1604681595
transform 1 0 22356 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_243
timestamp 1604681595
transform 1 0 23460 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_255
timestamp 1604681595
transform 1 0 24564 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_267
timestamp 1604681595
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1604681595
transform 1 0 27600 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_296
timestamp 1604681595
transform 1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 9936 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_84
timestamp 1604681595
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_88
timestamp 1604681595
transform 1 0 9200 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_100
timestamp 1604681595
transform 1 0 10304 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 12512 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_112
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_120
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_128
timestamp 1604681595
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_132
timestamp 1604681595
transform 1 0 13248 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_144
timestamp 1604681595
transform 1 0 14352 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 16284 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_156
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_164
timestamp 1604681595
transform 1 0 16192 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_173
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_196
timestamp 1604681595
transform 1 0 19136 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1604681595
transform 1 0 18768 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1604681595
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 19228 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1604681595
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_200
timestamp 1604681595
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 19688 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1604681595
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1604681595
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_214
timestamp 1604681595
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 20424 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_221
timestamp 1604681595
transform 1 0 21436 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_228
timestamp 1604681595
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 21712 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 21528 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_226
timestamp 1604681595
transform 1 0 21896 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_249
timestamp 1604681595
transform 1 0 24012 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_238
timestamp 1604681595
transform 1 0 23000 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_250
timestamp 1604681595
transform 1 0 24104 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 24196 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1604681595
transform 1 0 24380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1604681595
transform 1 0 25484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_262
timestamp 1604681595
transform 1 0 25208 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_277
timestamp 1604681595
transform 1 0 26588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_289
timestamp 1604681595
transform 1 0 27692 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1604681595
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604681595
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1604681595
transform 1 0 28428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604681595
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604681595
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604681595
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604681595
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604681595
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604681595
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 9770 0 9826 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 9678 23520 9734 24000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 10782 0 10838 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 11242 23520 11298 24000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 478 0 534 480 6 bottom_grid_pin_0_
port 4 nsew default tristate
rlabel metal2 s 5630 0 5686 480 6 bottom_grid_pin_10_
port 5 nsew default tristate
rlabel metal2 s 1490 0 1546 480 6 bottom_grid_pin_2_
port 6 nsew default tristate
rlabel metal2 s 2502 0 2558 480 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal2 s 3514 0 3570 480 6 bottom_grid_pin_6_
port 8 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 bottom_grid_pin_8_
port 9 nsew default tristate
rlabel metal2 s 6642 0 6698 480 6 ccff_head
port 10 nsew default input
rlabel metal2 s 7654 0 7710 480 6 ccff_tail
port 11 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 12 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 13 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 14 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 15 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 16 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 17 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 18 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 19 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 20 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 21 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 22 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 23 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 24 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 25 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 26 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 27 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 28 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 29 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 30 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 31 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 32 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 33 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 34 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 35 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 36 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 37 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 38 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 39 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 40 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 41 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 42 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 49 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 50 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 51 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 52 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 53 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 54 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 55 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 56 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 57 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 58 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 59 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 60 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 61 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 62 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 63 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 64 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 65 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 66 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 67 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 68 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 69 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 70 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 71 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 72 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 73 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 74 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 75 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 76 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 77 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 78 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 79 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 80 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 81 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 82 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 83 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 84 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 85 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 86 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 87 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 88 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 89 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 90 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 91 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
port 92 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
port 93 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
port 94 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
port 95 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
port 96 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
port 97 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[0]
port 98 nsew default input
rlabel metal2 s 19062 0 19118 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[1]
port 99 nsew default input
rlabel metal2 s 20074 0 20130 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[2]
port 100 nsew default input
rlabel metal2 s 21086 0 21142 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[3]
port 101 nsew default input
rlabel metal2 s 22190 0 22246 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[4]
port 102 nsew default input
rlabel metal2 s 23202 0 23258 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[5]
port 103 nsew default input
rlabel metal2 s 24214 0 24270 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
port 104 nsew default tristate
rlabel metal2 s 25226 0 25282 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
port 105 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
port 106 nsew default tristate
rlabel metal2 s 27342 0 27398 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
port 107 nsew default tristate
rlabel metal2 s 28354 0 28410 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
port 108 nsew default tristate
rlabel metal2 s 29366 0 29422 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
port 109 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 prog_clk
port 110 nsew default input
rlabel metal2 s 12714 23520 12770 24000 6 top_width_0_height_0__pin_0_
port 111 nsew default input
rlabel metal2 s 20166 23520 20222 24000 6 top_width_0_height_0__pin_10_
port 112 nsew default input
rlabel metal2 s 29182 23520 29238 24000 6 top_width_0_height_0__pin_11_lower
port 113 nsew default tristate
rlabel metal2 s 8206 23520 8262 24000 6 top_width_0_height_0__pin_11_upper
port 114 nsew default tristate
rlabel metal2 s 21730 23520 21786 24000 6 top_width_0_height_0__pin_1_lower
port 115 nsew default tristate
rlabel metal2 s 754 23520 810 24000 6 top_width_0_height_0__pin_1_upper
port 116 nsew default tristate
rlabel metal2 s 14186 23520 14242 24000 6 top_width_0_height_0__pin_2_
port 117 nsew default input
rlabel metal2 s 23202 23520 23258 24000 6 top_width_0_height_0__pin_3_lower
port 118 nsew default tristate
rlabel metal2 s 2226 23520 2282 24000 6 top_width_0_height_0__pin_3_upper
port 119 nsew default tristate
rlabel metal2 s 15750 23520 15806 24000 6 top_width_0_height_0__pin_4_
port 120 nsew default input
rlabel metal2 s 24674 23520 24730 24000 6 top_width_0_height_0__pin_5_lower
port 121 nsew default tristate
rlabel metal2 s 3698 23520 3754 24000 6 top_width_0_height_0__pin_5_upper
port 122 nsew default tristate
rlabel metal2 s 17222 23520 17278 24000 6 top_width_0_height_0__pin_6_
port 123 nsew default input
rlabel metal2 s 26238 23520 26294 24000 6 top_width_0_height_0__pin_7_lower
port 124 nsew default tristate
rlabel metal2 s 5170 23520 5226 24000 6 top_width_0_height_0__pin_7_upper
port 125 nsew default tristate
rlabel metal2 s 18694 23520 18750 24000 6 top_width_0_height_0__pin_8_
port 126 nsew default input
rlabel metal2 s 27710 23520 27766 24000 6 top_width_0_height_0__pin_9_lower
port 127 nsew default tristate
rlabel metal2 s 6734 23520 6790 24000 6 top_width_0_height_0__pin_9_upper
port 128 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 129 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 130 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
