magic
tech sky130A
magscale 1 2
timestamp 1608133486
<< obsli1 >>
rect 1104 2159 18860 14705
<< obsm1 >>
rect 382 1164 19490 15292
<< metal2 >>
rect 1674 16200 1730 17000
rect 4986 16200 5042 17000
rect 8298 16200 8354 17000
rect 11610 16200 11666 17000
rect 14922 16200 14978 17000
rect 18234 16200 18290 17000
rect 386 0 442 800
rect 1214 0 1270 800
rect 2134 0 2190 800
rect 3054 0 3110 800
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15750 0 15806 800
rect 16670 0 16726 800
rect 17590 0 17646 800
rect 18510 0 18566 800
rect 19430 0 19486 800
<< obsm2 >>
rect 388 16144 1618 16833
rect 1786 16144 4930 16833
rect 5098 16144 8242 16833
rect 8410 16144 11554 16833
rect 11722 16144 14866 16833
rect 15034 16144 18178 16833
rect 18346 16144 19484 16833
rect 388 856 19484 16144
rect 498 167 1158 856
rect 1326 167 2078 856
rect 2246 167 2998 856
rect 3166 167 3918 856
rect 4086 167 4838 856
rect 5006 167 5758 856
rect 5926 167 6678 856
rect 6846 167 7506 856
rect 7674 167 8426 856
rect 8594 167 9346 856
rect 9514 167 10266 856
rect 10434 167 11186 856
rect 11354 167 12106 856
rect 12274 167 13026 856
rect 13194 167 13854 856
rect 14022 167 14774 856
rect 14942 167 15694 856
rect 15862 167 16614 856
rect 16782 167 17534 856
rect 17702 167 18454 856
rect 18622 167 19374 856
<< metal3 >>
rect 0 16736 800 16856
rect 0 16464 800 16584
rect 19200 16736 20000 16856
rect 19200 16464 20000 16584
rect 0 16056 800 16176
rect 0 15784 800 15904
rect 19200 16056 20000 16176
rect 19200 15784 20000 15904
rect 0 15376 800 15496
rect 0 15104 800 15224
rect 19200 15376 20000 15496
rect 19200 15104 20000 15224
rect 0 14696 800 14816
rect 0 14424 800 14544
rect 19200 14696 20000 14816
rect 19200 14424 20000 14544
rect 0 14016 800 14136
rect 0 13744 800 13864
rect 0 13472 800 13592
rect 19200 14016 20000 14136
rect 19200 13744 20000 13864
rect 19200 13472 20000 13592
rect 0 13064 800 13184
rect 0 12792 800 12912
rect 19200 13064 20000 13184
rect 19200 12792 20000 12912
rect 0 12384 800 12504
rect 0 12112 800 12232
rect 19200 12384 20000 12504
rect 19200 12112 20000 12232
rect 0 11704 800 11824
rect 0 11432 800 11552
rect 19200 11704 20000 11824
rect 19200 11432 20000 11552
rect 0 11024 800 11144
rect 0 10752 800 10872
rect 19200 11024 20000 11144
rect 19200 10752 20000 10872
rect 0 10344 800 10464
rect 0 10072 800 10192
rect 0 9800 800 9920
rect 19200 10344 20000 10464
rect 19200 10072 20000 10192
rect 19200 9800 20000 9920
rect 0 9392 800 9512
rect 0 9120 800 9240
rect 19200 9392 20000 9512
rect 19200 9120 20000 9240
rect 0 8712 800 8832
rect 0 8440 800 8560
rect 19200 8712 20000 8832
rect 19200 8440 20000 8560
rect 0 8032 800 8152
rect 0 7760 800 7880
rect 19200 8032 20000 8152
rect 19200 7760 20000 7880
rect 0 7352 800 7472
rect 0 7080 800 7200
rect 0 6808 800 6928
rect 19200 7352 20000 7472
rect 19200 7080 20000 7200
rect 19200 6808 20000 6928
rect 0 6400 800 6520
rect 0 6128 800 6248
rect 19200 6400 20000 6520
rect 19200 6128 20000 6248
rect 0 5720 800 5840
rect 0 5448 800 5568
rect 19200 5720 20000 5840
rect 19200 5448 20000 5568
rect 0 5040 800 5160
rect 0 4768 800 4888
rect 19200 5040 20000 5160
rect 19200 4768 20000 4888
rect 0 4360 800 4480
rect 0 4088 800 4208
rect 19200 4360 20000 4480
rect 19200 4088 20000 4208
rect 0 3680 800 3800
rect 0 3408 800 3528
rect 0 3136 800 3256
rect 19200 3680 20000 3800
rect 19200 3408 20000 3528
rect 19200 3136 20000 3256
rect 0 2728 800 2848
rect 0 2456 800 2576
rect 19200 2728 20000 2848
rect 19200 2456 20000 2576
rect 0 2048 800 2168
rect 0 1776 800 1896
rect 19200 2048 20000 2168
rect 19200 1776 20000 1896
rect 0 1368 800 1488
rect 0 1096 800 1216
rect 19200 1368 20000 1488
rect 19200 1096 20000 1216
rect 0 688 800 808
rect 0 416 800 536
rect 0 144 800 264
rect 19200 688 20000 808
rect 19200 416 20000 536
rect 19200 144 20000 264
<< obsm3 >>
rect 880 16384 19120 16829
rect 800 16256 19200 16384
rect 880 15704 19120 16256
rect 800 15576 19200 15704
rect 880 15024 19120 15576
rect 800 14896 19200 15024
rect 880 14344 19120 14896
rect 800 14216 19200 14344
rect 880 13392 19120 14216
rect 800 13264 19200 13392
rect 880 12712 19120 13264
rect 800 12584 19200 12712
rect 880 12032 19120 12584
rect 800 11904 19200 12032
rect 880 11352 19120 11904
rect 800 11224 19200 11352
rect 880 10672 19120 11224
rect 800 10544 19200 10672
rect 880 9720 19120 10544
rect 800 9592 19200 9720
rect 880 9040 19120 9592
rect 800 8912 19200 9040
rect 880 8360 19120 8912
rect 800 8232 19200 8360
rect 880 7680 19120 8232
rect 800 7552 19200 7680
rect 880 6728 19120 7552
rect 800 6600 19200 6728
rect 880 6048 19120 6600
rect 800 5920 19200 6048
rect 880 5368 19120 5920
rect 800 5240 19200 5368
rect 880 4688 19120 5240
rect 800 4560 19200 4688
rect 880 4008 19120 4560
rect 800 3880 19200 4008
rect 880 3056 19120 3880
rect 800 2928 19200 3056
rect 880 2376 19120 2928
rect 800 2248 19200 2376
rect 880 1696 19120 2248
rect 800 1568 19200 1696
rect 880 1016 19120 1568
rect 800 888 19200 1016
rect 880 171 19120 888
<< metal4 >>
rect 3909 2128 4229 14736
rect 6875 2128 7195 14736
<< obsm4 >>
rect 3003 14816 16685 16829
rect 3003 2128 3829 14816
rect 4309 2128 6795 14816
rect 7275 2128 16685 14816
<< labels >>
rlabel metal3 s 0 16736 800 16856 6 REGIN_FEEDTHROUGH
port 1 nsew default input
rlabel metal2 s 18234 16200 18290 17000 6 REGOUT_FEEDTHROUGH
port 2 nsew default output
rlabel metal2 s 16670 0 16726 800 6 SC_IN_BOT
port 3 nsew default input
rlabel metal2 s 1674 16200 1730 17000 6 SC_IN_TOP
port 4 nsew default input
rlabel metal2 s 17590 0 17646 800 6 SC_OUT_BOT
port 5 nsew default output
rlabel metal2 s 4986 16200 5042 17000 6 SC_OUT_TOP
port 6 nsew default output
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_0_
port 7 nsew default output
rlabel metal2 s 11242 0 11298 800 6 bottom_grid_pin_10_
port 8 nsew default output
rlabel metal2 s 12162 0 12218 800 6 bottom_grid_pin_11_
port 9 nsew default output
rlabel metal2 s 13082 0 13138 800 6 bottom_grid_pin_12_
port 10 nsew default output
rlabel metal2 s 13910 0 13966 800 6 bottom_grid_pin_13_
port 11 nsew default output
rlabel metal2 s 14830 0 14886 800 6 bottom_grid_pin_14_
port 12 nsew default output
rlabel metal2 s 15750 0 15806 800 6 bottom_grid_pin_15_
port 13 nsew default output
rlabel metal2 s 3054 0 3110 800 6 bottom_grid_pin_1_
port 14 nsew default output
rlabel metal2 s 3974 0 4030 800 6 bottom_grid_pin_2_
port 15 nsew default output
rlabel metal2 s 4894 0 4950 800 6 bottom_grid_pin_3_
port 16 nsew default output
rlabel metal2 s 5814 0 5870 800 6 bottom_grid_pin_4_
port 17 nsew default output
rlabel metal2 s 6734 0 6790 800 6 bottom_grid_pin_5_
port 18 nsew default output
rlabel metal2 s 7562 0 7618 800 6 bottom_grid_pin_6_
port 19 nsew default output
rlabel metal2 s 8482 0 8538 800 6 bottom_grid_pin_7_
port 20 nsew default output
rlabel metal2 s 9402 0 9458 800 6 bottom_grid_pin_8_
port 21 nsew default output
rlabel metal2 s 10322 0 10378 800 6 bottom_grid_pin_9_
port 22 nsew default output
rlabel metal2 s 386 0 442 800 6 ccff_head
port 23 nsew default input
rlabel metal2 s 1214 0 1270 800 6 ccff_tail
port 24 nsew default output
rlabel metal3 s 0 6808 800 6928 6 chanx_left_in[0]
port 25 nsew default input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[10]
port 26 nsew default input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[11]
port 27 nsew default input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[12]
port 28 nsew default input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[13]
port 29 nsew default input
rlabel metal3 s 0 11432 800 11552 6 chanx_left_in[14]
port 30 nsew default input
rlabel metal3 s 0 11704 800 11824 6 chanx_left_in[15]
port 31 nsew default input
rlabel metal3 s 0 12112 800 12232 6 chanx_left_in[16]
port 32 nsew default input
rlabel metal3 s 0 12384 800 12504 6 chanx_left_in[17]
port 33 nsew default input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[18]
port 34 nsew default input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[19]
port 35 nsew default input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[1]
port 36 nsew default input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[2]
port 37 nsew default input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[3]
port 38 nsew default input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[4]
port 39 nsew default input
rlabel metal3 s 0 8440 800 8560 6 chanx_left_in[5]
port 40 nsew default input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[6]
port 41 nsew default input
rlabel metal3 s 0 9120 800 9240 6 chanx_left_in[7]
port 42 nsew default input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[8]
port 43 nsew default input
rlabel metal3 s 0 9800 800 9920 6 chanx_left_in[9]
port 44 nsew default input
rlabel metal3 s 0 144 800 264 6 chanx_left_out[0]
port 45 nsew default output
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[10]
port 46 nsew default output
rlabel metal3 s 0 3680 800 3800 6 chanx_left_out[11]
port 47 nsew default output
rlabel metal3 s 0 4088 800 4208 6 chanx_left_out[12]
port 48 nsew default output
rlabel metal3 s 0 4360 800 4480 6 chanx_left_out[13]
port 49 nsew default output
rlabel metal3 s 0 4768 800 4888 6 chanx_left_out[14]
port 50 nsew default output
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[15]
port 51 nsew default output
rlabel metal3 s 0 5448 800 5568 6 chanx_left_out[16]
port 52 nsew default output
rlabel metal3 s 0 5720 800 5840 6 chanx_left_out[17]
port 53 nsew default output
rlabel metal3 s 0 6128 800 6248 6 chanx_left_out[18]
port 54 nsew default output
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[19]
port 55 nsew default output
rlabel metal3 s 0 416 800 536 6 chanx_left_out[1]
port 56 nsew default output
rlabel metal3 s 0 688 800 808 6 chanx_left_out[2]
port 57 nsew default output
rlabel metal3 s 0 1096 800 1216 6 chanx_left_out[3]
port 58 nsew default output
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[4]
port 59 nsew default output
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[5]
port 60 nsew default output
rlabel metal3 s 0 2048 800 2168 6 chanx_left_out[6]
port 61 nsew default output
rlabel metal3 s 0 2456 800 2576 6 chanx_left_out[7]
port 62 nsew default output
rlabel metal3 s 0 2728 800 2848 6 chanx_left_out[8]
port 63 nsew default output
rlabel metal3 s 0 3136 800 3256 6 chanx_left_out[9]
port 64 nsew default output
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[0]
port 65 nsew default input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[10]
port 66 nsew default input
rlabel metal3 s 19200 14016 20000 14136 6 chanx_right_in[11]
port 67 nsew default input
rlabel metal3 s 19200 14424 20000 14544 6 chanx_right_in[12]
port 68 nsew default input
rlabel metal3 s 19200 14696 20000 14816 6 chanx_right_in[13]
port 69 nsew default input
rlabel metal3 s 19200 15104 20000 15224 6 chanx_right_in[14]
port 70 nsew default input
rlabel metal3 s 19200 15376 20000 15496 6 chanx_right_in[15]
port 71 nsew default input
rlabel metal3 s 19200 15784 20000 15904 6 chanx_right_in[16]
port 72 nsew default input
rlabel metal3 s 19200 16056 20000 16176 6 chanx_right_in[17]
port 73 nsew default input
rlabel metal3 s 19200 16464 20000 16584 6 chanx_right_in[18]
port 74 nsew default input
rlabel metal3 s 19200 16736 20000 16856 6 chanx_right_in[19]
port 75 nsew default input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[1]
port 76 nsew default input
rlabel metal3 s 19200 11024 20000 11144 6 chanx_right_in[2]
port 77 nsew default input
rlabel metal3 s 19200 11432 20000 11552 6 chanx_right_in[3]
port 78 nsew default input
rlabel metal3 s 19200 11704 20000 11824 6 chanx_right_in[4]
port 79 nsew default input
rlabel metal3 s 19200 12112 20000 12232 6 chanx_right_in[5]
port 80 nsew default input
rlabel metal3 s 19200 12384 20000 12504 6 chanx_right_in[6]
port 81 nsew default input
rlabel metal3 s 19200 12792 20000 12912 6 chanx_right_in[7]
port 82 nsew default input
rlabel metal3 s 19200 13064 20000 13184 6 chanx_right_in[8]
port 83 nsew default input
rlabel metal3 s 19200 13472 20000 13592 6 chanx_right_in[9]
port 84 nsew default input
rlabel metal3 s 19200 3680 20000 3800 6 chanx_right_out[0]
port 85 nsew default output
rlabel metal3 s 19200 7080 20000 7200 6 chanx_right_out[10]
port 86 nsew default output
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[11]
port 87 nsew default output
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[12]
port 88 nsew default output
rlabel metal3 s 19200 8032 20000 8152 6 chanx_right_out[13]
port 89 nsew default output
rlabel metal3 s 19200 8440 20000 8560 6 chanx_right_out[14]
port 90 nsew default output
rlabel metal3 s 19200 8712 20000 8832 6 chanx_right_out[15]
port 91 nsew default output
rlabel metal3 s 19200 9120 20000 9240 6 chanx_right_out[16]
port 92 nsew default output
rlabel metal3 s 19200 9392 20000 9512 6 chanx_right_out[17]
port 93 nsew default output
rlabel metal3 s 19200 9800 20000 9920 6 chanx_right_out[18]
port 94 nsew default output
rlabel metal3 s 19200 10072 20000 10192 6 chanx_right_out[19]
port 95 nsew default output
rlabel metal3 s 19200 4088 20000 4208 6 chanx_right_out[1]
port 96 nsew default output
rlabel metal3 s 19200 4360 20000 4480 6 chanx_right_out[2]
port 97 nsew default output
rlabel metal3 s 19200 4768 20000 4888 6 chanx_right_out[3]
port 98 nsew default output
rlabel metal3 s 19200 5040 20000 5160 6 chanx_right_out[4]
port 99 nsew default output
rlabel metal3 s 19200 5448 20000 5568 6 chanx_right_out[5]
port 100 nsew default output
rlabel metal3 s 19200 5720 20000 5840 6 chanx_right_out[6]
port 101 nsew default output
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[7]
port 102 nsew default output
rlabel metal3 s 19200 6400 20000 6520 6 chanx_right_out[8]
port 103 nsew default output
rlabel metal3 s 19200 6808 20000 6928 6 chanx_right_out[9]
port 104 nsew default output
rlabel metal3 s 19200 3408 20000 3528 6 clk_1_E_in
port 105 nsew default input
rlabel metal2 s 8298 16200 8354 17000 6 clk_1_N_out
port 106 nsew default output
rlabel metal2 s 18510 0 18566 800 6 clk_1_S_out
port 107 nsew default output
rlabel metal3 s 0 16464 800 16584 6 clk_1_W_in
port 108 nsew default input
rlabel metal3 s 19200 3136 20000 3256 6 clk_2_E_in
port 109 nsew default input
rlabel metal3 s 19200 1368 20000 1488 6 clk_2_E_out
port 110 nsew default output
rlabel metal3 s 0 16056 800 16176 6 clk_2_W_in
port 111 nsew default input
rlabel metal3 s 0 14424 800 14544 6 clk_2_W_out
port 112 nsew default output
rlabel metal3 s 19200 2728 20000 2848 6 clk_3_E_in
port 113 nsew default input
rlabel metal3 s 19200 1096 20000 1216 6 clk_3_E_out
port 114 nsew default output
rlabel metal3 s 0 15784 800 15904 6 clk_3_W_in
port 115 nsew default input
rlabel metal3 s 0 14016 800 14136 6 clk_3_W_out
port 116 nsew default output
rlabel metal2 s 11610 16200 11666 17000 6 prog_clk_0_N_in
port 117 nsew default input
rlabel metal2 s 14922 16200 14978 17000 6 prog_clk_0_W_out
port 118 nsew default output
rlabel metal3 s 19200 2456 20000 2576 6 prog_clk_1_E_in
port 119 nsew default input
rlabel metal3 s 19200 688 20000 808 6 prog_clk_1_N_out
port 120 nsew default output
rlabel metal2 s 19430 0 19486 800 6 prog_clk_1_S_out
port 121 nsew default output
rlabel metal3 s 0 15376 800 15496 6 prog_clk_1_W_in
port 122 nsew default input
rlabel metal3 s 19200 2048 20000 2168 6 prog_clk_2_E_in
port 123 nsew default input
rlabel metal3 s 19200 416 20000 536 6 prog_clk_2_E_out
port 124 nsew default output
rlabel metal3 s 0 15104 800 15224 6 prog_clk_2_W_in
port 125 nsew default input
rlabel metal3 s 0 13744 800 13864 6 prog_clk_2_W_out
port 126 nsew default output
rlabel metal3 s 19200 1776 20000 1896 6 prog_clk_3_E_in
port 127 nsew default input
rlabel metal3 s 19200 144 20000 264 6 prog_clk_3_E_out
port 128 nsew default output
rlabel metal3 s 0 14696 800 14816 6 prog_clk_3_W_in
port 129 nsew default input
rlabel metal3 s 0 13472 800 13592 6 prog_clk_3_W_out
port 130 nsew default output
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 131 nsew power input
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 132 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 20000 17000
string LEFview TRUE
<< end >>
