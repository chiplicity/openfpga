VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 2.400 ;
    END
  END Test_en
  PIN bottom_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END bottom_width_0_height_0__pin_16_
  PIN bottom_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.400 ;
    END
  END bottom_width_0_height_0__pin_17_
  PIN bottom_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.400 ;
    END
  END bottom_width_0_height_0__pin_18_
  PIN bottom_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 2.400 ;
    END
  END bottom_width_0_height_0__pin_19_
  PIN bottom_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END bottom_width_0_height_0__pin_20_
  PIN bottom_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 2.400 ;
    END
  END bottom_width_0_height_0__pin_21_
  PIN bottom_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.400 ;
    END
  END bottom_width_0_height_0__pin_22_
  PIN bottom_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 2.400 ;
    END
  END bottom_width_0_height_0__pin_23_
  PIN bottom_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 2.400 ;
    END
  END bottom_width_0_height_0__pin_24_
  PIN bottom_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END bottom_width_0_height_0__pin_25_
  PIN bottom_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 2.400 ;
    END
  END bottom_width_0_height_0__pin_26_
  PIN bottom_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.400 ;
    END
  END bottom_width_0_height_0__pin_27_
  PIN bottom_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.400 ;
    END
  END bottom_width_0_height_0__pin_28_
  PIN bottom_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 2.400 ;
    END
  END bottom_width_0_height_0__pin_29_
  PIN bottom_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 2.400 ;
    END
  END bottom_width_0_height_0__pin_30_
  PIN bottom_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 2.400 ;
    END
  END bottom_width_0_height_0__pin_31_
  PIN bottom_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 2.400 ;
    END
  END bottom_width_0_height_0__pin_42_lower
  PIN bottom_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 2.400 ;
    END
  END bottom_width_0_height_0__pin_42_upper
  PIN bottom_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 2.400 ;
    END
  END bottom_width_0_height_0__pin_43_lower
  PIN bottom_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 2.400 ;
    END
  END bottom_width_0_height_0__pin_43_upper
  PIN bottom_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 2.400 ;
    END
  END bottom_width_0_height_0__pin_44_lower
  PIN bottom_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 2.400 ;
    END
  END bottom_width_0_height_0__pin_44_upper
  PIN bottom_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 2.400 ;
    END
  END bottom_width_0_height_0__pin_45_lower
  PIN bottom_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 2.400 ;
    END
  END bottom_width_0_height_0__pin_45_upper
  PIN bottom_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 2.400 ;
    END
  END bottom_width_0_height_0__pin_46_lower
  PIN bottom_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.400 ;
    END
  END bottom_width_0_height_0__pin_46_upper
  PIN bottom_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 2.400 ;
    END
  END bottom_width_0_height_0__pin_47_lower
  PIN bottom_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 2.400 ;
    END
  END bottom_width_0_height_0__pin_47_upper
  PIN bottom_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 2.400 ;
    END
  END bottom_width_0_height_0__pin_48_lower
  PIN bottom_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.400 ;
    END
  END bottom_width_0_height_0__pin_48_upper
  PIN bottom_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 2.400 ;
    END
  END bottom_width_0_height_0__pin_49_lower
  PIN bottom_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 2.400 ;
    END
  END bottom_width_0_height_0__pin_49_upper
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 2.400 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 2.400 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 51.040 200.000 51.640 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 2.400 ;
    END
  END clk
  PIN left_width_0_height_0__pin_52_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 2.400 167.240 ;
    END
  END left_width_0_height_0__pin_52_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END prog_clk
  PIN right_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 57.160 200.000 57.760 ;
    END
  END right_width_0_height_0__pin_0_
  PIN right_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 117.680 200.000 118.280 ;
    END
  END right_width_0_height_0__pin_10_
  PIN right_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 123.800 200.000 124.400 ;
    END
  END right_width_0_height_0__pin_11_
  PIN right_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 129.920 200.000 130.520 ;
    END
  END right_width_0_height_0__pin_12_
  PIN right_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 136.040 200.000 136.640 ;
    END
  END right_width_0_height_0__pin_13_
  PIN right_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 141.480 200.000 142.080 ;
    END
  END right_width_0_height_0__pin_14_
  PIN right_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 147.600 200.000 148.200 ;
    END
  END right_width_0_height_0__pin_15_
  PIN right_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 63.280 200.000 63.880 ;
    END
  END right_width_0_height_0__pin_1_
  PIN right_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 69.400 200.000 70.000 ;
    END
  END right_width_0_height_0__pin_2_
  PIN right_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 14.320 200.000 14.920 ;
    END
  END right_width_0_height_0__pin_34_lower
  PIN right_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 153.720 200.000 154.320 ;
    END
  END right_width_0_height_0__pin_34_upper
  PIN right_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 20.440 200.000 21.040 ;
    END
  END right_width_0_height_0__pin_35_lower
  PIN right_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 159.840 200.000 160.440 ;
    END
  END right_width_0_height_0__pin_35_upper
  PIN right_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 26.560 200.000 27.160 ;
    END
  END right_width_0_height_0__pin_36_lower
  PIN right_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 165.960 200.000 166.560 ;
    END
  END right_width_0_height_0__pin_36_upper
  PIN right_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 32.680 200.000 33.280 ;
    END
  END right_width_0_height_0__pin_37_lower
  PIN right_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 172.080 200.000 172.680 ;
    END
  END right_width_0_height_0__pin_37_upper
  PIN right_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 38.800 200.000 39.400 ;
    END
  END right_width_0_height_0__pin_38_lower
  PIN right_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 178.200 200.000 178.800 ;
    END
  END right_width_0_height_0__pin_38_upper
  PIN right_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 44.920 200.000 45.520 ;
    END
  END right_width_0_height_0__pin_39_lower
  PIN right_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 184.320 200.000 184.920 ;
    END
  END right_width_0_height_0__pin_39_upper
  PIN right_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 74.840 200.000 75.440 ;
    END
  END right_width_0_height_0__pin_3_
  PIN right_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 2.760 200.000 3.360 ;
    END
  END right_width_0_height_0__pin_40_lower
  PIN right_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 190.440 200.000 191.040 ;
    END
  END right_width_0_height_0__pin_40_upper
  PIN right_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 8.200 200.000 8.800 ;
    END
  END right_width_0_height_0__pin_41_lower
  PIN right_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 196.560 200.000 197.160 ;
    END
  END right_width_0_height_0__pin_41_upper
  PIN right_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 80.960 200.000 81.560 ;
    END
  END right_width_0_height_0__pin_4_
  PIN right_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 87.080 200.000 87.680 ;
    END
  END right_width_0_height_0__pin_5_
  PIN right_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 93.200 200.000 93.800 ;
    END
  END right_width_0_height_0__pin_6_
  PIN right_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 99.320 200.000 99.920 ;
    END
  END right_width_0_height_0__pin_7_
  PIN right_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 105.440 200.000 106.040 ;
    END
  END right_width_0_height_0__pin_8_
  PIN right_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 111.560 200.000 112.160 ;
    END
  END right_width_0_height_0__pin_9_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 197.600 50.050 200.000 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.590 197.600 149.870 200.000 ;
    END
  END top_width_0_height_0__pin_33_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 2.830 2.760 194.120 187.920 ;
      LAYER met2 ;
        RECT 2.860 197.320 49.490 197.600 ;
        RECT 50.330 197.320 149.310 197.600 ;
        RECT 150.150 197.320 197.250 197.600 ;
        RECT 2.860 2.680 197.250 197.320 ;
        RECT 3.410 2.400 8.090 2.680 ;
        RECT 8.930 2.400 13.610 2.680 ;
        RECT 14.450 2.400 19.130 2.680 ;
        RECT 19.970 2.400 24.650 2.680 ;
        RECT 25.490 2.400 30.170 2.680 ;
        RECT 31.010 2.400 35.690 2.680 ;
        RECT 36.530 2.400 41.210 2.680 ;
        RECT 42.050 2.400 46.730 2.680 ;
        RECT 47.570 2.400 52.250 2.680 ;
        RECT 53.090 2.400 57.770 2.680 ;
        RECT 58.610 2.400 63.290 2.680 ;
        RECT 64.130 2.400 69.270 2.680 ;
        RECT 70.110 2.400 74.790 2.680 ;
        RECT 75.630 2.400 80.310 2.680 ;
        RECT 81.150 2.400 85.830 2.680 ;
        RECT 86.670 2.400 91.350 2.680 ;
        RECT 92.190 2.400 96.870 2.680 ;
        RECT 97.710 2.400 102.390 2.680 ;
        RECT 103.230 2.400 107.910 2.680 ;
        RECT 108.750 2.400 113.430 2.680 ;
        RECT 114.270 2.400 118.950 2.680 ;
        RECT 119.790 2.400 124.470 2.680 ;
        RECT 125.310 2.400 129.990 2.680 ;
        RECT 130.830 2.400 135.970 2.680 ;
        RECT 136.810 2.400 141.490 2.680 ;
        RECT 142.330 2.400 147.010 2.680 ;
        RECT 147.850 2.400 152.530 2.680 ;
        RECT 153.370 2.400 158.050 2.680 ;
        RECT 158.890 2.400 163.570 2.680 ;
        RECT 164.410 2.400 169.090 2.680 ;
        RECT 169.930 2.400 174.610 2.680 ;
        RECT 175.450 2.400 180.130 2.680 ;
        RECT 180.970 2.400 185.650 2.680 ;
        RECT 186.490 2.400 191.170 2.680 ;
        RECT 192.010 2.400 196.690 2.680 ;
      LAYER met3 ;
        RECT 2.400 196.160 197.200 197.025 ;
        RECT 2.400 191.440 197.600 196.160 ;
        RECT 2.400 190.040 197.200 191.440 ;
        RECT 2.400 185.320 197.600 190.040 ;
        RECT 2.400 183.920 197.200 185.320 ;
        RECT 2.400 179.200 197.600 183.920 ;
        RECT 2.400 177.800 197.200 179.200 ;
        RECT 2.400 173.080 197.600 177.800 ;
        RECT 2.400 171.680 197.200 173.080 ;
        RECT 2.400 167.640 197.600 171.680 ;
        RECT 2.800 166.960 197.600 167.640 ;
        RECT 2.800 166.240 197.200 166.960 ;
        RECT 2.400 165.560 197.200 166.240 ;
        RECT 2.400 160.840 197.600 165.560 ;
        RECT 2.400 159.440 197.200 160.840 ;
        RECT 2.400 154.720 197.600 159.440 ;
        RECT 2.400 153.320 197.200 154.720 ;
        RECT 2.400 148.600 197.600 153.320 ;
        RECT 2.400 147.200 197.200 148.600 ;
        RECT 2.400 142.480 197.600 147.200 ;
        RECT 2.400 141.080 197.200 142.480 ;
        RECT 2.400 137.040 197.600 141.080 ;
        RECT 2.400 135.640 197.200 137.040 ;
        RECT 2.400 130.920 197.600 135.640 ;
        RECT 2.400 129.520 197.200 130.920 ;
        RECT 2.400 124.800 197.600 129.520 ;
        RECT 2.400 123.400 197.200 124.800 ;
        RECT 2.400 118.680 197.600 123.400 ;
        RECT 2.400 117.280 197.200 118.680 ;
        RECT 2.400 112.560 197.600 117.280 ;
        RECT 2.400 111.160 197.200 112.560 ;
        RECT 2.400 106.440 197.600 111.160 ;
        RECT 2.400 105.040 197.200 106.440 ;
        RECT 2.400 101.000 197.600 105.040 ;
        RECT 2.800 100.320 197.600 101.000 ;
        RECT 2.800 99.600 197.200 100.320 ;
        RECT 2.400 98.920 197.200 99.600 ;
        RECT 2.400 94.200 197.600 98.920 ;
        RECT 2.400 92.800 197.200 94.200 ;
        RECT 2.400 88.080 197.600 92.800 ;
        RECT 2.400 86.680 197.200 88.080 ;
        RECT 2.400 81.960 197.600 86.680 ;
        RECT 2.400 80.560 197.200 81.960 ;
        RECT 2.400 75.840 197.600 80.560 ;
        RECT 2.400 74.440 197.200 75.840 ;
        RECT 2.400 70.400 197.600 74.440 ;
        RECT 2.400 69.000 197.200 70.400 ;
        RECT 2.400 64.280 197.600 69.000 ;
        RECT 2.400 62.880 197.200 64.280 ;
        RECT 2.400 58.160 197.600 62.880 ;
        RECT 2.400 56.760 197.200 58.160 ;
        RECT 2.400 52.040 197.600 56.760 ;
        RECT 2.400 50.640 197.200 52.040 ;
        RECT 2.400 45.920 197.600 50.640 ;
        RECT 2.400 44.520 197.200 45.920 ;
        RECT 2.400 39.800 197.600 44.520 ;
        RECT 2.400 38.400 197.200 39.800 ;
        RECT 2.400 34.360 197.600 38.400 ;
        RECT 2.800 33.680 197.600 34.360 ;
        RECT 2.800 32.960 197.200 33.680 ;
        RECT 2.400 32.280 197.200 32.960 ;
        RECT 2.400 27.560 197.600 32.280 ;
        RECT 2.400 26.160 197.200 27.560 ;
        RECT 2.400 21.440 197.600 26.160 ;
        RECT 2.400 20.040 197.200 21.440 ;
        RECT 2.400 15.320 197.600 20.040 ;
        RECT 2.400 13.920 197.200 15.320 ;
        RECT 2.400 9.200 197.600 13.920 ;
        RECT 2.400 7.800 197.200 9.200 ;
        RECT 2.400 3.760 197.600 7.800 ;
        RECT 2.400 2.895 197.200 3.760 ;
      LAYER met4 ;
        RECT 64.270 10.640 97.440 187.920 ;
        RECT 99.840 10.640 176.240 187.920 ;
      LAYER met5 ;
        RECT 64.060 14.500 145.700 16.100 ;
  END
END grid_clb
END LIBRARY

