VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__3_
  CLASS BLOCK ;
  FOREIGN sb_1__3_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 3.440 140.000 4.040 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 10.240 140.000 10.840 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 137.600 3.590 140.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 137.600 10.490 140.000 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 2.400 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 2.400 16.280 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 17.040 140.000 17.640 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 137.600 17.390 140.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 137.600 24.290 140.000 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 2.400 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 2.400 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 137.600 31.190 140.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 23.840 140.000 24.440 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 31.320 140.000 31.920 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.120 140.000 38.720 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.170 137.600 45.450 140.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.920 140.000 45.520 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.070 137.600 52.350 140.000 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 137.600 59.250 140.000 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 2.400 36.680 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 52.400 140.000 53.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.400 49.600 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.400 56.400 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 137.600 66.150 140.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 59.200 140.000 59.800 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 66.000 140.000 66.600 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 2.400 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 73.480 140.000 74.080 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.230 137.600 73.510 140.000 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 2.400 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.280 140.000 80.880 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 2.400 76.120 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 137.600 80.410 140.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 2.400 82.920 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.030 137.600 87.310 140.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 2.400 96.520 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 87.080 140.000 87.680 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 137.600 94.210 140.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 93.880 140.000 94.480 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 2.400 103.320 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 137.600 101.110 140.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 108.160 140.000 108.760 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 114.960 140.000 115.560 ;
    END
  END chany_bottom_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 2.400 ;
    END
  END left_top_grid_pin_11_
  PIN left_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 137.600 115.370 140.000 ;
    END
  END left_top_grid_pin_13_
  PIN left_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 137.600 122.270 140.000 ;
    END
  END left_top_grid_pin_15_
  PIN left_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 2.400 ;
    END
  END left_top_grid_pin_1_
  PIN left_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 2.400 123.040 ;
    END
  END left_top_grid_pin_3_
  PIN left_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 122.440 140.000 123.040 ;
    END
  END left_top_grid_pin_5_
  PIN left_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 137.600 108.470 140.000 ;
    END
  END left_top_grid_pin_7_
  PIN left_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END left_top_grid_pin_9_
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 137.600 129.170 140.000 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 137.600 136.070 140.000 ;
    END
  END right_top_grid_pin_11_
  PIN right_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.400 ;
    END
  END right_top_grid_pin_13_
  PIN right_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 2.400 ;
    END
  END right_top_grid_pin_15_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 2.400 129.840 ;
    END
  END right_top_grid_pin_1_
  PIN right_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.240 140.000 129.840 ;
    END
  END right_top_grid_pin_3_
  PIN right_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 2.400 ;
    END
  END right_top_grid_pin_5_
  PIN right_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.040 140.000 136.640 ;
    END
  END right_top_grid_pin_7_
  PIN right_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 2.400 136.640 ;
    END
  END right_top_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.070 0.380 138.390 137.660 ;
      LAYER met2 ;
        RECT 0.100 137.320 3.030 137.770 ;
        RECT 3.870 137.320 9.930 137.770 ;
        RECT 10.770 137.320 16.830 137.770 ;
        RECT 17.670 137.320 23.730 137.770 ;
        RECT 24.570 137.320 30.630 137.770 ;
        RECT 31.470 137.320 37.990 137.770 ;
        RECT 38.830 137.320 44.890 137.770 ;
        RECT 45.730 137.320 51.790 137.770 ;
        RECT 52.630 137.320 58.690 137.770 ;
        RECT 59.530 137.320 65.590 137.770 ;
        RECT 66.430 137.320 72.950 137.770 ;
        RECT 73.790 137.320 79.850 137.770 ;
        RECT 80.690 137.320 86.750 137.770 ;
        RECT 87.590 137.320 93.650 137.770 ;
        RECT 94.490 137.320 100.550 137.770 ;
        RECT 101.390 137.320 107.910 137.770 ;
        RECT 108.750 137.320 114.810 137.770 ;
        RECT 115.650 137.320 121.710 137.770 ;
        RECT 122.550 137.320 128.610 137.770 ;
        RECT 129.450 137.320 135.510 137.770 ;
        RECT 136.350 137.320 138.370 137.770 ;
        RECT 0.100 2.680 138.370 137.320 ;
        RECT 0.100 0.270 2.570 2.680 ;
        RECT 3.410 0.270 8.550 2.680 ;
        RECT 9.390 0.270 14.990 2.680 ;
        RECT 15.830 0.270 21.430 2.680 ;
        RECT 22.270 0.270 27.870 2.680 ;
        RECT 28.710 0.270 34.310 2.680 ;
        RECT 35.150 0.270 40.290 2.680 ;
        RECT 41.130 0.270 46.730 2.680 ;
        RECT 47.570 0.270 53.170 2.680 ;
        RECT 54.010 0.270 59.610 2.680 ;
        RECT 60.450 0.270 66.050 2.680 ;
        RECT 66.890 0.270 72.490 2.680 ;
        RECT 73.330 0.270 78.470 2.680 ;
        RECT 79.310 0.270 84.910 2.680 ;
        RECT 85.750 0.270 91.350 2.680 ;
        RECT 92.190 0.270 97.790 2.680 ;
        RECT 98.630 0.270 104.230 2.680 ;
        RECT 105.070 0.270 110.210 2.680 ;
        RECT 111.050 0.270 116.650 2.680 ;
        RECT 117.490 0.270 123.090 2.680 ;
        RECT 123.930 0.270 129.530 2.680 ;
        RECT 130.370 0.270 135.970 2.680 ;
        RECT 136.810 0.270 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 135.640 137.200 136.040 ;
        RECT 0.270 130.240 138.650 135.640 ;
        RECT 2.800 128.840 137.200 130.240 ;
        RECT 0.270 123.440 138.650 128.840 ;
        RECT 2.800 122.040 137.200 123.440 ;
        RECT 0.270 116.640 138.650 122.040 ;
        RECT 2.800 115.960 138.650 116.640 ;
        RECT 2.800 115.240 137.200 115.960 ;
        RECT 0.270 114.560 137.200 115.240 ;
        RECT 0.270 109.840 138.650 114.560 ;
        RECT 2.800 109.160 138.650 109.840 ;
        RECT 2.800 108.440 137.200 109.160 ;
        RECT 0.270 107.760 137.200 108.440 ;
        RECT 0.270 103.720 138.650 107.760 ;
        RECT 2.800 102.360 138.650 103.720 ;
        RECT 2.800 102.320 137.200 102.360 ;
        RECT 0.270 100.960 137.200 102.320 ;
        RECT 0.270 96.920 138.650 100.960 ;
        RECT 2.800 95.520 138.650 96.920 ;
        RECT 0.270 94.880 138.650 95.520 ;
        RECT 0.270 93.480 137.200 94.880 ;
        RECT 0.270 90.120 138.650 93.480 ;
        RECT 2.800 88.720 138.650 90.120 ;
        RECT 0.270 88.080 138.650 88.720 ;
        RECT 0.270 86.680 137.200 88.080 ;
        RECT 0.270 83.320 138.650 86.680 ;
        RECT 2.800 81.920 138.650 83.320 ;
        RECT 0.270 81.280 138.650 81.920 ;
        RECT 0.270 79.880 137.200 81.280 ;
        RECT 0.270 76.520 138.650 79.880 ;
        RECT 2.800 75.120 138.650 76.520 ;
        RECT 0.270 74.480 138.650 75.120 ;
        RECT 0.270 73.080 137.200 74.480 ;
        RECT 0.270 70.400 138.650 73.080 ;
        RECT 2.800 69.000 138.650 70.400 ;
        RECT 0.270 67.000 138.650 69.000 ;
        RECT 0.270 65.600 137.200 67.000 ;
        RECT 0.270 63.600 138.650 65.600 ;
        RECT 2.800 62.200 138.650 63.600 ;
        RECT 0.270 60.200 138.650 62.200 ;
        RECT 0.270 58.800 137.200 60.200 ;
        RECT 0.270 56.800 138.650 58.800 ;
        RECT 2.800 55.400 138.650 56.800 ;
        RECT 0.270 53.400 138.650 55.400 ;
        RECT 0.270 52.000 137.200 53.400 ;
        RECT 0.270 50.000 138.650 52.000 ;
        RECT 2.800 48.600 138.650 50.000 ;
        RECT 0.270 45.920 138.650 48.600 ;
        RECT 0.270 44.520 137.200 45.920 ;
        RECT 0.270 43.200 138.650 44.520 ;
        RECT 2.800 41.800 138.650 43.200 ;
        RECT 0.270 39.120 138.650 41.800 ;
        RECT 0.270 37.720 137.200 39.120 ;
        RECT 0.270 37.080 138.650 37.720 ;
        RECT 2.800 35.680 138.650 37.080 ;
        RECT 0.270 32.320 138.650 35.680 ;
        RECT 0.270 30.920 137.200 32.320 ;
        RECT 0.270 30.280 138.650 30.920 ;
        RECT 2.800 28.880 138.650 30.280 ;
        RECT 0.270 24.840 138.650 28.880 ;
        RECT 0.270 23.480 137.200 24.840 ;
        RECT 2.800 23.440 137.200 23.480 ;
        RECT 2.800 22.080 138.650 23.440 ;
        RECT 0.270 18.040 138.650 22.080 ;
        RECT 0.270 16.680 137.200 18.040 ;
        RECT 2.800 16.640 137.200 16.680 ;
        RECT 2.800 15.280 138.650 16.640 ;
        RECT 0.270 11.240 138.650 15.280 ;
        RECT 0.270 9.880 137.200 11.240 ;
        RECT 2.800 9.840 137.200 9.880 ;
        RECT 2.800 8.480 138.650 9.840 ;
        RECT 0.270 4.440 138.650 8.480 ;
        RECT 0.270 3.760 137.200 4.440 ;
        RECT 2.800 3.040 137.200 3.760 ;
        RECT 2.800 2.360 138.650 3.040 ;
        RECT 0.270 0.855 138.650 2.360 ;
      LAYER met4 ;
        RECT 0.295 128.480 138.625 129.705 ;
        RECT 0.295 10.640 27.655 128.480 ;
        RECT 30.055 10.640 50.985 128.480 ;
        RECT 53.385 10.640 138.625 128.480 ;
      LAYER met5 ;
        RECT 19.900 65.500 118.100 67.100 ;
  END
END sb_1__3_
END LIBRARY

