magic
tech EFS8A
magscale 1 2
timestamp 1604399260
<< locali >>
rect 12449 26095 12483 26265
rect 15577 25755 15611 26265
rect 12173 25347 12207 25449
rect 3341 25143 3375 25313
rect 3893 21947 3927 22185
rect 3709 20927 3743 21097
rect 3249 20791 3283 20893
rect 17233 18615 17267 18853
rect 11989 18071 12023 18377
rect 9321 13855 9355 14025
rect 16313 12767 16347 12937
rect 17693 11543 17727 11645
<< viali >>
rect 12449 26265 12483 26299
rect 12449 26061 12483 26095
rect 15577 26265 15611 26299
rect 15577 25721 15611 25755
rect 1961 25449 1995 25483
rect 2881 25449 2915 25483
rect 4813 25449 4847 25483
rect 7113 25449 7147 25483
rect 7481 25449 7515 25483
rect 10977 25449 11011 25483
rect 12081 25449 12115 25483
rect 12173 25449 12207 25483
rect 12633 25449 12667 25483
rect 14473 25449 14507 25483
rect 18521 25449 18555 25483
rect 20177 25449 20211 25483
rect 22661 25449 22695 25483
rect 23029 25449 23063 25483
rect 23765 25449 23799 25483
rect 24225 25449 24259 25483
rect 11345 25381 11379 25415
rect 15853 25381 15887 25415
rect 21557 25381 21591 25415
rect 1409 25313 1443 25347
rect 2789 25313 2823 25347
rect 3341 25313 3375 25347
rect 4721 25313 4755 25347
rect 6929 25313 6963 25347
rect 8493 25313 8527 25347
rect 9965 25313 9999 25347
rect 12173 25313 12207 25347
rect 12449 25313 12483 25347
rect 13001 25313 13035 25347
rect 14289 25313 14323 25347
rect 17141 25313 17175 25347
rect 18337 25313 18371 25347
rect 19993 25313 20027 25347
rect 20545 25313 20579 25347
rect 21741 25313 21775 25347
rect 22845 25313 22879 25347
rect 24041 25313 24075 25347
rect 25145 25313 25179 25347
rect 2973 25245 3007 25279
rect 1593 25177 1627 25211
rect 4997 25245 5031 25279
rect 8585 25245 8619 25279
rect 8769 25245 8803 25279
rect 9137 25245 9171 25279
rect 11437 25245 11471 25279
rect 11529 25245 11563 25279
rect 13093 25245 13127 25279
rect 13277 25245 13311 25279
rect 15945 25245 15979 25279
rect 16129 25245 16163 25279
rect 6009 25177 6043 25211
rect 10149 25177 10183 25211
rect 15117 25177 15151 25211
rect 17325 25177 17359 25211
rect 21925 25177 21959 25211
rect 2329 25109 2363 25143
rect 2421 25109 2455 25143
rect 3341 25109 3375 25143
rect 3433 25109 3467 25143
rect 3801 25109 3835 25143
rect 4353 25109 4387 25143
rect 5641 25109 5675 25143
rect 6469 25109 6503 25143
rect 7849 25109 7883 25143
rect 8125 25109 8159 25143
rect 10517 25109 10551 25143
rect 15485 25109 15519 25143
rect 16589 25109 16623 25143
rect 18061 25109 18095 25143
rect 22385 25109 22419 25143
rect 25329 25109 25363 25143
rect 18521 24905 18555 24939
rect 18889 24905 18923 24939
rect 2697 24837 2731 24871
rect 5089 24837 5123 24871
rect 5457 24837 5491 24871
rect 10701 24837 10735 24871
rect 11529 24837 11563 24871
rect 16129 24837 16163 24871
rect 25789 24837 25823 24871
rect 2053 24769 2087 24803
rect 2237 24769 2271 24803
rect 7481 24769 7515 24803
rect 11897 24769 11931 24803
rect 13645 24769 13679 24803
rect 14381 24769 14415 24803
rect 15669 24769 15703 24803
rect 20085 24769 20119 24803
rect 20729 24769 20763 24803
rect 21557 24769 21591 24803
rect 22661 24769 22695 24803
rect 23489 24769 23523 24803
rect 24317 24769 24351 24803
rect 1961 24701 1995 24735
rect 3157 24701 3191 24735
rect 3424 24701 3458 24735
rect 5641 24701 5675 24735
rect 7389 24701 7423 24735
rect 8585 24701 8619 24735
rect 11345 24701 11379 24735
rect 12909 24701 12943 24735
rect 13461 24701 13495 24735
rect 14933 24701 14967 24735
rect 16589 24701 16623 24735
rect 17141 24701 17175 24735
rect 18061 24701 18095 24735
rect 19073 24701 19107 24735
rect 24041 24701 24075 24735
rect 25145 24701 25179 24735
rect 25237 24701 25271 24735
rect 6285 24633 6319 24667
rect 8830 24633 8864 24667
rect 12265 24633 12299 24667
rect 15393 24633 15427 24667
rect 20637 24633 20671 24667
rect 21833 24633 21867 24667
rect 22385 24633 22419 24667
rect 24685 24633 24719 24667
rect 1593 24565 1627 24599
rect 3065 24565 3099 24599
rect 4537 24565 4571 24599
rect 5825 24565 5859 24599
rect 6561 24565 6595 24599
rect 6929 24565 6963 24599
rect 7297 24565 7331 24599
rect 8125 24565 8159 24599
rect 9965 24565 9999 24599
rect 11069 24565 11103 24599
rect 13001 24565 13035 24599
rect 13369 24565 13403 24599
rect 14013 24565 14047 24599
rect 15025 24565 15059 24599
rect 15485 24565 15519 24599
rect 16405 24565 16439 24599
rect 16773 24565 16807 24599
rect 17601 24565 17635 24599
rect 18245 24565 18279 24599
rect 19257 24565 19291 24599
rect 19625 24565 19659 24599
rect 20177 24565 20211 24599
rect 20545 24565 20579 24599
rect 22017 24565 22051 24599
rect 22477 24565 22511 24599
rect 23029 24565 23063 24599
rect 23673 24565 23707 24599
rect 24133 24565 24167 24599
rect 25421 24565 25455 24599
rect 1593 24361 1627 24395
rect 1961 24361 1995 24395
rect 2329 24361 2363 24395
rect 2881 24361 2915 24395
rect 3433 24361 3467 24395
rect 3893 24361 3927 24395
rect 4445 24361 4479 24395
rect 8677 24361 8711 24395
rect 10149 24361 10183 24395
rect 10701 24361 10735 24395
rect 11161 24361 11195 24395
rect 11713 24361 11747 24395
rect 17049 24361 17083 24395
rect 17233 24361 17267 24395
rect 18245 24361 18279 24395
rect 19257 24361 19291 24395
rect 20361 24361 20395 24395
rect 23213 24361 23247 24395
rect 23765 24361 23799 24395
rect 25237 24361 25271 24395
rect 25329 24361 25363 24395
rect 9045 24293 9079 24327
rect 11069 24293 11103 24327
rect 12633 24293 12667 24327
rect 20637 24293 20671 24327
rect 22017 24293 22051 24327
rect 1409 24225 1443 24259
rect 2789 24225 2823 24259
rect 4537 24225 4571 24259
rect 5641 24225 5675 24259
rect 5908 24225 5942 24259
rect 8125 24225 8159 24259
rect 12725 24225 12759 24259
rect 14105 24225 14139 24259
rect 16037 24225 16071 24259
rect 17601 24225 17635 24259
rect 19625 24225 19659 24259
rect 21925 24225 21959 24259
rect 23673 24225 23707 24259
rect 3065 24157 3099 24191
rect 4629 24157 4663 24191
rect 5181 24157 5215 24191
rect 9689 24157 9723 24191
rect 11345 24157 11379 24191
rect 12173 24157 12207 24191
rect 12817 24157 12851 24191
rect 16129 24157 16163 24191
rect 16313 24157 16347 24191
rect 17693 24157 17727 24191
rect 17785 24157 17819 24191
rect 19717 24157 19751 24191
rect 19901 24157 19935 24191
rect 21465 24157 21499 24191
rect 22109 24157 22143 24191
rect 23857 24157 23891 24191
rect 24317 24157 24351 24191
rect 25421 24157 25455 24191
rect 7941 24089 7975 24123
rect 14289 24089 14323 24123
rect 15025 24089 15059 24123
rect 15577 24089 15611 24123
rect 19165 24089 19199 24123
rect 22661 24089 22695 24123
rect 2421 24021 2455 24055
rect 4077 24021 4111 24055
rect 5549 24021 5583 24055
rect 7021 24021 7055 24055
rect 7573 24021 7607 24055
rect 8309 24021 8343 24055
rect 9505 24021 9539 24055
rect 12265 24021 12299 24055
rect 13277 24021 13311 24055
rect 14657 24021 14691 24055
rect 15669 24021 15703 24055
rect 21557 24021 21591 24055
rect 23305 24021 23339 24055
rect 24869 24021 24903 24055
rect 1593 23817 1627 23851
rect 3433 23817 3467 23851
rect 5365 23817 5399 23851
rect 9321 23817 9355 23851
rect 9597 23817 9631 23851
rect 12173 23817 12207 23851
rect 12725 23817 12759 23851
rect 14933 23817 14967 23851
rect 18153 23817 18187 23851
rect 19901 23817 19935 23851
rect 25421 23817 25455 23851
rect 25789 23817 25823 23851
rect 1961 23749 1995 23783
rect 6377 23749 6411 23783
rect 16865 23749 16899 23783
rect 20361 23749 20395 23783
rect 24961 23749 24995 23783
rect 3065 23681 3099 23715
rect 3985 23681 4019 23715
rect 8861 23681 8895 23715
rect 9781 23681 9815 23715
rect 15485 23681 15519 23715
rect 18797 23681 18831 23715
rect 24225 23681 24259 23715
rect 1409 23613 1443 23647
rect 2789 23613 2823 23647
rect 3801 23613 3835 23647
rect 6837 23613 6871 23647
rect 8125 23613 8159 23647
rect 8585 23613 8619 23647
rect 13001 23613 13035 23647
rect 17417 23613 17451 23647
rect 18521 23613 18555 23647
rect 19717 23613 19751 23647
rect 20913 23613 20947 23647
rect 21169 23613 21203 23647
rect 25237 23613 25271 23647
rect 26157 23613 26191 23647
rect 2329 23545 2363 23579
rect 4230 23545 4264 23579
rect 10026 23545 10060 23579
rect 13268 23545 13302 23579
rect 15301 23545 15335 23579
rect 15752 23545 15786 23579
rect 17785 23545 17819 23579
rect 18613 23545 18647 23579
rect 24041 23545 24075 23579
rect 2421 23477 2455 23511
rect 2881 23477 2915 23511
rect 5917 23477 5951 23511
rect 7021 23477 7055 23511
rect 7481 23477 7515 23511
rect 8217 23477 8251 23511
rect 8677 23477 8711 23511
rect 11161 23477 11195 23511
rect 11805 23477 11839 23511
rect 14381 23477 14415 23511
rect 19349 23477 19383 23511
rect 20821 23477 20855 23511
rect 22293 23477 22327 23511
rect 23029 23477 23063 23511
rect 23489 23477 23523 23511
rect 23673 23477 23707 23511
rect 24133 23477 24167 23511
rect 3801 23273 3835 23307
rect 4629 23273 4663 23307
rect 7573 23273 7607 23307
rect 8401 23273 8435 23307
rect 8493 23273 8527 23307
rect 9689 23273 9723 23307
rect 10793 23273 10827 23307
rect 11161 23273 11195 23307
rect 12909 23273 12943 23307
rect 18429 23273 18463 23307
rect 21097 23273 21131 23307
rect 23949 23273 23983 23307
rect 24317 23273 24351 23307
rect 24961 23273 24995 23307
rect 3525 23205 3559 23239
rect 7849 23205 7883 23239
rect 9137 23205 9171 23239
rect 16304 23205 16338 23239
rect 17969 23205 18003 23239
rect 18705 23205 18739 23239
rect 24409 23205 24443 23239
rect 2789 23137 2823 23171
rect 2881 23137 2915 23171
rect 4905 23137 4939 23171
rect 5172 23137 5206 23171
rect 6929 23137 6963 23171
rect 10057 23137 10091 23171
rect 11529 23137 11563 23171
rect 11796 23137 11830 23171
rect 14105 23137 14139 23171
rect 19625 23137 19659 23171
rect 21732 23137 21766 23171
rect 1409 23069 1443 23103
rect 3065 23069 3099 23103
rect 8677 23069 8711 23103
rect 9413 23069 9447 23103
rect 10149 23069 10183 23103
rect 10241 23069 10275 23103
rect 15485 23069 15519 23103
rect 16037 23069 16071 23103
rect 19165 23069 19199 23103
rect 19717 23069 19751 23103
rect 19901 23069 19935 23103
rect 21465 23069 21499 23103
rect 24501 23069 24535 23103
rect 8033 23001 8067 23035
rect 13553 23001 13587 23035
rect 14289 23001 14323 23035
rect 17417 23001 17451 23035
rect 20269 23001 20303 23035
rect 1961 22933 1995 22967
rect 2329 22933 2363 22967
rect 2421 22933 2455 22967
rect 4261 22933 4295 22967
rect 6285 22933 6319 22967
rect 13829 22933 13863 22967
rect 14657 22933 14691 22967
rect 15945 22933 15979 22967
rect 19257 22933 19291 22967
rect 20729 22933 20763 22967
rect 22845 22933 22879 22967
rect 23673 22933 23707 22967
rect 25329 22933 25363 22967
rect 2881 22729 2915 22763
rect 4997 22729 5031 22763
rect 5181 22729 5215 22763
rect 7481 22729 7515 22763
rect 7941 22729 7975 22763
rect 9413 22729 9447 22763
rect 11529 22729 11563 22763
rect 13093 22729 13127 22763
rect 15301 22729 15335 22763
rect 16037 22729 16071 22763
rect 17785 22729 17819 22763
rect 18521 22729 18555 22763
rect 20913 22729 20947 22763
rect 25053 22729 25087 22763
rect 25421 22729 25455 22763
rect 4445 22661 4479 22695
rect 10517 22661 10551 22695
rect 13737 22661 13771 22695
rect 21833 22661 21867 22695
rect 2421 22593 2455 22627
rect 3893 22593 3927 22627
rect 5825 22593 5859 22627
rect 8033 22593 8067 22627
rect 9965 22593 9999 22627
rect 10977 22593 11011 22627
rect 11069 22593 11103 22627
rect 13921 22593 13955 22627
rect 16957 22593 16991 22627
rect 22569 22593 22603 22627
rect 24225 22593 24259 22627
rect 24685 22593 24719 22627
rect 2237 22525 2271 22559
rect 3249 22525 3283 22559
rect 5641 22525 5675 22559
rect 6193 22525 6227 22559
rect 6837 22525 6871 22559
rect 11989 22525 12023 22559
rect 12909 22525 12943 22559
rect 18337 22525 18371 22559
rect 19533 22525 19567 22559
rect 21465 22525 21499 22559
rect 22477 22525 22511 22559
rect 24041 22525 24075 22559
rect 25237 22525 25271 22559
rect 2145 22457 2179 22491
rect 3801 22457 3835 22491
rect 8300 22457 8334 22491
rect 10885 22457 10919 22491
rect 13369 22457 13403 22491
rect 14188 22457 14222 22491
rect 19800 22457 19834 22491
rect 24133 22457 24167 22491
rect 25789 22457 25823 22491
rect 1593 22389 1627 22423
rect 1777 22389 1811 22423
rect 3341 22389 3375 22423
rect 3709 22389 3743 22423
rect 5549 22389 5583 22423
rect 6561 22389 6595 22423
rect 7021 22389 7055 22423
rect 10333 22389 10367 22423
rect 12633 22389 12667 22423
rect 16405 22389 16439 22423
rect 16773 22389 16807 22423
rect 16865 22389 16899 22423
rect 17417 22389 17451 22423
rect 18889 22389 18923 22423
rect 19349 22389 19383 22423
rect 22017 22389 22051 22423
rect 22385 22389 22419 22423
rect 23305 22389 23339 22423
rect 23673 22389 23707 22423
rect 1961 22185 1995 22219
rect 3065 22185 3099 22219
rect 3893 22185 3927 22219
rect 5917 22185 5951 22219
rect 8677 22185 8711 22219
rect 9413 22185 9447 22219
rect 10333 22185 10367 22219
rect 10885 22185 10919 22219
rect 16313 22185 16347 22219
rect 21925 22185 21959 22219
rect 22937 22185 22971 22219
rect 2053 22117 2087 22151
rect 2237 21981 2271 22015
rect 3341 21981 3375 22015
rect 4445 22117 4479 22151
rect 10241 22117 10275 22151
rect 11704 22117 11738 22151
rect 14013 22117 14047 22151
rect 17141 22117 17175 22151
rect 20913 22117 20947 22151
rect 5549 22049 5583 22083
rect 6541 22049 6575 22083
rect 11345 22049 11379 22083
rect 14105 22049 14139 22083
rect 15669 22049 15703 22083
rect 17233 22049 17267 22083
rect 18593 22049 18627 22083
rect 20361 22049 20395 22083
rect 22293 22049 22327 22083
rect 23857 22049 23891 22083
rect 24869 22049 24903 22083
rect 25053 22049 25087 22083
rect 25605 22049 25639 22083
rect 4537 21981 4571 22015
rect 4721 21981 4755 22015
rect 6285 21981 6319 22015
rect 9137 21981 9171 22015
rect 10517 21981 10551 22015
rect 11437 21981 11471 22015
rect 17417 21981 17451 22015
rect 18337 21981 18371 22015
rect 20729 21981 20763 22015
rect 22385 21981 22419 22015
rect 22477 21981 22511 22015
rect 23949 21981 23983 22015
rect 24041 21981 24075 22015
rect 24501 21981 24535 22015
rect 3893 21913 3927 21947
rect 5181 21913 5215 21947
rect 9873 21913 9907 21947
rect 14289 21913 14323 21947
rect 15853 21913 15887 21947
rect 16773 21913 16807 21947
rect 17785 21913 17819 21947
rect 19717 21913 19751 21947
rect 23489 21913 23523 21947
rect 1593 21845 1627 21879
rect 2605 21845 2639 21879
rect 3709 21845 3743 21879
rect 4077 21845 4111 21879
rect 7665 21845 7699 21879
rect 8309 21845 8343 21879
rect 12817 21845 12851 21879
rect 13369 21845 13403 21879
rect 14749 21845 14783 21879
rect 15577 21845 15611 21879
rect 16589 21845 16623 21879
rect 18245 21845 18279 21879
rect 21557 21845 21591 21879
rect 23397 21845 23431 21879
rect 25237 21845 25271 21879
rect 2605 21641 2639 21675
rect 4721 21641 4755 21675
rect 5365 21641 5399 21675
rect 5917 21641 5951 21675
rect 10333 21641 10367 21675
rect 10701 21641 10735 21675
rect 11805 21641 11839 21675
rect 12265 21641 12299 21675
rect 14657 21641 14691 21675
rect 16405 21641 16439 21675
rect 17877 21641 17911 21675
rect 22661 21641 22695 21675
rect 25605 21641 25639 21675
rect 13093 21573 13127 21607
rect 23857 21573 23891 21607
rect 2237 21505 2271 21539
rect 7297 21505 7331 21539
rect 7481 21505 7515 21539
rect 7849 21505 7883 21539
rect 8309 21505 8343 21539
rect 9137 21505 9171 21539
rect 9781 21505 9815 21539
rect 11345 21505 11379 21539
rect 13277 21505 13311 21539
rect 15577 21505 15611 21539
rect 17049 21505 17083 21539
rect 22017 21505 22051 21539
rect 24501 21505 24535 21539
rect 3249 21437 3283 21471
rect 3341 21437 3375 21471
rect 6193 21437 6227 21471
rect 9597 21437 9631 21471
rect 11161 21437 11195 21471
rect 12633 21437 12667 21471
rect 13544 21437 13578 21471
rect 16865 21437 16899 21471
rect 18981 21437 19015 21471
rect 21833 21437 21867 21471
rect 23121 21437 23155 21471
rect 24225 21437 24259 21471
rect 25421 21437 25455 21471
rect 25973 21437 26007 21471
rect 2053 21369 2087 21403
rect 3608 21369 3642 21403
rect 6653 21369 6687 21403
rect 11253 21369 11287 21403
rect 15945 21369 15979 21403
rect 19226 21369 19260 21403
rect 21925 21369 21959 21403
rect 24317 21369 24351 21403
rect 1593 21301 1627 21335
rect 1961 21301 1995 21335
rect 6837 21301 6871 21335
rect 7205 21301 7239 21335
rect 8585 21301 8619 21335
rect 9229 21301 9263 21335
rect 9689 21301 9723 21335
rect 10793 21301 10827 21335
rect 16313 21301 16347 21335
rect 16773 21301 16807 21335
rect 17417 21301 17451 21335
rect 18337 21301 18371 21335
rect 18797 21301 18831 21335
rect 20361 21301 20395 21335
rect 20913 21301 20947 21335
rect 21281 21301 21315 21335
rect 21465 21301 21499 21335
rect 23489 21301 23523 21335
rect 25053 21301 25087 21335
rect 1869 21097 1903 21131
rect 2421 21097 2455 21131
rect 3709 21097 3743 21131
rect 3893 21097 3927 21131
rect 6009 21097 6043 21131
rect 6377 21097 6411 21131
rect 7389 21097 7423 21131
rect 9965 21097 9999 21131
rect 10517 21097 10551 21131
rect 11529 21097 11563 21131
rect 12081 21097 12115 21131
rect 13369 21097 13403 21131
rect 13645 21097 13679 21131
rect 15669 21097 15703 21131
rect 16405 21097 16439 21131
rect 18981 21097 19015 21131
rect 19165 21097 19199 21131
rect 22753 21097 22787 21131
rect 23213 21097 23247 21131
rect 2329 21029 2363 21063
rect 2789 21029 2823 21063
rect 2881 20961 2915 20995
rect 8033 21029 8067 21063
rect 10977 21029 11011 21063
rect 11989 21029 12023 21063
rect 14013 21029 14047 21063
rect 16948 21029 16982 21063
rect 18613 21029 18647 21063
rect 22017 21029 22051 21063
rect 22385 21029 22419 21063
rect 4333 20961 4367 20995
rect 7481 20961 7515 20995
rect 10885 20961 10919 20995
rect 12449 20961 12483 20995
rect 14105 20961 14139 20995
rect 15485 20961 15519 20995
rect 16681 20961 16715 20995
rect 19533 20961 19567 20995
rect 20177 20961 20211 20995
rect 21281 20961 21315 20995
rect 22569 20961 22603 20995
rect 24317 20961 24351 20995
rect 24409 20961 24443 20995
rect 1409 20893 1443 20927
rect 3065 20893 3099 20927
rect 3249 20893 3283 20927
rect 3709 20893 3743 20927
rect 4077 20893 4111 20927
rect 7573 20893 7607 20927
rect 8585 20893 8619 20927
rect 11069 20893 11103 20927
rect 12541 20893 12575 20927
rect 12725 20893 12759 20927
rect 14197 20893 14231 20927
rect 19625 20893 19659 20927
rect 19717 20893 19751 20927
rect 20729 20893 20763 20927
rect 21373 20893 21407 20927
rect 21465 20893 21499 20927
rect 24501 20893 24535 20927
rect 6929 20825 6963 20859
rect 9413 20825 9447 20859
rect 3249 20757 3283 20791
rect 3525 20757 3559 20791
rect 5457 20757 5491 20791
rect 7021 20757 7055 20791
rect 8401 20757 8435 20791
rect 9045 20757 9079 20791
rect 10241 20757 10275 20791
rect 14657 20757 14691 20791
rect 15117 20757 15151 20791
rect 16037 20757 16071 20791
rect 18061 20757 18095 20791
rect 20913 20757 20947 20791
rect 23581 20757 23615 20791
rect 23949 20757 23983 20791
rect 24961 20757 24995 20791
rect 1961 20553 1995 20587
rect 2329 20553 2363 20587
rect 2881 20553 2915 20587
rect 4169 20553 4203 20587
rect 4445 20553 4479 20587
rect 6837 20553 6871 20587
rect 9965 20553 9999 20587
rect 10609 20553 10643 20587
rect 14381 20553 14415 20587
rect 14841 20553 14875 20587
rect 15301 20553 15335 20587
rect 17325 20553 17359 20587
rect 17877 20553 17911 20587
rect 18245 20553 18279 20587
rect 19165 20553 19199 20587
rect 22293 20553 22327 20587
rect 22845 20553 22879 20587
rect 25421 20553 25455 20587
rect 5825 20485 5859 20519
rect 6285 20485 6319 20519
rect 3341 20417 3375 20451
rect 3433 20417 3467 20451
rect 4905 20417 4939 20451
rect 5089 20417 5123 20451
rect 7297 20417 7331 20451
rect 7389 20417 7423 20451
rect 15393 20417 15427 20451
rect 19717 20417 19751 20451
rect 20913 20417 20947 20451
rect 24317 20417 24351 20451
rect 24685 20417 24719 20451
rect 1409 20349 1443 20383
rect 2789 20349 2823 20383
rect 8585 20349 8619 20383
rect 11069 20349 11103 20383
rect 12449 20349 12483 20383
rect 12705 20349 12739 20383
rect 15660 20349 15694 20383
rect 18061 20349 18095 20383
rect 18705 20349 18739 20383
rect 19533 20349 19567 20383
rect 24041 20349 24075 20383
rect 25237 20349 25271 20383
rect 25789 20349 25823 20383
rect 3249 20281 3283 20315
rect 8852 20281 8886 20315
rect 12081 20281 12115 20315
rect 20361 20281 20395 20315
rect 21158 20281 21192 20315
rect 23489 20281 23523 20315
rect 1593 20213 1627 20247
rect 4813 20213 4847 20247
rect 5457 20213 5491 20247
rect 6653 20213 6687 20247
rect 7205 20213 7239 20247
rect 7941 20213 7975 20247
rect 8493 20213 8527 20247
rect 10885 20213 10919 20247
rect 11253 20213 11287 20247
rect 11621 20213 11655 20247
rect 13829 20213 13863 20247
rect 16773 20213 16807 20247
rect 18981 20213 19015 20247
rect 19625 20213 19659 20247
rect 20821 20213 20855 20247
rect 23673 20213 23707 20247
rect 24133 20213 24167 20247
rect 25145 20213 25179 20247
rect 1593 20009 1627 20043
rect 2421 20009 2455 20043
rect 2881 20009 2915 20043
rect 4077 20009 4111 20043
rect 4445 20009 4479 20043
rect 7849 20009 7883 20043
rect 8953 20009 8987 20043
rect 11069 20009 11103 20043
rect 12357 20009 12391 20043
rect 13645 20009 13679 20043
rect 14657 20009 14691 20043
rect 16313 20009 16347 20043
rect 17233 20009 17267 20043
rect 18061 20009 18095 20043
rect 19717 20009 19751 20043
rect 21925 20009 21959 20043
rect 24685 20009 24719 20043
rect 25237 20009 25271 20043
rect 6184 19941 6218 19975
rect 8217 19941 8251 19975
rect 11713 19941 11747 19975
rect 13461 19941 13495 19975
rect 16773 19941 16807 19975
rect 1409 19873 1443 19907
rect 2789 19873 2823 19907
rect 5089 19873 5123 19907
rect 5457 19873 5491 19907
rect 5917 19873 5951 19907
rect 8401 19873 8435 19907
rect 9945 19873 9979 19907
rect 12173 19873 12207 19907
rect 14013 19873 14047 19907
rect 15025 19873 15059 19907
rect 15669 19873 15703 19907
rect 17693 19873 17727 19907
rect 18337 19873 18371 19907
rect 18604 19873 18638 19907
rect 21281 19873 21315 19907
rect 22652 19873 22686 19907
rect 24317 19873 24351 19907
rect 2329 19805 2363 19839
rect 2973 19805 3007 19839
rect 4537 19805 4571 19839
rect 4629 19805 4663 19839
rect 9689 19805 9723 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 15761 19805 15795 19839
rect 15945 19805 15979 19839
rect 22385 19805 22419 19839
rect 25329 19805 25363 19839
rect 25513 19805 25547 19839
rect 7297 19737 7331 19771
rect 15301 19737 15335 19771
rect 1869 19669 1903 19703
rect 3709 19669 3743 19703
rect 8585 19669 8619 19703
rect 9413 19669 9447 19703
rect 11989 19669 12023 19703
rect 12725 19669 12759 19703
rect 13185 19669 13219 19703
rect 20729 19669 20763 19703
rect 21189 19669 21223 19703
rect 21465 19669 21499 19703
rect 23765 19669 23799 19703
rect 24869 19669 24903 19703
rect 2789 19465 2823 19499
rect 4629 19465 4663 19499
rect 5181 19465 5215 19499
rect 6193 19465 6227 19499
rect 10425 19465 10459 19499
rect 16497 19465 16531 19499
rect 16865 19465 16899 19499
rect 17785 19465 17819 19499
rect 20821 19465 20855 19499
rect 25973 19465 26007 19499
rect 25605 19397 25639 19431
rect 1961 19329 1995 19363
rect 4261 19329 4295 19363
rect 5733 19329 5767 19363
rect 7481 19329 7515 19363
rect 9413 19329 9447 19363
rect 10977 19329 11011 19363
rect 13553 19329 13587 19363
rect 18061 19329 18095 19363
rect 21005 19329 21039 19363
rect 1777 19261 1811 19295
rect 2513 19261 2547 19295
rect 4077 19261 4111 19295
rect 5549 19261 5583 19295
rect 6653 19261 6687 19295
rect 9321 19261 9355 19295
rect 10241 19261 10275 19295
rect 10793 19261 10827 19295
rect 11805 19261 11839 19295
rect 13369 19261 13403 19295
rect 14381 19261 14415 19295
rect 14565 19261 14599 19295
rect 14832 19261 14866 19295
rect 23673 19261 23707 19295
rect 3525 19193 3559 19227
rect 5641 19193 5675 19227
rect 18306 19193 18340 19227
rect 20545 19193 20579 19227
rect 21250 19193 21284 19227
rect 22937 19193 22971 19227
rect 23397 19193 23431 19227
rect 23940 19193 23974 19227
rect 1409 19125 1443 19159
rect 1869 19125 1903 19159
rect 3617 19125 3651 19159
rect 3985 19125 4019 19159
rect 5089 19125 5123 19159
rect 6837 19125 6871 19159
rect 7205 19125 7239 19159
rect 7297 19125 7331 19159
rect 7849 19125 7883 19159
rect 8493 19125 8527 19159
rect 8861 19125 8895 19159
rect 9229 19125 9263 19159
rect 9965 19125 9999 19159
rect 10885 19125 10919 19159
rect 11437 19125 11471 19159
rect 12265 19125 12299 19159
rect 12817 19125 12851 19159
rect 13001 19125 13035 19159
rect 13461 19125 13495 19159
rect 14013 19125 14047 19159
rect 15945 19125 15979 19159
rect 17417 19125 17451 19159
rect 19441 19125 19475 19159
rect 22385 19125 22419 19159
rect 25053 19125 25087 19159
rect 1409 18921 1443 18955
rect 3709 18921 3743 18955
rect 4445 18921 4479 18955
rect 7389 18921 7423 18955
rect 10885 18921 10919 18955
rect 11253 18921 11287 18955
rect 13829 18921 13863 18955
rect 14197 18921 14231 18955
rect 17509 18921 17543 18955
rect 19073 18921 19107 18955
rect 21833 18921 21867 18955
rect 23857 18921 23891 18955
rect 24869 18921 24903 18955
rect 25145 18921 25179 18955
rect 2789 18853 2823 18887
rect 6929 18853 6963 18887
rect 7297 18853 7331 18887
rect 15025 18853 15059 18887
rect 17233 18853 17267 18887
rect 17969 18853 18003 18887
rect 19533 18853 19567 18887
rect 21741 18853 21775 18887
rect 23213 18853 23247 18887
rect 24501 18853 24535 18887
rect 6193 18785 6227 18819
rect 7757 18785 7791 18819
rect 10241 18785 10275 18819
rect 11704 18785 11738 18819
rect 13461 18785 13495 18819
rect 14749 18785 14783 18819
rect 16313 18785 16347 18819
rect 2881 18717 2915 18751
rect 2973 18717 3007 18751
rect 4537 18717 4571 18751
rect 4629 18717 4663 18751
rect 6285 18717 6319 18751
rect 6469 18717 6503 18751
rect 7849 18717 7883 18751
rect 7941 18717 7975 18751
rect 10333 18717 10367 18751
rect 10517 18717 10551 18751
rect 11437 18717 11471 18751
rect 16405 18717 16439 18751
rect 16589 18717 16623 18751
rect 2329 18649 2363 18683
rect 4077 18649 4111 18683
rect 5181 18649 5215 18683
rect 5733 18649 5767 18683
rect 9505 18649 9539 18683
rect 15945 18649 15979 18683
rect 16957 18649 16991 18683
rect 17877 18785 17911 18819
rect 19441 18785 19475 18819
rect 22201 18785 22235 18819
rect 23765 18785 23799 18819
rect 24961 18785 24995 18819
rect 25513 18785 25547 18819
rect 18061 18717 18095 18751
rect 18521 18717 18555 18751
rect 19625 18717 19659 18751
rect 22293 18717 22327 18751
rect 22385 18717 22419 18751
rect 23949 18717 23983 18751
rect 1961 18581 1995 18615
rect 2421 18581 2455 18615
rect 5825 18581 5859 18615
rect 8493 18581 8527 18615
rect 8953 18581 8987 18615
rect 9873 18581 9907 18615
rect 12817 18581 12851 18615
rect 15485 18581 15519 18615
rect 17233 18581 17267 18615
rect 17325 18581 17359 18615
rect 20085 18581 20119 18615
rect 21373 18581 21407 18615
rect 22845 18581 22879 18615
rect 23397 18581 23431 18615
rect 2973 18377 3007 18411
rect 5089 18377 5123 18411
rect 6653 18377 6687 18411
rect 11805 18377 11839 18411
rect 11989 18377 12023 18411
rect 14197 18377 14231 18411
rect 16589 18377 16623 18411
rect 17601 18377 17635 18411
rect 18429 18377 18463 18411
rect 23489 18377 23523 18411
rect 25421 18377 25455 18411
rect 26249 18377 26283 18411
rect 4537 18309 4571 18343
rect 5549 18309 5583 18343
rect 7849 18309 7883 18343
rect 2053 18241 2087 18275
rect 8493 18241 8527 18275
rect 3157 18173 3191 18207
rect 3413 18173 3447 18207
rect 5641 18173 5675 18207
rect 8309 18173 8343 18207
rect 9413 18173 9447 18207
rect 9680 18173 9714 18207
rect 1869 18105 1903 18139
rect 2605 18105 2639 18139
rect 6285 18105 6319 18139
rect 9229 18105 9263 18139
rect 25053 18309 25087 18343
rect 12909 18241 12943 18275
rect 13093 18241 13127 18275
rect 13461 18241 13495 18275
rect 14289 18241 14323 18275
rect 16957 18241 16991 18275
rect 22661 18241 22695 18275
rect 24133 18241 24167 18275
rect 24225 18241 24259 18275
rect 12817 18173 12851 18207
rect 14556 18173 14590 18207
rect 19533 18173 19567 18207
rect 22385 18173 22419 18207
rect 24041 18173 24075 18207
rect 24685 18173 24719 18207
rect 25237 18173 25271 18207
rect 25789 18173 25823 18207
rect 12173 18105 12207 18139
rect 16221 18105 16255 18139
rect 19778 18105 19812 18139
rect 21557 18105 21591 18139
rect 1501 18037 1535 18071
rect 1961 18037 1995 18071
rect 5825 18037 5859 18071
rect 6837 18037 6871 18071
rect 7389 18037 7423 18071
rect 8217 18037 8251 18071
rect 8861 18037 8895 18071
rect 10793 18037 10827 18071
rect 11529 18037 11563 18071
rect 11989 18037 12023 18071
rect 12449 18037 12483 18071
rect 15669 18037 15703 18071
rect 18521 18037 18555 18071
rect 19073 18037 19107 18071
rect 20913 18037 20947 18071
rect 21833 18037 21867 18071
rect 22017 18037 22051 18071
rect 22477 18037 22511 18071
rect 23029 18037 23063 18071
rect 23673 18037 23707 18071
rect 2881 17833 2915 17867
rect 3801 17833 3835 17867
rect 4721 17833 4755 17867
rect 6745 17833 6779 17867
rect 7113 17833 7147 17867
rect 9505 17833 9539 17867
rect 10793 17833 10827 17867
rect 11345 17833 11379 17867
rect 12817 17833 12851 17867
rect 13829 17833 13863 17867
rect 14657 17833 14691 17867
rect 19165 17833 19199 17867
rect 19901 17833 19935 17867
rect 22293 17833 22327 17867
rect 22845 17833 22879 17867
rect 1768 17765 1802 17799
rect 7757 17765 7791 17799
rect 10057 17765 10091 17799
rect 13369 17765 13403 17799
rect 17224 17765 17258 17799
rect 23765 17765 23799 17799
rect 24777 17765 24811 17799
rect 3433 17697 3467 17731
rect 5080 17697 5114 17731
rect 7665 17697 7699 17731
rect 9045 17697 9079 17731
rect 11704 17697 11738 17731
rect 15117 17697 15151 17731
rect 15761 17697 15795 17731
rect 16957 17697 16991 17731
rect 19717 17697 19751 17731
rect 21180 17697 21214 17731
rect 24961 17697 24995 17731
rect 1501 17629 1535 17663
rect 4813 17629 4847 17663
rect 7941 17629 7975 17663
rect 10149 17629 10183 17663
rect 10333 17629 10367 17663
rect 11437 17629 11471 17663
rect 14197 17629 14231 17663
rect 15853 17629 15887 17663
rect 16037 17629 16071 17663
rect 20913 17629 20947 17663
rect 23857 17629 23891 17663
rect 24041 17629 24075 17663
rect 7297 17561 7331 17595
rect 9689 17561 9723 17595
rect 15393 17561 15427 17595
rect 23305 17561 23339 17595
rect 4353 17493 4387 17527
rect 6193 17493 6227 17527
rect 8309 17493 8343 17527
rect 8677 17493 8711 17527
rect 16497 17493 16531 17527
rect 16865 17493 16899 17527
rect 18337 17493 18371 17527
rect 19533 17493 19567 17527
rect 23397 17493 23431 17527
rect 24409 17493 24443 17527
rect 25145 17493 25179 17527
rect 25605 17493 25639 17527
rect 3433 17289 3467 17323
rect 4077 17289 4111 17323
rect 4721 17289 4755 17323
rect 7021 17289 7055 17323
rect 7849 17289 7883 17323
rect 10057 17289 10091 17323
rect 11805 17289 11839 17323
rect 12173 17289 12207 17323
rect 12633 17289 12667 17323
rect 13645 17289 13679 17323
rect 15761 17289 15795 17323
rect 16405 17289 16439 17323
rect 17417 17289 17451 17323
rect 18521 17289 18555 17323
rect 1869 17221 1903 17255
rect 4353 17221 4387 17255
rect 6653 17221 6687 17255
rect 9413 17221 9447 17255
rect 12909 17221 12943 17255
rect 20913 17221 20947 17255
rect 23397 17221 23431 17255
rect 2053 17153 2087 17187
rect 5365 17153 5399 17187
rect 5549 17153 5583 17187
rect 11437 17153 11471 17187
rect 13737 17153 13771 17187
rect 16957 17153 16991 17187
rect 18705 17153 18739 17187
rect 21833 17153 21867 17187
rect 22477 17153 22511 17187
rect 23673 17153 23707 17187
rect 2320 17085 2354 17119
rect 5273 17085 5307 17119
rect 6837 17085 6871 17119
rect 8033 17085 8067 17119
rect 11161 17085 11195 17119
rect 11253 17085 11287 17119
rect 12449 17085 12483 17119
rect 14004 17085 14038 17119
rect 16313 17085 16347 17119
rect 16773 17085 16807 17119
rect 22293 17085 22327 17119
rect 8300 17017 8334 17051
rect 10701 17017 10735 17051
rect 16865 17017 16899 17051
rect 18950 17017 18984 17051
rect 22385 17017 22419 17051
rect 23121 17017 23155 17051
rect 23940 17017 23974 17051
rect 4905 16949 4939 16983
rect 6009 16949 6043 16983
rect 7481 16949 7515 16983
rect 10793 16949 10827 16983
rect 15117 16949 15151 16983
rect 17877 16949 17911 16983
rect 20085 16949 20119 16983
rect 21373 16949 21407 16983
rect 21925 16949 21959 16983
rect 25053 16949 25087 16983
rect 25697 16949 25731 16983
rect 1593 16745 1627 16779
rect 1961 16745 1995 16779
rect 2237 16745 2271 16779
rect 2421 16745 2455 16779
rect 4261 16745 4295 16779
rect 4997 16745 5031 16779
rect 6837 16745 6871 16779
rect 7481 16745 7515 16779
rect 8033 16745 8067 16779
rect 8401 16745 8435 16779
rect 9137 16745 9171 16779
rect 10977 16745 11011 16779
rect 13369 16745 13403 16779
rect 13829 16745 13863 16779
rect 15301 16745 15335 16779
rect 15945 16745 15979 16779
rect 17785 16745 17819 16779
rect 18705 16745 18739 16779
rect 18889 16745 18923 16779
rect 19257 16745 19291 16779
rect 19349 16745 19383 16779
rect 20729 16745 20763 16779
rect 20913 16745 20947 16779
rect 21925 16745 21959 16779
rect 22293 16745 22327 16779
rect 22937 16745 22971 16779
rect 24409 16745 24443 16779
rect 2789 16677 2823 16711
rect 5365 16677 5399 16711
rect 5702 16677 5736 16711
rect 7757 16677 7791 16711
rect 9413 16677 9447 16711
rect 23296 16677 23330 16711
rect 1409 16609 1443 16643
rect 3433 16609 3467 16643
rect 3893 16609 3927 16643
rect 4077 16609 4111 16643
rect 5457 16609 5491 16643
rect 8493 16609 8527 16643
rect 10241 16609 10275 16643
rect 11693 16609 11727 16643
rect 13921 16609 13955 16643
rect 14381 16609 14415 16643
rect 15117 16609 15151 16643
rect 16313 16609 16347 16643
rect 16672 16609 16706 16643
rect 19901 16609 19935 16643
rect 21281 16609 21315 16643
rect 23029 16609 23063 16643
rect 2881 16541 2915 16575
rect 3065 16541 3099 16575
rect 8677 16541 8711 16575
rect 10333 16541 10367 16575
rect 10517 16541 10551 16575
rect 11437 16541 11471 16575
rect 16405 16541 16439 16575
rect 19533 16541 19567 16575
rect 21373 16541 21407 16575
rect 21557 16541 21591 16575
rect 9873 16473 9907 16507
rect 11253 16405 11287 16439
rect 12817 16405 12851 16439
rect 18429 16405 18463 16439
rect 20361 16405 20395 16439
rect 2421 16201 2455 16235
rect 5181 16201 5215 16235
rect 6193 16201 6227 16235
rect 6561 16201 6595 16235
rect 9321 16201 9355 16235
rect 9781 16201 9815 16235
rect 11805 16201 11839 16235
rect 14013 16201 14047 16235
rect 15485 16201 15519 16235
rect 16405 16201 16439 16235
rect 18061 16201 18095 16235
rect 19441 16201 19475 16235
rect 19993 16201 20027 16235
rect 21557 16201 21591 16235
rect 23121 16201 23155 16235
rect 23397 16201 23431 16235
rect 5089 16133 5123 16167
rect 21097 16133 21131 16167
rect 22753 16133 22787 16167
rect 2605 16065 2639 16099
rect 4721 16065 4755 16099
rect 5733 16065 5767 16099
rect 6837 16065 6871 16099
rect 13001 16065 13035 16099
rect 13461 16065 13495 16099
rect 14565 16065 14599 16099
rect 17049 16065 17083 16099
rect 18613 16065 18647 16099
rect 19901 16065 19935 16099
rect 20545 16065 20579 16099
rect 21373 16065 21407 16099
rect 22109 16065 22143 16099
rect 23673 16065 23707 16099
rect 1409 15997 1443 16031
rect 5641 15997 5675 16031
rect 9873 15997 9907 16031
rect 13829 15997 13863 16031
rect 14381 15997 14415 16031
rect 16773 15997 16807 16031
rect 17509 15997 17543 16031
rect 20361 15997 20395 16031
rect 21925 15997 21959 16031
rect 2872 15929 2906 15963
rect 5549 15929 5583 15963
rect 7082 15929 7116 15963
rect 10140 15929 10174 15963
rect 12265 15929 12299 15963
rect 12817 15929 12851 15963
rect 19165 15929 19199 15963
rect 22017 15929 22051 15963
rect 23918 15929 23952 15963
rect 1593 15861 1627 15895
rect 2053 15861 2087 15895
rect 3985 15861 4019 15895
rect 8217 15861 8251 15895
rect 8861 15861 8895 15895
rect 11253 15861 11287 15895
rect 12449 15861 12483 15895
rect 12909 15861 12943 15895
rect 14473 15861 14507 15895
rect 15945 15861 15979 15895
rect 16313 15861 16347 15895
rect 16865 15861 16899 15895
rect 17785 15861 17819 15895
rect 18429 15861 18463 15895
rect 18521 15861 18555 15895
rect 20453 15861 20487 15895
rect 25053 15861 25087 15895
rect 1869 15657 1903 15691
rect 2973 15657 3007 15691
rect 3341 15657 3375 15691
rect 4353 15657 4387 15691
rect 4721 15657 4755 15691
rect 5549 15657 5583 15691
rect 8125 15657 8159 15691
rect 8769 15657 8803 15691
rect 9505 15657 9539 15691
rect 9873 15657 9907 15691
rect 10241 15657 10275 15691
rect 10885 15657 10919 15691
rect 11345 15657 11379 15691
rect 12817 15657 12851 15691
rect 16405 15657 16439 15691
rect 17877 15657 17911 15691
rect 18521 15657 18555 15691
rect 19349 15657 19383 15691
rect 21373 15657 21407 15691
rect 22937 15657 22971 15691
rect 23489 15657 23523 15691
rect 23857 15657 23891 15691
rect 6184 15589 6218 15623
rect 8493 15589 8527 15623
rect 11704 15589 11738 15623
rect 13737 15589 13771 15623
rect 20729 15589 20763 15623
rect 2237 15521 2271 15555
rect 2329 15521 2363 15555
rect 3709 15521 3743 15555
rect 4813 15521 4847 15555
rect 5917 15521 5951 15555
rect 8585 15521 8619 15555
rect 11437 15521 11471 15555
rect 13921 15521 13955 15555
rect 16764 15521 16798 15555
rect 21813 15521 21847 15555
rect 24409 15521 24443 15555
rect 24501 15521 24535 15555
rect 1777 15453 1811 15487
rect 2421 15453 2455 15487
rect 4905 15453 4939 15487
rect 10333 15453 10367 15487
rect 10517 15453 10551 15487
rect 15301 15453 15335 15487
rect 16497 15453 16531 15487
rect 19441 15453 19475 15487
rect 19533 15453 19567 15487
rect 21557 15453 21591 15487
rect 24685 15453 24719 15487
rect 9137 15385 9171 15419
rect 14105 15385 14139 15419
rect 18889 15385 18923 15419
rect 7297 15317 7331 15351
rect 13369 15317 13403 15351
rect 14381 15317 14415 15351
rect 18981 15317 19015 15351
rect 19993 15317 20027 15351
rect 24041 15317 24075 15351
rect 4997 15113 5031 15147
rect 6193 15113 6227 15147
rect 6561 15113 6595 15147
rect 7021 15113 7055 15147
rect 9965 15113 9999 15147
rect 10333 15113 10367 15147
rect 10793 15113 10827 15147
rect 11805 15113 11839 15147
rect 12725 15113 12759 15147
rect 16957 15113 16991 15147
rect 17785 15113 17819 15147
rect 21005 15113 21039 15147
rect 21925 15113 21959 15147
rect 22293 15113 22327 15147
rect 22661 15113 22695 15147
rect 23489 15113 23523 15147
rect 23857 15113 23891 15147
rect 25605 15113 25639 15147
rect 3617 15045 3651 15079
rect 7573 15045 7607 15079
rect 24869 15045 24903 15079
rect 25237 15045 25271 15079
rect 1961 14977 1995 15011
rect 2513 14977 2547 15011
rect 2605 14977 2639 15011
rect 3157 14977 3191 15011
rect 4169 14977 4203 15011
rect 4721 14977 4755 15011
rect 5825 14977 5859 15011
rect 7757 14977 7791 15011
rect 11253 14977 11287 15011
rect 11437 14977 11471 15011
rect 13277 14977 13311 15011
rect 18613 14977 18647 15011
rect 24317 14977 24351 15011
rect 24409 14977 24443 15011
rect 5549 14909 5583 14943
rect 5641 14909 5675 14943
rect 14657 14909 14691 14943
rect 16589 14909 16623 14943
rect 18521 14909 18555 14943
rect 19625 14909 19659 14943
rect 22477 14909 22511 14943
rect 23029 14909 23063 14943
rect 24225 14909 24259 14943
rect 25421 14909 25455 14943
rect 25973 14909 26007 14943
rect 3985 14841 4019 14875
rect 8002 14841 8036 14875
rect 12265 14841 12299 14875
rect 13185 14841 13219 14875
rect 14473 14841 14507 14875
rect 14902 14841 14936 14875
rect 17509 14841 17543 14875
rect 18429 14841 18463 14875
rect 19073 14841 19107 14875
rect 19892 14841 19926 14875
rect 2053 14773 2087 14807
rect 2421 14773 2455 14807
rect 3525 14773 3559 14807
rect 4077 14773 4111 14807
rect 5181 14773 5215 14807
rect 9137 14773 9171 14807
rect 10609 14773 10643 14807
rect 11161 14773 11195 14807
rect 13093 14773 13127 14807
rect 14013 14773 14047 14807
rect 16037 14773 16071 14807
rect 18061 14773 18095 14807
rect 19441 14773 19475 14807
rect 21557 14773 21591 14807
rect 2421 14569 2455 14603
rect 2881 14569 2915 14603
rect 3709 14569 3743 14603
rect 4721 14569 4755 14603
rect 6285 14569 6319 14603
rect 9505 14569 9539 14603
rect 11713 14569 11747 14603
rect 11989 14569 12023 14603
rect 12357 14569 12391 14603
rect 13185 14569 13219 14603
rect 13645 14569 13679 14603
rect 17601 14569 17635 14603
rect 18245 14569 18279 14603
rect 18705 14569 18739 14603
rect 20729 14569 20763 14603
rect 23857 14569 23891 14603
rect 24869 14569 24903 14603
rect 25605 14569 25639 14603
rect 4353 14501 4387 14535
rect 21158 14501 21192 14535
rect 24225 14501 24259 14535
rect 1409 14433 1443 14467
rect 2789 14433 2823 14467
rect 5273 14433 5307 14467
rect 6725 14433 6759 14467
rect 9956 14433 9990 14467
rect 12173 14433 12207 14467
rect 14013 14433 14047 14467
rect 16221 14433 16255 14467
rect 16488 14433 16522 14467
rect 19073 14433 19107 14467
rect 23397 14433 23431 14467
rect 25421 14433 25455 14467
rect 2973 14365 3007 14399
rect 5365 14365 5399 14399
rect 5457 14365 5491 14399
rect 6469 14365 6503 14399
rect 9689 14365 9723 14399
rect 14105 14365 14139 14399
rect 14197 14365 14231 14399
rect 19165 14365 19199 14399
rect 19257 14365 19291 14399
rect 20913 14365 20947 14399
rect 24317 14365 24351 14399
rect 24409 14365 24443 14399
rect 4905 14297 4939 14331
rect 5917 14297 5951 14331
rect 7849 14297 7883 14331
rect 8401 14297 8435 14331
rect 22293 14297 22327 14331
rect 1593 14229 1627 14263
rect 2145 14229 2179 14263
rect 9137 14229 9171 14263
rect 11069 14229 11103 14263
rect 12725 14229 12759 14263
rect 13461 14229 13495 14263
rect 14657 14229 14691 14263
rect 16037 14229 16071 14263
rect 18613 14229 18647 14263
rect 19717 14229 19751 14263
rect 23029 14229 23063 14263
rect 23765 14229 23799 14263
rect 1593 14025 1627 14059
rect 2421 14025 2455 14059
rect 2697 14025 2731 14059
rect 6469 14025 6503 14059
rect 7481 14025 7515 14059
rect 9045 14025 9079 14059
rect 9321 14025 9355 14059
rect 9413 14025 9447 14059
rect 11529 14025 11563 14059
rect 13001 14025 13035 14059
rect 13369 14025 13403 14059
rect 15853 14025 15887 14059
rect 17877 14025 17911 14059
rect 21281 14025 21315 14059
rect 21465 14025 21499 14059
rect 23489 14025 23523 14059
rect 2053 13957 2087 13991
rect 5181 13957 5215 13991
rect 8033 13957 8067 13991
rect 3433 13889 3467 13923
rect 4169 13889 4203 13923
rect 5825 13889 5859 13923
rect 8677 13889 8711 13923
rect 14841 13957 14875 13991
rect 16957 13957 16991 13991
rect 19993 13957 20027 13991
rect 23029 13957 23063 13991
rect 23673 13957 23707 13991
rect 16497 13889 16531 13923
rect 20913 13889 20947 13923
rect 21925 13889 21959 13923
rect 22017 13889 22051 13923
rect 24225 13889 24259 13923
rect 26157 13889 26191 13923
rect 1409 13821 1443 13855
rect 2513 13821 2547 13855
rect 4721 13821 4755 13855
rect 7849 13821 7883 13855
rect 8493 13821 8527 13855
rect 9321 13821 9355 13855
rect 9597 13821 9631 13855
rect 9864 13821 9898 13855
rect 13461 13821 13495 13855
rect 15393 13821 15427 13855
rect 16405 13821 16439 13855
rect 18613 13821 18647 13855
rect 24133 13821 24167 13855
rect 25053 13821 25087 13855
rect 25237 13821 25271 13855
rect 25789 13821 25823 13855
rect 3157 13753 3191 13787
rect 4077 13753 4111 13787
rect 5549 13753 5583 13787
rect 6837 13753 6871 13787
rect 8401 13753 8435 13787
rect 12173 13753 12207 13787
rect 13706 13753 13740 13787
rect 18429 13753 18463 13787
rect 18858 13753 18892 13787
rect 24041 13753 24075 13787
rect 3617 13685 3651 13719
rect 3985 13685 4019 13719
rect 4997 13685 5031 13719
rect 5641 13685 5675 13719
rect 10977 13685 11011 13719
rect 12449 13685 12483 13719
rect 15945 13685 15979 13719
rect 16313 13685 16347 13719
rect 20637 13685 20671 13719
rect 21833 13685 21867 13719
rect 22477 13685 22511 13719
rect 24685 13685 24719 13719
rect 25421 13685 25455 13719
rect 1593 13481 1627 13515
rect 1961 13481 1995 13515
rect 2329 13481 2363 13515
rect 3617 13481 3651 13515
rect 4261 13481 4295 13515
rect 4445 13481 4479 13515
rect 4905 13481 4939 13515
rect 6469 13481 6503 13515
rect 7941 13481 7975 13515
rect 8493 13481 8527 13515
rect 13829 13481 13863 13515
rect 14381 13481 14415 13515
rect 18705 13481 18739 13515
rect 21097 13481 21131 13515
rect 22753 13481 22787 13515
rect 23765 13481 23799 13515
rect 24225 13481 24259 13515
rect 25605 13481 25639 13515
rect 5917 13413 5951 13447
rect 7389 13413 7423 13447
rect 9321 13413 9355 13447
rect 12716 13413 12750 13447
rect 17018 13413 17052 13447
rect 24317 13413 24351 13447
rect 1409 13345 1443 13379
rect 2513 13345 2547 13379
rect 4813 13345 4847 13379
rect 5549 13345 5583 13379
rect 6377 13345 6411 13379
rect 8401 13345 8435 13379
rect 9965 13345 9999 13379
rect 10232 13345 10266 13379
rect 12449 13345 12483 13379
rect 16773 13345 16807 13379
rect 19625 13345 19659 13379
rect 21373 13345 21407 13379
rect 21640 13345 21674 13379
rect 25421 13345 25455 13379
rect 4997 13277 5031 13311
rect 6561 13277 6595 13311
rect 7021 13277 7055 13311
rect 8677 13277 8711 13311
rect 15761 13277 15795 13311
rect 19073 13277 19107 13311
rect 19717 13277 19751 13311
rect 19809 13277 19843 13311
rect 24409 13277 24443 13311
rect 2697 13209 2731 13243
rect 8033 13209 8067 13243
rect 3157 13141 3191 13175
rect 6009 13141 6043 13175
rect 11345 13141 11379 13175
rect 12173 13141 12207 13175
rect 15485 13141 15519 13175
rect 16313 13141 16347 13175
rect 18153 13141 18187 13175
rect 19257 13141 19291 13175
rect 20361 13141 20395 13175
rect 23397 13141 23431 13175
rect 23857 13141 23891 13175
rect 1593 12937 1627 12971
rect 3065 12937 3099 12971
rect 3525 12937 3559 12971
rect 4261 12937 4295 12971
rect 4721 12937 4755 12971
rect 5181 12937 5215 12971
rect 6193 12937 6227 12971
rect 6837 12937 6871 12971
rect 8125 12937 8159 12971
rect 8493 12937 8527 12971
rect 8769 12937 8803 12971
rect 9321 12937 9355 12971
rect 10333 12937 10367 12971
rect 10793 12937 10827 12971
rect 13553 12937 13587 12971
rect 15025 12937 15059 12971
rect 16313 12937 16347 12971
rect 16405 12937 16439 12971
rect 16865 12937 16899 12971
rect 17141 12937 17175 12971
rect 18061 12937 18095 12971
rect 19349 12937 19383 12971
rect 20177 12937 20211 12971
rect 21373 12937 21407 12971
rect 21925 12937 21959 12971
rect 23673 12937 23707 12971
rect 24685 12937 24719 12971
rect 25053 12937 25087 12971
rect 2421 12869 2455 12903
rect 3801 12869 3835 12903
rect 15117 12869 15151 12903
rect 5733 12801 5767 12835
rect 6561 12801 6595 12835
rect 7389 12801 7423 12835
rect 9873 12801 9907 12835
rect 12541 12801 12575 12835
rect 14197 12801 14231 12835
rect 14657 12801 14691 12835
rect 15761 12801 15795 12835
rect 23489 12869 23523 12903
rect 26157 12869 26191 12903
rect 17509 12801 17543 12835
rect 18613 12801 18647 12835
rect 20729 12801 20763 12835
rect 22385 12801 22419 12835
rect 22569 12801 22603 12835
rect 23121 12801 23155 12835
rect 24225 12801 24259 12835
rect 1409 12733 1443 12767
rect 2513 12733 2547 12767
rect 3617 12733 3651 12767
rect 5549 12733 5583 12767
rect 7205 12733 7239 12767
rect 9781 12733 9815 12767
rect 13461 12733 13495 12767
rect 14013 12733 14047 12767
rect 15485 12733 15519 12767
rect 15577 12733 15611 12767
rect 16313 12733 16347 12767
rect 16957 12733 16991 12767
rect 17877 12733 17911 12767
rect 18521 12733 18555 12767
rect 19717 12733 19751 12767
rect 20637 12733 20671 12767
rect 24041 12733 24075 12767
rect 25237 12733 25271 12767
rect 25789 12733 25823 12767
rect 7297 12665 7331 12699
rect 10977 12665 11011 12699
rect 12173 12665 12207 12699
rect 13921 12665 13955 12699
rect 20085 12665 20119 12699
rect 20545 12665 20579 12699
rect 2053 12597 2087 12631
rect 2697 12597 2731 12631
rect 4997 12597 5031 12631
rect 5641 12597 5675 12631
rect 9137 12597 9171 12631
rect 9689 12597 9723 12631
rect 13001 12597 13035 12631
rect 18429 12597 18463 12631
rect 21833 12597 21867 12631
rect 22293 12597 22327 12631
rect 24133 12597 24167 12631
rect 25421 12597 25455 12631
rect 1593 12393 1627 12427
rect 2053 12393 2087 12427
rect 2329 12393 2363 12427
rect 2697 12393 2731 12427
rect 2973 12393 3007 12427
rect 3893 12393 3927 12427
rect 4813 12393 4847 12427
rect 5641 12393 5675 12427
rect 6929 12393 6963 12427
rect 8953 12393 8987 12427
rect 9413 12393 9447 12427
rect 12909 12393 12943 12427
rect 13553 12393 13587 12427
rect 20361 12393 20395 12427
rect 21189 12393 21223 12427
rect 24685 12393 24719 12427
rect 24869 12393 24903 12427
rect 25237 12393 25271 12427
rect 4537 12325 4571 12359
rect 7665 12325 7699 12359
rect 10149 12325 10183 12359
rect 21925 12325 21959 12359
rect 25329 12325 25363 12359
rect 1409 12257 1443 12291
rect 2513 12257 2547 12291
rect 5273 12257 5307 12291
rect 6009 12257 6043 12291
rect 6101 12257 6135 12291
rect 7573 12257 7607 12291
rect 10057 12257 10091 12291
rect 11796 12257 11830 12291
rect 15301 12257 15335 12291
rect 15568 12257 15602 12291
rect 18604 12257 18638 12291
rect 21281 12257 21315 12291
rect 22293 12257 22327 12291
rect 22652 12257 22686 12291
rect 6193 12189 6227 12223
rect 7757 12189 7791 12223
rect 10241 12189 10275 12223
rect 11529 12189 11563 12223
rect 14197 12189 14231 12223
rect 18337 12189 18371 12223
rect 20729 12189 20763 12223
rect 22385 12189 22419 12223
rect 25421 12189 25455 12223
rect 7205 12121 7239 12155
rect 8677 12121 8711 12155
rect 9689 12121 9723 12155
rect 10885 12121 10919 12155
rect 21465 12121 21499 12155
rect 23765 12121 23799 12155
rect 24317 12121 24351 12155
rect 8309 12053 8343 12087
rect 11253 12053 11287 12087
rect 14013 12053 14047 12087
rect 15117 12053 15151 12087
rect 16681 12053 16715 12087
rect 17325 12053 17359 12087
rect 18153 12053 18187 12087
rect 19717 12053 19751 12087
rect 1593 11849 1627 11883
rect 1869 11849 1903 11883
rect 2605 11849 2639 11883
rect 4997 11849 5031 11883
rect 6101 11849 6135 11883
rect 7205 11849 7239 11883
rect 7573 11849 7607 11883
rect 9229 11849 9263 11883
rect 10241 11849 10275 11883
rect 10793 11849 10827 11883
rect 11805 11849 11839 11883
rect 15761 11849 15795 11883
rect 21833 11849 21867 11883
rect 22661 11849 22695 11883
rect 23029 11849 23063 11883
rect 23673 11849 23707 11883
rect 25421 11849 25455 11883
rect 26157 11849 26191 11883
rect 4629 11781 4663 11815
rect 7665 11781 7699 11815
rect 14657 11781 14691 11815
rect 24961 11781 24995 11815
rect 5273 11713 5307 11747
rect 6653 11713 6687 11747
rect 8125 11713 8159 11747
rect 8309 11713 8343 11747
rect 9137 11713 9171 11747
rect 9781 11713 9815 11747
rect 11253 11713 11287 11747
rect 11437 11713 11471 11747
rect 16221 11713 16255 11747
rect 16405 11713 16439 11747
rect 16865 11713 16899 11747
rect 17509 11713 17543 11747
rect 18613 11713 18647 11747
rect 24225 11713 24259 11747
rect 1409 11645 1443 11679
rect 2237 11645 2271 11679
rect 5733 11645 5767 11679
rect 8033 11645 8067 11679
rect 8769 11645 8803 11679
rect 9597 11645 9631 11679
rect 10701 11645 10735 11679
rect 11161 11645 11195 11679
rect 13093 11645 13127 11679
rect 13277 11645 13311 11679
rect 17693 11645 17727 11679
rect 18521 11645 18555 11679
rect 19901 11645 19935 11679
rect 22477 11645 22511 11679
rect 24041 11645 24075 11679
rect 25237 11645 25271 11679
rect 25789 11645 25823 11679
rect 9689 11577 9723 11611
rect 12173 11577 12207 11611
rect 12817 11577 12851 11611
rect 13522 11577 13556 11611
rect 16129 11577 16163 11611
rect 19073 11577 19107 11611
rect 19717 11577 19751 11611
rect 20168 11577 20202 11611
rect 24133 11577 24167 11611
rect 15301 11509 15335 11543
rect 17693 11509 17727 11543
rect 17785 11509 17819 11543
rect 18061 11509 18095 11543
rect 18429 11509 18463 11543
rect 21281 11509 21315 11543
rect 22385 11509 22419 11543
rect 23489 11509 23523 11543
rect 1685 11305 1719 11339
rect 5181 11305 5215 11339
rect 6101 11305 6135 11339
rect 7297 11305 7331 11339
rect 8401 11305 8435 11339
rect 9321 11305 9355 11339
rect 10149 11305 10183 11339
rect 11069 11305 11103 11339
rect 14381 11305 14415 11339
rect 16681 11305 16715 11339
rect 17325 11305 17359 11339
rect 18153 11305 18187 11339
rect 21189 11305 21223 11339
rect 23489 11305 23523 11339
rect 24041 11305 24075 11339
rect 25605 11305 25639 11339
rect 7665 11237 7699 11271
rect 9689 11237 9723 11271
rect 11529 11237 11563 11271
rect 15117 11237 15151 11271
rect 15568 11237 15602 11271
rect 17785 11237 17819 11271
rect 22017 11237 22051 11271
rect 22354 11237 22388 11271
rect 8493 11169 8527 11203
rect 11437 11169 11471 11203
rect 13001 11169 13035 11203
rect 14197 11169 14231 11203
rect 15301 11169 15335 11203
rect 18604 11169 18638 11203
rect 21005 11169 21039 11203
rect 24961 11169 24995 11203
rect 8585 11101 8619 11135
rect 11713 11101 11747 11135
rect 12173 11101 12207 11135
rect 13093 11101 13127 11135
rect 13185 11101 13219 11135
rect 18337 11101 18371 11135
rect 22109 11101 22143 11135
rect 25053 11101 25087 11135
rect 25145 11101 25179 11135
rect 5733 11033 5767 11067
rect 8033 11033 8067 11067
rect 10885 11033 10919 11067
rect 12633 11033 12667 11067
rect 19717 11033 19751 11067
rect 20269 11033 20303 11067
rect 21649 11033 21683 11067
rect 12541 10965 12575 10999
rect 24593 10965 24627 10999
rect 8125 10761 8159 10795
rect 8493 10761 8527 10795
rect 9229 10761 9263 10795
rect 10793 10761 10827 10795
rect 12265 10761 12299 10795
rect 13829 10761 13863 10795
rect 14381 10761 14415 10795
rect 17049 10761 17083 10795
rect 18245 10761 18279 10795
rect 19625 10761 19659 10795
rect 20913 10761 20947 10795
rect 23029 10761 23063 10795
rect 23489 10761 23523 10795
rect 25053 10761 25087 10795
rect 25421 10761 25455 10795
rect 7757 10693 7791 10727
rect 10333 10693 10367 10727
rect 17509 10693 17543 10727
rect 19993 10693 20027 10727
rect 23673 10693 23707 10727
rect 9781 10625 9815 10659
rect 11253 10625 11287 10659
rect 11437 10625 11471 10659
rect 12449 10625 12483 10659
rect 15485 10625 15519 10659
rect 18705 10625 18739 10659
rect 18797 10625 18831 10659
rect 21097 10625 21131 10659
rect 24225 10625 24259 10659
rect 9137 10557 9171 10591
rect 9597 10557 9631 10591
rect 12705 10557 12739 10591
rect 14841 10557 14875 10591
rect 16865 10557 16899 10591
rect 17877 10557 17911 10591
rect 19809 10557 19843 10591
rect 24041 10557 24075 10591
rect 25237 10557 25271 10591
rect 25789 10557 25823 10591
rect 10609 10489 10643 10523
rect 11161 10489 11195 10523
rect 15301 10489 15335 10523
rect 16313 10489 16347 10523
rect 20637 10489 20671 10523
rect 21364 10489 21398 10523
rect 9689 10421 9723 10455
rect 11805 10421 11839 10455
rect 14933 10421 14967 10455
rect 15393 10421 15427 10455
rect 16037 10421 16071 10455
rect 16681 10421 16715 10455
rect 18613 10421 18647 10455
rect 19257 10421 19291 10455
rect 22477 10421 22511 10455
rect 24133 10421 24167 10455
rect 24685 10421 24719 10455
rect 9321 10217 9355 10251
rect 10149 10217 10183 10251
rect 11621 10217 11655 10251
rect 14197 10217 14231 10251
rect 15025 10217 15059 10251
rect 15577 10217 15611 10251
rect 23305 10217 23339 10251
rect 24225 10217 24259 10251
rect 25421 10217 25455 10251
rect 10517 10149 10551 10183
rect 12440 10149 12474 10183
rect 16304 10149 16338 10183
rect 20913 10149 20947 10183
rect 24777 10149 24811 10183
rect 10977 10081 11011 10115
rect 11069 10081 11103 10115
rect 12173 10081 12207 10115
rect 16037 10081 16071 10115
rect 19165 10081 19199 10115
rect 21741 10081 21775 10115
rect 22192 10081 22226 10115
rect 11253 10013 11287 10047
rect 18061 10013 18095 10047
rect 19257 10013 19291 10047
rect 19441 10013 19475 10047
rect 21925 10013 21959 10047
rect 24869 10013 24903 10047
rect 24961 10013 24995 10047
rect 8953 9945 8987 9979
rect 10609 9945 10643 9979
rect 11989 9945 12023 9979
rect 18797 9945 18831 9979
rect 19809 9945 19843 9979
rect 24409 9945 24443 9979
rect 13553 9877 13587 9911
rect 17417 9877 17451 9911
rect 18337 9877 18371 9911
rect 20269 9877 20303 9911
rect 23857 9877 23891 9911
rect 12173 9673 12207 9707
rect 13553 9673 13587 9707
rect 15117 9673 15151 9707
rect 22661 9673 22695 9707
rect 24133 9673 24167 9707
rect 10057 9605 10091 9639
rect 11161 9605 11195 9639
rect 16221 9605 16255 9639
rect 17233 9605 17267 9639
rect 20269 9605 20303 9639
rect 24777 9605 24811 9639
rect 25145 9605 25179 9639
rect 10701 9537 10735 9571
rect 13737 9537 13771 9571
rect 16865 9537 16899 9571
rect 22201 9537 22235 9571
rect 10517 9469 10551 9503
rect 15761 9469 15795 9503
rect 16589 9469 16623 9503
rect 18337 9469 18371 9503
rect 21557 9469 21591 9503
rect 22017 9469 22051 9503
rect 24593 9469 24627 9503
rect 25513 9469 25547 9503
rect 13277 9401 13311 9435
rect 14004 9401 14038 9435
rect 16129 9401 16163 9435
rect 18582 9401 18616 9435
rect 21189 9401 21223 9435
rect 22109 9401 22143 9435
rect 24409 9401 24443 9435
rect 9873 9333 9907 9367
rect 10425 9333 10459 9367
rect 11529 9333 11563 9367
rect 11897 9333 11931 9367
rect 12541 9333 12575 9367
rect 16681 9333 16715 9367
rect 17785 9333 17819 9367
rect 19717 9333 19751 9367
rect 21649 9333 21683 9367
rect 10057 9129 10091 9163
rect 10701 9129 10735 9163
rect 11989 9129 12023 9163
rect 12449 9129 12483 9163
rect 13093 9129 13127 9163
rect 13921 9129 13955 9163
rect 15577 9129 15611 9163
rect 16957 9129 16991 9163
rect 19533 9129 19567 9163
rect 20545 9129 20579 9163
rect 20913 9129 20947 9163
rect 22477 9129 22511 9163
rect 22845 9129 22879 9163
rect 24777 9129 24811 9163
rect 14565 9061 14599 9095
rect 22017 9061 22051 9095
rect 22937 9061 22971 9095
rect 10977 8993 11011 9027
rect 12357 8993 12391 9027
rect 14013 8993 14047 9027
rect 15945 8993 15979 9027
rect 17408 8993 17442 9027
rect 21281 8993 21315 9027
rect 24593 8993 24627 9027
rect 12633 8925 12667 8959
rect 14197 8925 14231 8959
rect 15117 8925 15151 8959
rect 16037 8925 16071 8959
rect 16129 8925 16163 8959
rect 17141 8925 17175 8959
rect 19625 8925 19659 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 23121 8925 23155 8959
rect 13553 8857 13587 8891
rect 18521 8857 18555 8891
rect 19073 8857 19107 8891
rect 13369 8789 13403 8823
rect 16589 8789 16623 8823
rect 12633 8585 12667 8619
rect 12909 8585 12943 8619
rect 13921 8585 13955 8619
rect 15669 8585 15703 8619
rect 17417 8585 17451 8619
rect 18981 8585 19015 8619
rect 20545 8585 20579 8619
rect 21557 8585 21591 8619
rect 22937 8585 22971 8619
rect 23397 8585 23431 8619
rect 24133 8585 24167 8619
rect 24869 8585 24903 8619
rect 25145 8585 25179 8619
rect 14473 8517 14507 8551
rect 16405 8517 16439 8551
rect 19993 8517 20027 8551
rect 22661 8517 22695 8551
rect 23857 8517 23891 8551
rect 11345 8449 11379 8483
rect 13461 8449 13495 8483
rect 15025 8449 15059 8483
rect 16957 8449 16991 8483
rect 17785 8449 17819 8483
rect 19533 8449 19567 8483
rect 21005 8449 21039 8483
rect 21097 8449 21131 8483
rect 22109 8449 22143 8483
rect 13277 8381 13311 8415
rect 14933 8381 14967 8415
rect 16773 8381 16807 8415
rect 18521 8381 18555 8415
rect 19349 8381 19383 8415
rect 23673 8381 23707 8415
rect 24685 8381 24719 8415
rect 25513 8381 25547 8415
rect 11989 8313 12023 8347
rect 14381 8313 14415 8347
rect 14841 8313 14875 8347
rect 16865 8313 16899 8347
rect 18797 8313 18831 8347
rect 19441 8313 19475 8347
rect 20453 8313 20487 8347
rect 20913 8313 20947 8347
rect 11253 8245 11287 8279
rect 13369 8245 13403 8279
rect 16313 8245 16347 8279
rect 11897 8041 11931 8075
rect 13001 8041 13035 8075
rect 13645 8041 13679 8075
rect 14197 8041 14231 8075
rect 14749 8041 14783 8075
rect 15117 8041 15151 8075
rect 16405 8041 16439 8075
rect 18981 8041 19015 8075
rect 20637 8041 20671 8075
rect 21465 8041 21499 8075
rect 22937 8041 22971 8075
rect 23949 8041 23983 8075
rect 24961 8041 24995 8075
rect 16037 7973 16071 8007
rect 19349 7973 19383 8007
rect 12265 7905 12299 7939
rect 16764 7905 16798 7939
rect 20913 7905 20947 7939
rect 22753 7905 22787 7939
rect 23765 7905 23799 7939
rect 24777 7905 24811 7939
rect 12357 7837 12391 7871
rect 12449 7837 12483 7871
rect 15485 7837 15519 7871
rect 16497 7837 16531 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 17877 7769 17911 7803
rect 21097 7769 21131 7803
rect 14013 7701 14047 7735
rect 11529 7497 11563 7531
rect 14841 7497 14875 7531
rect 15301 7497 15335 7531
rect 15577 7497 15611 7531
rect 16405 7497 16439 7531
rect 18061 7497 18095 7531
rect 19073 7497 19107 7531
rect 19625 7497 19659 7531
rect 20637 7497 20671 7531
rect 21005 7497 21039 7531
rect 22937 7497 22971 7531
rect 24501 7497 24535 7531
rect 25145 7497 25179 7531
rect 16221 7429 16255 7463
rect 23857 7429 23891 7463
rect 15945 7361 15979 7395
rect 16957 7361 16991 7395
rect 17509 7361 17543 7395
rect 18705 7361 18739 7395
rect 20085 7361 20119 7395
rect 20269 7361 20303 7395
rect 21189 7361 21223 7395
rect 22385 7361 22419 7395
rect 24685 7361 24719 7395
rect 12725 7293 12759 7327
rect 15393 7293 15427 7327
rect 16773 7293 16807 7327
rect 23673 7293 23707 7327
rect 24133 7293 24167 7327
rect 17785 7225 17819 7259
rect 18521 7225 18555 7259
rect 19533 7225 19567 7259
rect 19993 7225 20027 7259
rect 11897 7157 11931 7191
rect 16865 7157 16899 7191
rect 18429 7157 18463 7191
rect 17509 6953 17543 6987
rect 20085 6953 20119 6987
rect 15945 6885 15979 6919
rect 17601 6885 17635 6919
rect 16037 6817 16071 6851
rect 16681 6817 16715 6851
rect 19073 6817 19107 6851
rect 19717 6817 19751 6851
rect 23673 6817 23707 6851
rect 16221 6749 16255 6783
rect 17693 6749 17727 6783
rect 15577 6681 15611 6715
rect 16957 6681 16991 6715
rect 23857 6681 23891 6715
rect 17141 6613 17175 6647
rect 18245 6613 18279 6647
rect 15577 6409 15611 6443
rect 15945 6409 15979 6443
rect 16405 6409 16439 6443
rect 16773 6409 16807 6443
rect 17509 6409 17543 6443
rect 23857 6409 23891 6443
rect 17141 6069 17175 6103
rect 14289 2601 14323 2635
rect 12449 2533 12483 2567
rect 13176 2465 13210 2499
rect 11989 2397 12023 2431
rect 12909 2397 12943 2431
<< metal1 >>
rect 13446 27004 13452 27056
rect 13504 27044 13510 27056
rect 15378 27044 15384 27056
rect 13504 27016 15384 27044
rect 13504 27004 13510 27016
rect 15378 27004 15384 27016
rect 15436 27004 15442 27056
rect 12437 26299 12495 26305
rect 12437 26265 12449 26299
rect 12483 26296 12495 26299
rect 15565 26299 15623 26305
rect 15565 26296 15577 26299
rect 12483 26268 15577 26296
rect 12483 26265 12495 26268
rect 12437 26259 12495 26265
rect 15565 26265 15577 26268
rect 15611 26265 15623 26299
rect 15565 26259 15623 26265
rect 10042 26188 10048 26240
rect 10100 26228 10106 26240
rect 14826 26228 14832 26240
rect 10100 26200 14832 26228
rect 10100 26188 10106 26200
rect 14826 26188 14832 26200
rect 14884 26188 14890 26240
rect 11606 26120 11612 26172
rect 11664 26160 11670 26172
rect 19978 26160 19984 26172
rect 11664 26132 19984 26160
rect 11664 26120 11670 26132
rect 19978 26120 19984 26132
rect 20036 26120 20042 26172
rect 12066 26052 12072 26104
rect 12124 26092 12130 26104
rect 12437 26095 12495 26101
rect 12437 26092 12449 26095
rect 12124 26064 12449 26092
rect 12124 26052 12130 26064
rect 12437 26061 12449 26064
rect 12483 26061 12495 26095
rect 12437 26055 12495 26061
rect 9582 25984 9588 26036
rect 9640 26024 9646 26036
rect 18138 26024 18144 26036
rect 9640 25996 18144 26024
rect 9640 25984 9646 25996
rect 18138 25984 18144 25996
rect 18196 25984 18202 26036
rect 2682 25916 2688 25968
rect 2740 25956 2746 25968
rect 17494 25956 17500 25968
rect 2740 25928 17500 25956
rect 2740 25916 2746 25928
rect 17494 25916 17500 25928
rect 17552 25916 17558 25968
rect 2222 25848 2228 25900
rect 2280 25888 2286 25900
rect 6270 25888 6276 25900
rect 2280 25860 6276 25888
rect 2280 25848 2286 25860
rect 6270 25848 6276 25860
rect 6328 25848 6334 25900
rect 10962 25848 10968 25900
rect 11020 25888 11026 25900
rect 20898 25888 20904 25900
rect 11020 25860 20904 25888
rect 11020 25848 11026 25860
rect 20898 25848 20904 25860
rect 20956 25848 20962 25900
rect 3786 25780 3792 25832
rect 3844 25820 3850 25832
rect 6454 25820 6460 25832
rect 3844 25792 6460 25820
rect 3844 25780 3850 25792
rect 6454 25780 6460 25792
rect 6512 25780 6518 25832
rect 8662 25780 8668 25832
rect 8720 25820 8726 25832
rect 11974 25820 11980 25832
rect 8720 25792 11980 25820
rect 8720 25780 8726 25792
rect 11974 25780 11980 25792
rect 12032 25780 12038 25832
rect 12802 25780 12808 25832
rect 12860 25820 12866 25832
rect 22646 25820 22652 25832
rect 12860 25792 22652 25820
rect 12860 25780 12866 25792
rect 22646 25780 22652 25792
rect 22704 25780 22710 25832
rect 1946 25712 1952 25764
rect 2004 25752 2010 25764
rect 15565 25755 15623 25761
rect 2004 25724 12572 25752
rect 2004 25712 2010 25724
rect 3142 25644 3148 25696
rect 3200 25684 3206 25696
rect 12434 25684 12440 25696
rect 3200 25656 12440 25684
rect 3200 25644 3206 25656
rect 12434 25644 12440 25656
rect 12492 25644 12498 25696
rect 12544 25684 12572 25724
rect 15565 25721 15577 25755
rect 15611 25752 15623 25755
rect 19058 25752 19064 25764
rect 15611 25724 19064 25752
rect 15611 25721 15623 25724
rect 15565 25715 15623 25721
rect 19058 25712 19064 25724
rect 19116 25712 19122 25764
rect 17218 25684 17224 25696
rect 12544 25656 17224 25684
rect 17218 25644 17224 25656
rect 17276 25644 17282 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1946 25480 1952 25492
rect 1907 25452 1952 25480
rect 1946 25440 1952 25452
rect 2004 25440 2010 25492
rect 2869 25483 2927 25489
rect 2869 25449 2881 25483
rect 2915 25480 2927 25483
rect 3602 25480 3608 25492
rect 2915 25452 3608 25480
rect 2915 25449 2927 25452
rect 2869 25443 2927 25449
rect 3602 25440 3608 25452
rect 3660 25440 3666 25492
rect 4798 25480 4804 25492
rect 4759 25452 4804 25480
rect 4798 25440 4804 25452
rect 4856 25440 4862 25492
rect 7101 25483 7159 25489
rect 7101 25449 7113 25483
rect 7147 25449 7159 25483
rect 7101 25443 7159 25449
rect 3050 25372 3056 25424
rect 3108 25412 3114 25424
rect 7116 25412 7144 25443
rect 7282 25440 7288 25492
rect 7340 25480 7346 25492
rect 7469 25483 7527 25489
rect 7469 25480 7481 25483
rect 7340 25452 7481 25480
rect 7340 25440 7346 25452
rect 7469 25449 7481 25452
rect 7515 25449 7527 25483
rect 10962 25480 10968 25492
rect 10923 25452 10968 25480
rect 7469 25443 7527 25449
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 12066 25480 12072 25492
rect 12027 25452 12072 25480
rect 12066 25440 12072 25452
rect 12124 25440 12130 25492
rect 12161 25483 12219 25489
rect 12161 25449 12173 25483
rect 12207 25480 12219 25483
rect 12621 25483 12679 25489
rect 12621 25480 12633 25483
rect 12207 25452 12633 25480
rect 12207 25449 12219 25452
rect 12161 25443 12219 25449
rect 12621 25449 12633 25452
rect 12667 25449 12679 25483
rect 12621 25443 12679 25449
rect 14461 25483 14519 25489
rect 14461 25449 14473 25483
rect 14507 25480 14519 25483
rect 17770 25480 17776 25492
rect 14507 25452 17776 25480
rect 14507 25449 14519 25452
rect 14461 25443 14519 25449
rect 17770 25440 17776 25452
rect 17828 25440 17834 25492
rect 18509 25483 18567 25489
rect 18509 25449 18521 25483
rect 18555 25480 18567 25483
rect 20070 25480 20076 25492
rect 18555 25452 20076 25480
rect 18555 25449 18567 25452
rect 18509 25443 18567 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 20165 25483 20223 25489
rect 20165 25449 20177 25483
rect 20211 25480 20223 25483
rect 21818 25480 21824 25492
rect 20211 25452 21824 25480
rect 20211 25449 20223 25452
rect 20165 25443 20223 25449
rect 21818 25440 21824 25452
rect 21876 25440 21882 25492
rect 22646 25480 22652 25492
rect 22607 25452 22652 25480
rect 22646 25440 22652 25452
rect 22704 25440 22710 25492
rect 23017 25483 23075 25489
rect 23017 25449 23029 25483
rect 23063 25449 23075 25483
rect 23750 25480 23756 25492
rect 23711 25452 23756 25480
rect 23017 25443 23075 25449
rect 3108 25384 7144 25412
rect 11333 25415 11391 25421
rect 3108 25372 3114 25384
rect 11333 25381 11345 25415
rect 11379 25412 11391 25415
rect 11698 25412 11704 25424
rect 11379 25384 11704 25412
rect 11379 25381 11391 25384
rect 11333 25375 11391 25381
rect 11698 25372 11704 25384
rect 11756 25412 11762 25424
rect 11756 25384 12388 25412
rect 11756 25372 11762 25384
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2498 25344 2504 25356
rect 1443 25316 2504 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2498 25304 2504 25316
rect 2556 25304 2562 25356
rect 2774 25344 2780 25356
rect 2735 25316 2780 25344
rect 2774 25304 2780 25316
rect 2832 25304 2838 25356
rect 3329 25347 3387 25353
rect 3329 25313 3341 25347
rect 3375 25344 3387 25347
rect 4709 25347 4767 25353
rect 4709 25344 4721 25347
rect 3375 25316 4721 25344
rect 3375 25313 3387 25316
rect 3329 25307 3387 25313
rect 4709 25313 4721 25316
rect 4755 25344 4767 25347
rect 5442 25344 5448 25356
rect 4755 25316 5448 25344
rect 4755 25313 4767 25316
rect 4709 25307 4767 25313
rect 5442 25304 5448 25316
rect 5500 25304 5506 25356
rect 6546 25304 6552 25356
rect 6604 25344 6610 25356
rect 6917 25347 6975 25353
rect 6917 25344 6929 25347
rect 6604 25316 6929 25344
rect 6604 25304 6610 25316
rect 6917 25313 6929 25316
rect 6963 25313 6975 25347
rect 8478 25344 8484 25356
rect 8439 25316 8484 25344
rect 6917 25307 6975 25313
rect 8478 25304 8484 25316
rect 8536 25344 8542 25356
rect 9582 25344 9588 25356
rect 8536 25316 9588 25344
rect 8536 25304 8542 25316
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 9953 25347 10011 25353
rect 9953 25313 9965 25347
rect 9999 25344 10011 25347
rect 12161 25347 12219 25353
rect 12161 25344 12173 25347
rect 9999 25316 10548 25344
rect 9999 25313 10011 25316
rect 9953 25307 10011 25313
rect 2958 25276 2964 25288
rect 2919 25248 2964 25276
rect 2958 25236 2964 25248
rect 3016 25236 3022 25288
rect 4985 25279 5043 25285
rect 4985 25245 4997 25279
rect 5031 25245 5043 25279
rect 4985 25239 5043 25245
rect 1581 25211 1639 25217
rect 1581 25177 1593 25211
rect 1627 25208 1639 25211
rect 5000 25208 5028 25239
rect 8294 25236 8300 25288
rect 8352 25276 8358 25288
rect 8573 25279 8631 25285
rect 8573 25276 8585 25279
rect 8352 25248 8585 25276
rect 8352 25236 8358 25248
rect 8573 25245 8585 25248
rect 8619 25245 8631 25279
rect 8754 25276 8760 25288
rect 8715 25248 8760 25276
rect 8573 25239 8631 25245
rect 8754 25236 8760 25248
rect 8812 25276 8818 25288
rect 9125 25279 9183 25285
rect 9125 25276 9137 25279
rect 8812 25248 9137 25276
rect 8812 25236 8818 25248
rect 9125 25245 9137 25248
rect 9171 25245 9183 25279
rect 9125 25239 9183 25245
rect 5166 25208 5172 25220
rect 1627 25180 4660 25208
rect 5000 25180 5172 25208
rect 1627 25177 1639 25180
rect 1581 25171 1639 25177
rect 1946 25100 1952 25152
rect 2004 25140 2010 25152
rect 2317 25143 2375 25149
rect 2317 25140 2329 25143
rect 2004 25112 2329 25140
rect 2004 25100 2010 25112
rect 2317 25109 2329 25112
rect 2363 25140 2375 25143
rect 2409 25143 2467 25149
rect 2409 25140 2421 25143
rect 2363 25112 2421 25140
rect 2363 25109 2375 25112
rect 2317 25103 2375 25109
rect 2409 25109 2421 25112
rect 2455 25109 2467 25143
rect 2409 25103 2467 25109
rect 2498 25100 2504 25152
rect 2556 25140 2562 25152
rect 3329 25143 3387 25149
rect 3329 25140 3341 25143
rect 2556 25112 3341 25140
rect 2556 25100 2562 25112
rect 3329 25109 3341 25112
rect 3375 25109 3387 25143
rect 3329 25103 3387 25109
rect 3418 25100 3424 25152
rect 3476 25140 3482 25152
rect 3476 25112 3521 25140
rect 3476 25100 3482 25112
rect 3694 25100 3700 25152
rect 3752 25140 3758 25152
rect 3789 25143 3847 25149
rect 3789 25140 3801 25143
rect 3752 25112 3801 25140
rect 3752 25100 3758 25112
rect 3789 25109 3801 25112
rect 3835 25140 3847 25143
rect 4341 25143 4399 25149
rect 4341 25140 4353 25143
rect 3835 25112 4353 25140
rect 3835 25109 3847 25112
rect 3789 25103 3847 25109
rect 4341 25109 4353 25112
rect 4387 25109 4399 25143
rect 4632 25140 4660 25180
rect 5166 25168 5172 25180
rect 5224 25168 5230 25220
rect 5902 25168 5908 25220
rect 5960 25208 5966 25220
rect 5997 25211 6055 25217
rect 5997 25208 6009 25211
rect 5960 25180 6009 25208
rect 5960 25168 5966 25180
rect 5997 25177 6009 25180
rect 6043 25208 6055 25211
rect 8018 25208 8024 25220
rect 6043 25180 8024 25208
rect 6043 25177 6055 25180
rect 5997 25171 6055 25177
rect 8018 25168 8024 25180
rect 8076 25168 8082 25220
rect 10137 25211 10195 25217
rect 10137 25177 10149 25211
rect 10183 25208 10195 25211
rect 10410 25208 10416 25220
rect 10183 25180 10416 25208
rect 10183 25177 10195 25180
rect 10137 25171 10195 25177
rect 10410 25168 10416 25180
rect 10468 25168 10474 25220
rect 5534 25140 5540 25152
rect 4632 25112 5540 25140
rect 4341 25103 4399 25109
rect 5534 25100 5540 25112
rect 5592 25140 5598 25152
rect 5629 25143 5687 25149
rect 5629 25140 5641 25143
rect 5592 25112 5641 25140
rect 5592 25100 5598 25112
rect 5629 25109 5641 25112
rect 5675 25109 5687 25143
rect 5629 25103 5687 25109
rect 6457 25143 6515 25149
rect 6457 25109 6469 25143
rect 6503 25140 6515 25143
rect 6638 25140 6644 25152
rect 6503 25112 6644 25140
rect 6503 25109 6515 25112
rect 6457 25103 6515 25109
rect 6638 25100 6644 25112
rect 6696 25100 6702 25152
rect 7006 25100 7012 25152
rect 7064 25140 7070 25152
rect 7650 25140 7656 25152
rect 7064 25112 7656 25140
rect 7064 25100 7070 25112
rect 7650 25100 7656 25112
rect 7708 25140 7714 25152
rect 7837 25143 7895 25149
rect 7837 25140 7849 25143
rect 7708 25112 7849 25140
rect 7708 25100 7714 25112
rect 7837 25109 7849 25112
rect 7883 25109 7895 25143
rect 7837 25103 7895 25109
rect 8113 25143 8171 25149
rect 8113 25109 8125 25143
rect 8159 25140 8171 25143
rect 8938 25140 8944 25152
rect 8159 25112 8944 25140
rect 8159 25109 8171 25112
rect 8113 25103 8171 25109
rect 8938 25100 8944 25112
rect 8996 25100 9002 25152
rect 10520 25149 10548 25316
rect 11440 25316 12173 25344
rect 10686 25236 10692 25288
rect 10744 25276 10750 25288
rect 11440 25285 11468 25316
rect 12161 25313 12173 25316
rect 12207 25313 12219 25347
rect 12161 25307 12219 25313
rect 11425 25279 11483 25285
rect 11425 25276 11437 25279
rect 10744 25248 11437 25276
rect 10744 25236 10750 25248
rect 11425 25245 11437 25248
rect 11471 25245 11483 25279
rect 11425 25239 11483 25245
rect 11514 25236 11520 25288
rect 11572 25276 11578 25288
rect 11572 25248 11617 25276
rect 11572 25236 11578 25248
rect 10505 25143 10563 25149
rect 10505 25109 10517 25143
rect 10551 25140 10563 25143
rect 11974 25140 11980 25152
rect 10551 25112 11980 25140
rect 10551 25109 10563 25112
rect 10505 25103 10563 25109
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12360 25140 12388 25384
rect 13262 25372 13268 25424
rect 13320 25412 13326 25424
rect 13320 25384 15148 25412
rect 13320 25372 13326 25384
rect 12437 25347 12495 25353
rect 12437 25313 12449 25347
rect 12483 25344 12495 25347
rect 12802 25344 12808 25356
rect 12483 25316 12808 25344
rect 12483 25313 12495 25316
rect 12437 25307 12495 25313
rect 12802 25304 12808 25316
rect 12860 25344 12866 25356
rect 12989 25347 13047 25353
rect 12989 25344 13001 25347
rect 12860 25316 13001 25344
rect 12860 25304 12866 25316
rect 12989 25313 13001 25316
rect 13035 25313 13047 25347
rect 12989 25307 13047 25313
rect 14277 25347 14335 25353
rect 14277 25313 14289 25347
rect 14323 25344 14335 25347
rect 14458 25344 14464 25356
rect 14323 25316 14464 25344
rect 14323 25313 14335 25316
rect 14277 25307 14335 25313
rect 14458 25304 14464 25316
rect 14516 25304 14522 25356
rect 15120 25344 15148 25384
rect 15470 25372 15476 25424
rect 15528 25412 15534 25424
rect 15841 25415 15899 25421
rect 15841 25412 15853 25415
rect 15528 25384 15853 25412
rect 15528 25372 15534 25384
rect 15841 25381 15853 25384
rect 15887 25412 15899 25415
rect 16942 25412 16948 25424
rect 15887 25384 16948 25412
rect 15887 25381 15899 25384
rect 15841 25375 15899 25381
rect 16942 25372 16948 25384
rect 17000 25372 17006 25424
rect 21545 25415 21603 25421
rect 21545 25412 21557 25415
rect 17052 25384 21557 25412
rect 17052 25344 17080 25384
rect 21545 25381 21557 25384
rect 21591 25412 21603 25415
rect 21591 25384 21772 25412
rect 21591 25381 21603 25384
rect 21545 25375 21603 25381
rect 15120 25316 17080 25344
rect 17129 25347 17187 25353
rect 17129 25313 17141 25347
rect 17175 25344 17187 25347
rect 17678 25344 17684 25356
rect 17175 25316 17684 25344
rect 17175 25313 17187 25316
rect 17129 25307 17187 25313
rect 17678 25304 17684 25316
rect 17736 25304 17742 25356
rect 18322 25344 18328 25356
rect 18283 25316 18328 25344
rect 18322 25304 18328 25316
rect 18380 25304 18386 25356
rect 19978 25344 19984 25356
rect 19939 25316 19984 25344
rect 19978 25304 19984 25316
rect 20036 25344 20042 25356
rect 21744 25353 21772 25384
rect 20533 25347 20591 25353
rect 20533 25344 20545 25347
rect 20036 25316 20545 25344
rect 20036 25304 20042 25316
rect 20533 25313 20545 25316
rect 20579 25313 20591 25347
rect 20533 25307 20591 25313
rect 21729 25347 21787 25353
rect 21729 25313 21741 25347
rect 21775 25313 21787 25347
rect 22664 25344 22692 25440
rect 23032 25412 23060 25443
rect 23750 25440 23756 25452
rect 23808 25440 23814 25492
rect 24213 25483 24271 25489
rect 24213 25449 24225 25483
rect 24259 25480 24271 25483
rect 25866 25480 25872 25492
rect 24259 25452 25872 25480
rect 24259 25449 24271 25452
rect 24213 25443 24271 25449
rect 25866 25440 25872 25452
rect 25924 25440 25930 25492
rect 25314 25412 25320 25424
rect 23032 25384 25320 25412
rect 25314 25372 25320 25384
rect 25372 25372 25378 25424
rect 22833 25347 22891 25353
rect 22833 25344 22845 25347
rect 22664 25316 22845 25344
rect 21729 25307 21787 25313
rect 22833 25313 22845 25316
rect 22879 25313 22891 25347
rect 22833 25307 22891 25313
rect 23842 25304 23848 25356
rect 23900 25344 23906 25356
rect 24029 25347 24087 25353
rect 24029 25344 24041 25347
rect 23900 25316 24041 25344
rect 23900 25304 23906 25316
rect 24029 25313 24041 25316
rect 24075 25313 24087 25347
rect 25130 25344 25136 25356
rect 25091 25316 25136 25344
rect 24029 25307 24087 25313
rect 25130 25304 25136 25316
rect 25188 25304 25194 25356
rect 12894 25236 12900 25288
rect 12952 25276 12958 25288
rect 13081 25279 13139 25285
rect 13081 25276 13093 25279
rect 12952 25248 13093 25276
rect 12952 25236 12958 25248
rect 13081 25245 13093 25248
rect 13127 25245 13139 25279
rect 13081 25239 13139 25245
rect 13170 25236 13176 25288
rect 13228 25276 13234 25288
rect 13265 25279 13323 25285
rect 13265 25276 13277 25279
rect 13228 25248 13277 25276
rect 13228 25236 13234 25248
rect 13265 25245 13277 25248
rect 13311 25276 13323 25279
rect 15930 25276 15936 25288
rect 13311 25248 15424 25276
rect 15891 25248 15936 25276
rect 13311 25245 13323 25248
rect 13265 25239 13323 25245
rect 15105 25211 15163 25217
rect 15105 25177 15117 25211
rect 15151 25208 15163 25211
rect 15286 25208 15292 25220
rect 15151 25180 15292 25208
rect 15151 25177 15163 25180
rect 15105 25171 15163 25177
rect 15286 25168 15292 25180
rect 15344 25168 15350 25220
rect 15396 25208 15424 25248
rect 15930 25236 15936 25248
rect 15988 25236 15994 25288
rect 16114 25276 16120 25288
rect 16075 25248 16120 25276
rect 16114 25236 16120 25248
rect 16172 25236 16178 25288
rect 16132 25208 16160 25236
rect 15396 25180 16160 25208
rect 17313 25211 17371 25217
rect 17313 25177 17325 25211
rect 17359 25208 17371 25211
rect 19518 25208 19524 25220
rect 17359 25180 19524 25208
rect 17359 25177 17371 25180
rect 17313 25171 17371 25177
rect 19518 25168 19524 25180
rect 19576 25168 19582 25220
rect 21913 25211 21971 25217
rect 21913 25177 21925 25211
rect 21959 25208 21971 25211
rect 24762 25208 24768 25220
rect 21959 25180 24768 25208
rect 21959 25177 21971 25180
rect 21913 25171 21971 25177
rect 24762 25168 24768 25180
rect 24820 25168 24826 25220
rect 15473 25143 15531 25149
rect 15473 25140 15485 25143
rect 12360 25112 15485 25140
rect 15473 25109 15485 25112
rect 15519 25109 15531 25143
rect 16574 25140 16580 25152
rect 16535 25112 16580 25140
rect 15473 25103 15531 25109
rect 16574 25100 16580 25112
rect 16632 25100 16638 25152
rect 18046 25140 18052 25152
rect 18007 25112 18052 25140
rect 18046 25100 18052 25112
rect 18104 25100 18110 25152
rect 22373 25143 22431 25149
rect 22373 25109 22385 25143
rect 22419 25140 22431 25143
rect 22922 25140 22928 25152
rect 22419 25112 22928 25140
rect 22419 25109 22431 25112
rect 22373 25103 22431 25109
rect 22922 25100 22928 25112
rect 22980 25100 22986 25152
rect 24670 25100 24676 25152
rect 24728 25140 24734 25152
rect 25317 25143 25375 25149
rect 25317 25140 25329 25143
rect 24728 25112 25329 25140
rect 24728 25100 24734 25112
rect 25317 25109 25329 25112
rect 25363 25109 25375 25143
rect 25317 25103 25375 25109
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1578 24896 1584 24948
rect 1636 24936 1642 24948
rect 18322 24936 18328 24948
rect 1636 24908 18328 24936
rect 1636 24896 1642 24908
rect 18322 24896 18328 24908
rect 18380 24936 18386 24948
rect 18509 24939 18567 24945
rect 18509 24936 18521 24939
rect 18380 24908 18521 24936
rect 18380 24896 18386 24908
rect 18509 24905 18521 24908
rect 18555 24905 18567 24939
rect 18874 24936 18880 24948
rect 18835 24908 18880 24936
rect 18509 24899 18567 24905
rect 18874 24896 18880 24908
rect 18932 24896 18938 24948
rect 1486 24828 1492 24880
rect 1544 24868 1550 24880
rect 2498 24868 2504 24880
rect 1544 24840 2504 24868
rect 1544 24828 1550 24840
rect 2498 24828 2504 24840
rect 2556 24828 2562 24880
rect 2685 24871 2743 24877
rect 2685 24837 2697 24871
rect 2731 24868 2743 24871
rect 2774 24868 2780 24880
rect 2731 24840 2780 24868
rect 2731 24837 2743 24840
rect 2685 24831 2743 24837
rect 2774 24828 2780 24840
rect 2832 24828 2838 24880
rect 4798 24828 4804 24880
rect 4856 24868 4862 24880
rect 5077 24871 5135 24877
rect 5077 24868 5089 24871
rect 4856 24840 5089 24868
rect 4856 24828 4862 24840
rect 5077 24837 5089 24840
rect 5123 24837 5135 24871
rect 5442 24868 5448 24880
rect 5403 24840 5448 24868
rect 5077 24831 5135 24837
rect 5442 24828 5448 24840
rect 5500 24828 5506 24880
rect 10686 24868 10692 24880
rect 10647 24840 10692 24868
rect 10686 24828 10692 24840
rect 10744 24828 10750 24880
rect 11517 24871 11575 24877
rect 11517 24837 11529 24871
rect 11563 24868 11575 24871
rect 11606 24868 11612 24880
rect 11563 24840 11612 24868
rect 11563 24837 11575 24840
rect 11517 24831 11575 24837
rect 11606 24828 11612 24840
rect 11664 24828 11670 24880
rect 12894 24828 12900 24880
rect 12952 24868 12958 24880
rect 16114 24868 16120 24880
rect 12952 24840 13768 24868
rect 16075 24840 16120 24868
rect 12952 24828 12958 24840
rect 2038 24800 2044 24812
rect 1999 24772 2044 24800
rect 2038 24760 2044 24772
rect 2096 24760 2102 24812
rect 2222 24800 2228 24812
rect 2183 24772 2228 24800
rect 2222 24760 2228 24772
rect 2280 24760 2286 24812
rect 7466 24800 7472 24812
rect 7427 24772 7472 24800
rect 7466 24760 7472 24772
rect 7524 24760 7530 24812
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24800 11943 24803
rect 13170 24800 13176 24812
rect 11931 24772 13176 24800
rect 11931 24769 11943 24772
rect 11885 24763 11943 24769
rect 13170 24760 13176 24772
rect 13228 24760 13234 24812
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24769 13691 24803
rect 13740 24800 13768 24840
rect 16114 24828 16120 24840
rect 16172 24828 16178 24880
rect 16850 24828 16856 24880
rect 16908 24868 16914 24880
rect 25130 24868 25136 24880
rect 16908 24840 25136 24868
rect 16908 24828 16914 24840
rect 25130 24828 25136 24840
rect 25188 24868 25194 24880
rect 25777 24871 25835 24877
rect 25777 24868 25789 24871
rect 25188 24840 25789 24868
rect 25188 24828 25194 24840
rect 25777 24837 25789 24840
rect 25823 24837 25835 24871
rect 25777 24831 25835 24837
rect 14369 24803 14427 24809
rect 14369 24800 14381 24803
rect 13740 24772 14381 24800
rect 13633 24763 13691 24769
rect 14369 24769 14381 24772
rect 14415 24769 14427 24803
rect 15194 24800 15200 24812
rect 14369 24763 14427 24769
rect 14476 24772 15200 24800
rect 1946 24732 1952 24744
rect 1907 24704 1952 24732
rect 1946 24692 1952 24704
rect 2004 24692 2010 24744
rect 3145 24735 3203 24741
rect 3145 24701 3157 24735
rect 3191 24732 3203 24735
rect 3234 24732 3240 24744
rect 3191 24704 3240 24732
rect 3191 24701 3203 24704
rect 3145 24695 3203 24701
rect 3234 24692 3240 24704
rect 3292 24692 3298 24744
rect 3418 24741 3424 24744
rect 3412 24732 3424 24741
rect 3379 24704 3424 24732
rect 3412 24695 3424 24704
rect 3418 24692 3424 24695
rect 3476 24692 3482 24744
rect 5534 24692 5540 24744
rect 5592 24732 5598 24744
rect 5629 24735 5687 24741
rect 5629 24732 5641 24735
rect 5592 24704 5641 24732
rect 5592 24692 5598 24704
rect 5629 24701 5641 24704
rect 5675 24701 5687 24735
rect 5629 24695 5687 24701
rect 7282 24692 7288 24744
rect 7340 24732 7346 24744
rect 7377 24735 7435 24741
rect 7377 24732 7389 24735
rect 7340 24704 7389 24732
rect 7340 24692 7346 24704
rect 7377 24701 7389 24704
rect 7423 24701 7435 24735
rect 8570 24732 8576 24744
rect 8531 24704 8576 24732
rect 7377 24695 7435 24701
rect 8570 24692 8576 24704
rect 8628 24692 8634 24744
rect 11333 24735 11391 24741
rect 11333 24701 11345 24735
rect 11379 24732 11391 24735
rect 12066 24732 12072 24744
rect 11379 24704 12072 24732
rect 11379 24701 11391 24704
rect 11333 24695 11391 24701
rect 12066 24692 12072 24704
rect 12124 24692 12130 24744
rect 12897 24735 12955 24741
rect 12897 24701 12909 24735
rect 12943 24732 12955 24735
rect 12986 24732 12992 24744
rect 12943 24704 12992 24732
rect 12943 24701 12955 24704
rect 12897 24695 12955 24701
rect 12986 24692 12992 24704
rect 13044 24732 13050 24744
rect 13446 24732 13452 24744
rect 13044 24704 13452 24732
rect 13044 24692 13050 24704
rect 13446 24692 13452 24704
rect 13504 24692 13510 24744
rect 13648 24732 13676 24763
rect 13648 24704 14044 24732
rect 2866 24624 2872 24676
rect 2924 24664 2930 24676
rect 6086 24664 6092 24676
rect 2924 24636 6092 24664
rect 2924 24624 2930 24636
rect 6086 24624 6092 24636
rect 6144 24624 6150 24676
rect 6273 24667 6331 24673
rect 6273 24633 6285 24667
rect 6319 24664 6331 24667
rect 6319 24636 7328 24664
rect 6319 24633 6331 24636
rect 6273 24627 6331 24633
rect 7300 24608 7328 24636
rect 7926 24624 7932 24676
rect 7984 24664 7990 24676
rect 8754 24664 8760 24676
rect 7984 24636 8760 24664
rect 7984 24624 7990 24636
rect 8754 24624 8760 24636
rect 8812 24673 8818 24676
rect 8812 24667 8876 24673
rect 8812 24633 8830 24667
rect 8864 24664 8876 24667
rect 9858 24664 9864 24676
rect 8864 24636 9864 24664
rect 8864 24633 8876 24636
rect 8812 24627 8876 24633
rect 8812 24624 8818 24627
rect 9858 24624 9864 24636
rect 9916 24624 9922 24676
rect 12253 24667 12311 24673
rect 12253 24633 12265 24667
rect 12299 24664 12311 24667
rect 12299 24636 13400 24664
rect 12299 24633 12311 24636
rect 12253 24627 12311 24633
rect 13372 24608 13400 24636
rect 14016 24608 14044 24704
rect 14366 24624 14372 24676
rect 14424 24664 14430 24676
rect 14476 24664 14504 24772
rect 15194 24760 15200 24772
rect 15252 24800 15258 24812
rect 15657 24803 15715 24809
rect 15657 24800 15669 24803
rect 15252 24772 15669 24800
rect 15252 24760 15258 24772
rect 15657 24769 15669 24772
rect 15703 24800 15715 24803
rect 18322 24800 18328 24812
rect 15703 24772 18328 24800
rect 15703 24769 15715 24772
rect 15657 24763 15715 24769
rect 18322 24760 18328 24772
rect 18380 24760 18386 24812
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24800 20131 24803
rect 20717 24803 20775 24809
rect 20717 24800 20729 24803
rect 20119 24772 20729 24800
rect 20119 24769 20131 24772
rect 20073 24763 20131 24769
rect 20717 24769 20729 24772
rect 20763 24800 20775 24803
rect 20990 24800 20996 24812
rect 20763 24772 20996 24800
rect 20763 24769 20775 24772
rect 20717 24763 20775 24769
rect 20990 24760 20996 24772
rect 21048 24760 21054 24812
rect 21542 24800 21548 24812
rect 21455 24772 21548 24800
rect 21542 24760 21548 24772
rect 21600 24800 21606 24812
rect 22649 24803 22707 24809
rect 21600 24772 22600 24800
rect 21600 24760 21606 24772
rect 14921 24735 14979 24741
rect 14921 24701 14933 24735
rect 14967 24732 14979 24735
rect 16574 24732 16580 24744
rect 14967 24704 15516 24732
rect 16487 24704 16580 24732
rect 14967 24701 14979 24704
rect 14921 24695 14979 24701
rect 14424 24636 14504 24664
rect 14424 24624 14430 24636
rect 14550 24624 14556 24676
rect 14608 24664 14614 24676
rect 15378 24664 15384 24676
rect 14608 24636 15056 24664
rect 15339 24636 15384 24664
rect 14608 24624 14614 24636
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 1854 24596 1860 24608
rect 1627 24568 1860 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 1854 24556 1860 24568
rect 1912 24556 1918 24608
rect 1946 24556 1952 24608
rect 2004 24596 2010 24608
rect 2774 24596 2780 24608
rect 2004 24568 2780 24596
rect 2004 24556 2010 24568
rect 2774 24556 2780 24568
rect 2832 24556 2838 24608
rect 3053 24599 3111 24605
rect 3053 24565 3065 24599
rect 3099 24596 3111 24599
rect 3602 24596 3608 24608
rect 3099 24568 3608 24596
rect 3099 24565 3111 24568
rect 3053 24559 3111 24565
rect 3602 24556 3608 24568
rect 3660 24556 3666 24608
rect 3878 24556 3884 24608
rect 3936 24596 3942 24608
rect 4525 24599 4583 24605
rect 4525 24596 4537 24599
rect 3936 24568 4537 24596
rect 3936 24556 3942 24568
rect 4525 24565 4537 24568
rect 4571 24565 4583 24599
rect 4525 24559 4583 24565
rect 5813 24599 5871 24605
rect 5813 24565 5825 24599
rect 5859 24596 5871 24599
rect 5994 24596 6000 24608
rect 5859 24568 6000 24596
rect 5859 24565 5871 24568
rect 5813 24559 5871 24565
rect 5994 24556 6000 24568
rect 6052 24556 6058 24608
rect 6546 24596 6552 24608
rect 6507 24568 6552 24596
rect 6546 24556 6552 24568
rect 6604 24556 6610 24608
rect 6917 24599 6975 24605
rect 6917 24565 6929 24599
rect 6963 24596 6975 24599
rect 7190 24596 7196 24608
rect 6963 24568 7196 24596
rect 6963 24565 6975 24568
rect 6917 24559 6975 24565
rect 7190 24556 7196 24568
rect 7248 24556 7254 24608
rect 7282 24556 7288 24608
rect 7340 24596 7346 24608
rect 8110 24596 8116 24608
rect 7340 24568 7385 24596
rect 8071 24568 8116 24596
rect 7340 24556 7346 24568
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 9950 24596 9956 24608
rect 9911 24568 9956 24596
rect 9950 24556 9956 24568
rect 10008 24556 10014 24608
rect 11057 24599 11115 24605
rect 11057 24565 11069 24599
rect 11103 24596 11115 24599
rect 11422 24596 11428 24608
rect 11103 24568 11428 24596
rect 11103 24565 11115 24568
rect 11057 24559 11115 24565
rect 11422 24556 11428 24568
rect 11480 24556 11486 24608
rect 12802 24556 12808 24608
rect 12860 24596 12866 24608
rect 12989 24599 13047 24605
rect 12989 24596 13001 24599
rect 12860 24568 13001 24596
rect 12860 24556 12866 24568
rect 12989 24565 13001 24568
rect 13035 24565 13047 24599
rect 13354 24596 13360 24608
rect 13315 24568 13360 24596
rect 12989 24559 13047 24565
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 13998 24596 14004 24608
rect 13959 24568 14004 24596
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 15028 24605 15056 24636
rect 15378 24624 15384 24636
rect 15436 24624 15442 24676
rect 15488 24608 15516 24704
rect 16574 24692 16580 24704
rect 16632 24692 16638 24744
rect 16942 24692 16948 24744
rect 17000 24732 17006 24744
rect 17129 24735 17187 24741
rect 17129 24732 17141 24735
rect 17000 24704 17141 24732
rect 17000 24692 17006 24704
rect 17129 24701 17141 24704
rect 17175 24701 17187 24735
rect 18046 24732 18052 24744
rect 18007 24704 18052 24732
rect 17129 24695 17187 24701
rect 18046 24692 18052 24704
rect 18104 24692 18110 24744
rect 18874 24692 18880 24744
rect 18932 24732 18938 24744
rect 19061 24735 19119 24741
rect 19061 24732 19073 24735
rect 18932 24704 19073 24732
rect 18932 24692 18938 24704
rect 19061 24701 19073 24704
rect 19107 24701 19119 24735
rect 19061 24695 19119 24701
rect 16592 24664 16620 24692
rect 20625 24667 20683 24673
rect 20625 24664 20637 24667
rect 16592 24636 18276 24664
rect 15013 24599 15071 24605
rect 15013 24565 15025 24599
rect 15059 24565 15071 24599
rect 15470 24596 15476 24608
rect 15431 24568 15476 24596
rect 15013 24559 15071 24565
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 15930 24556 15936 24608
rect 15988 24596 15994 24608
rect 16393 24599 16451 24605
rect 16393 24596 16405 24599
rect 15988 24568 16405 24596
rect 15988 24556 15994 24568
rect 16393 24565 16405 24568
rect 16439 24565 16451 24599
rect 16758 24596 16764 24608
rect 16719 24568 16764 24596
rect 16393 24559 16451 24565
rect 16758 24556 16764 24568
rect 16816 24556 16822 24608
rect 17589 24599 17647 24605
rect 17589 24565 17601 24599
rect 17635 24596 17647 24599
rect 17678 24596 17684 24608
rect 17635 24568 17684 24596
rect 17635 24565 17647 24568
rect 17589 24559 17647 24565
rect 17678 24556 17684 24568
rect 17736 24556 17742 24608
rect 18248 24605 18276 24636
rect 19628 24636 20637 24664
rect 18233 24599 18291 24605
rect 18233 24565 18245 24599
rect 18279 24565 18291 24599
rect 19242 24596 19248 24608
rect 19203 24568 19248 24596
rect 18233 24559 18291 24565
rect 19242 24556 19248 24568
rect 19300 24556 19306 24608
rect 19518 24556 19524 24608
rect 19576 24596 19582 24608
rect 19628 24605 19656 24636
rect 20625 24633 20637 24636
rect 20671 24633 20683 24667
rect 20625 24627 20683 24633
rect 20806 24624 20812 24676
rect 20864 24664 20870 24676
rect 21821 24667 21879 24673
rect 21821 24664 21833 24667
rect 20864 24636 21833 24664
rect 20864 24624 20870 24636
rect 21821 24633 21833 24636
rect 21867 24664 21879 24667
rect 22373 24667 22431 24673
rect 21867 24636 22324 24664
rect 21867 24633 21879 24636
rect 21821 24627 21879 24633
rect 19613 24599 19671 24605
rect 19613 24596 19625 24599
rect 19576 24568 19625 24596
rect 19576 24556 19582 24568
rect 19613 24565 19625 24568
rect 19659 24565 19671 24599
rect 20162 24596 20168 24608
rect 20123 24568 20168 24596
rect 19613 24559 19671 24565
rect 20162 24556 20168 24568
rect 20220 24556 20226 24608
rect 20530 24596 20536 24608
rect 20491 24568 20536 24596
rect 20530 24556 20536 24568
rect 20588 24556 20594 24608
rect 21910 24556 21916 24608
rect 21968 24596 21974 24608
rect 22005 24599 22063 24605
rect 22005 24596 22017 24599
rect 21968 24568 22017 24596
rect 21968 24556 21974 24568
rect 22005 24565 22017 24568
rect 22051 24565 22063 24599
rect 22296 24596 22324 24636
rect 22373 24633 22385 24667
rect 22419 24664 22431 24667
rect 22572 24664 22600 24772
rect 22649 24769 22661 24803
rect 22695 24800 22707 24803
rect 22922 24800 22928 24812
rect 22695 24772 22928 24800
rect 22695 24769 22707 24772
rect 22649 24763 22707 24769
rect 22922 24760 22928 24772
rect 22980 24760 22986 24812
rect 23474 24800 23480 24812
rect 23387 24772 23480 24800
rect 23474 24760 23480 24772
rect 23532 24800 23538 24812
rect 24302 24800 24308 24812
rect 23532 24772 24164 24800
rect 24263 24772 24308 24800
rect 23532 24760 23538 24772
rect 24136 24744 24164 24772
rect 24302 24760 24308 24772
rect 24360 24760 24366 24812
rect 23750 24692 23756 24744
rect 23808 24732 23814 24744
rect 24029 24735 24087 24741
rect 24029 24732 24041 24735
rect 23808 24704 24041 24732
rect 23808 24692 23814 24704
rect 24029 24701 24041 24704
rect 24075 24701 24087 24735
rect 24029 24695 24087 24701
rect 24118 24692 24124 24744
rect 24176 24692 24182 24744
rect 25133 24735 25191 24741
rect 25133 24701 25145 24735
rect 25179 24732 25191 24735
rect 25225 24735 25283 24741
rect 25225 24732 25237 24735
rect 25179 24704 25237 24732
rect 25179 24701 25191 24704
rect 25133 24695 25191 24701
rect 25225 24701 25237 24704
rect 25271 24732 25283 24735
rect 25774 24732 25780 24744
rect 25271 24704 25780 24732
rect 25271 24701 25283 24704
rect 25225 24695 25283 24701
rect 25774 24692 25780 24704
rect 25832 24692 25838 24744
rect 22646 24664 22652 24676
rect 22419 24636 22652 24664
rect 22419 24633 22431 24636
rect 22373 24627 22431 24633
rect 22646 24624 22652 24636
rect 22704 24664 22710 24676
rect 23198 24664 23204 24676
rect 22704 24636 23204 24664
rect 22704 24624 22710 24636
rect 23198 24624 23204 24636
rect 23256 24624 23262 24676
rect 23842 24624 23848 24676
rect 23900 24664 23906 24676
rect 24673 24667 24731 24673
rect 24673 24664 24685 24667
rect 23900 24636 24685 24664
rect 23900 24624 23906 24636
rect 24673 24633 24685 24636
rect 24719 24633 24731 24667
rect 24673 24627 24731 24633
rect 22462 24596 22468 24608
rect 22296 24568 22468 24596
rect 22005 24559 22063 24565
rect 22462 24556 22468 24568
rect 22520 24556 22526 24608
rect 22922 24556 22928 24608
rect 22980 24596 22986 24608
rect 23017 24599 23075 24605
rect 23017 24596 23029 24599
rect 22980 24568 23029 24596
rect 22980 24556 22986 24568
rect 23017 24565 23029 24568
rect 23063 24565 23075 24599
rect 23017 24559 23075 24565
rect 23661 24599 23719 24605
rect 23661 24565 23673 24599
rect 23707 24596 23719 24599
rect 23750 24596 23756 24608
rect 23707 24568 23756 24596
rect 23707 24565 23719 24568
rect 23661 24559 23719 24565
rect 23750 24556 23756 24568
rect 23808 24556 23814 24608
rect 24121 24599 24179 24605
rect 24121 24565 24133 24599
rect 24167 24596 24179 24599
rect 24210 24596 24216 24608
rect 24167 24568 24216 24596
rect 24167 24565 24179 24568
rect 24121 24559 24179 24565
rect 24210 24556 24216 24568
rect 24268 24556 24274 24608
rect 25406 24596 25412 24608
rect 25367 24568 25412 24596
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1578 24392 1584 24404
rect 1539 24364 1584 24392
rect 1578 24352 1584 24364
rect 1636 24352 1642 24404
rect 1949 24395 2007 24401
rect 1949 24361 1961 24395
rect 1995 24392 2007 24395
rect 2038 24392 2044 24404
rect 1995 24364 2044 24392
rect 1995 24361 2007 24364
rect 1949 24355 2007 24361
rect 2038 24352 2044 24364
rect 2096 24352 2102 24404
rect 2314 24392 2320 24404
rect 2275 24364 2320 24392
rect 2314 24352 2320 24364
rect 2372 24352 2378 24404
rect 2866 24392 2872 24404
rect 2827 24364 2872 24392
rect 2866 24352 2872 24364
rect 2924 24352 2930 24404
rect 3234 24352 3240 24404
rect 3292 24392 3298 24404
rect 3421 24395 3479 24401
rect 3421 24392 3433 24395
rect 3292 24364 3433 24392
rect 3292 24352 3298 24364
rect 3421 24361 3433 24364
rect 3467 24361 3479 24395
rect 3878 24392 3884 24404
rect 3839 24364 3884 24392
rect 3421 24355 3479 24361
rect 3878 24352 3884 24364
rect 3936 24352 3942 24404
rect 4430 24392 4436 24404
rect 4391 24364 4436 24392
rect 4430 24352 4436 24364
rect 4488 24352 4494 24404
rect 7006 24392 7012 24404
rect 4908 24364 7012 24392
rect 2130 24284 2136 24336
rect 2188 24324 2194 24336
rect 4908 24324 4936 24364
rect 7006 24352 7012 24364
rect 7064 24352 7070 24404
rect 8478 24352 8484 24404
rect 8536 24392 8542 24404
rect 8665 24395 8723 24401
rect 8665 24392 8677 24395
rect 8536 24364 8677 24392
rect 8536 24352 8542 24364
rect 8665 24361 8677 24364
rect 8711 24361 8723 24395
rect 8665 24355 8723 24361
rect 9950 24352 9956 24404
rect 10008 24392 10014 24404
rect 10137 24395 10195 24401
rect 10137 24392 10149 24395
rect 10008 24364 10149 24392
rect 10008 24352 10014 24364
rect 10137 24361 10149 24364
rect 10183 24361 10195 24395
rect 10686 24392 10692 24404
rect 10647 24364 10692 24392
rect 10137 24355 10195 24361
rect 10686 24352 10692 24364
rect 10744 24352 10750 24404
rect 11146 24392 11152 24404
rect 11107 24364 11152 24392
rect 11146 24352 11152 24364
rect 11204 24352 11210 24404
rect 11698 24392 11704 24404
rect 11659 24364 11704 24392
rect 11698 24352 11704 24364
rect 11756 24352 11762 24404
rect 13446 24352 13452 24404
rect 13504 24392 13510 24404
rect 16850 24392 16856 24404
rect 13504 24364 16856 24392
rect 13504 24352 13510 24364
rect 16850 24352 16856 24364
rect 16908 24352 16914 24404
rect 17034 24392 17040 24404
rect 16995 24364 17040 24392
rect 17034 24352 17040 24364
rect 17092 24352 17098 24404
rect 17218 24392 17224 24404
rect 17179 24364 17224 24392
rect 17218 24352 17224 24364
rect 17276 24352 17282 24404
rect 18138 24352 18144 24404
rect 18196 24392 18202 24404
rect 18233 24395 18291 24401
rect 18233 24392 18245 24395
rect 18196 24364 18245 24392
rect 18196 24352 18202 24364
rect 18233 24361 18245 24364
rect 18279 24361 18291 24395
rect 18233 24355 18291 24361
rect 19245 24395 19303 24401
rect 19245 24361 19257 24395
rect 19291 24392 19303 24395
rect 20349 24395 20407 24401
rect 20349 24392 20361 24395
rect 19291 24364 20361 24392
rect 19291 24361 19303 24364
rect 19245 24355 19303 24361
rect 20349 24361 20361 24364
rect 20395 24392 20407 24395
rect 20530 24392 20536 24404
rect 20395 24364 20536 24392
rect 20395 24361 20407 24364
rect 20349 24355 20407 24361
rect 20530 24352 20536 24364
rect 20588 24352 20594 24404
rect 23106 24352 23112 24404
rect 23164 24392 23170 24404
rect 23201 24395 23259 24401
rect 23201 24392 23213 24395
rect 23164 24364 23213 24392
rect 23164 24352 23170 24364
rect 23201 24361 23213 24364
rect 23247 24392 23259 24395
rect 23753 24395 23811 24401
rect 23753 24392 23765 24395
rect 23247 24364 23765 24392
rect 23247 24361 23259 24364
rect 23201 24355 23259 24361
rect 23753 24361 23765 24364
rect 23799 24392 23811 24395
rect 23934 24392 23940 24404
rect 23799 24364 23940 24392
rect 23799 24361 23811 24364
rect 23753 24355 23811 24361
rect 23934 24352 23940 24364
rect 23992 24352 23998 24404
rect 25222 24392 25228 24404
rect 25183 24364 25228 24392
rect 25222 24352 25228 24364
rect 25280 24352 25286 24404
rect 25317 24395 25375 24401
rect 25317 24361 25329 24395
rect 25363 24392 25375 24395
rect 25498 24392 25504 24404
rect 25363 24364 25504 24392
rect 25363 24361 25375 24364
rect 25317 24355 25375 24361
rect 25498 24352 25504 24364
rect 25556 24352 25562 24404
rect 6086 24324 6092 24336
rect 2188 24296 4936 24324
rect 5644 24296 6092 24324
rect 2188 24284 2194 24296
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 2038 24256 2044 24268
rect 1443 24228 2044 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 2038 24216 2044 24228
rect 2096 24216 2102 24268
rect 2314 24216 2320 24268
rect 2372 24256 2378 24268
rect 2590 24256 2596 24268
rect 2372 24228 2596 24256
rect 2372 24216 2378 24228
rect 2590 24216 2596 24228
rect 2648 24216 2654 24268
rect 2777 24259 2835 24265
rect 2777 24225 2789 24259
rect 2823 24256 2835 24259
rect 3326 24256 3332 24268
rect 2823 24228 3332 24256
rect 2823 24225 2835 24228
rect 2777 24219 2835 24225
rect 3326 24216 3332 24228
rect 3384 24216 3390 24268
rect 4522 24256 4528 24268
rect 4483 24228 4528 24256
rect 4522 24216 4528 24228
rect 4580 24216 4586 24268
rect 5644 24265 5672 24296
rect 6086 24284 6092 24296
rect 6144 24284 6150 24336
rect 8570 24284 8576 24336
rect 8628 24324 8634 24336
rect 9033 24327 9091 24333
rect 9033 24324 9045 24327
rect 8628 24296 9045 24324
rect 8628 24284 8634 24296
rect 9033 24293 9045 24296
rect 9079 24324 9091 24327
rect 9582 24324 9588 24336
rect 9079 24296 9588 24324
rect 9079 24293 9091 24296
rect 9033 24287 9091 24293
rect 9582 24284 9588 24296
rect 9640 24284 9646 24336
rect 10962 24284 10968 24336
rect 11020 24324 11026 24336
rect 11057 24327 11115 24333
rect 11057 24324 11069 24327
rect 11020 24296 11069 24324
rect 11020 24284 11026 24296
rect 11057 24293 11069 24296
rect 11103 24324 11115 24327
rect 11238 24324 11244 24336
rect 11103 24296 11244 24324
rect 11103 24293 11115 24296
rect 11057 24287 11115 24293
rect 11238 24284 11244 24296
rect 11296 24284 11302 24336
rect 12066 24284 12072 24336
rect 12124 24324 12130 24336
rect 12621 24327 12679 24333
rect 12621 24324 12633 24327
rect 12124 24296 12633 24324
rect 12124 24284 12130 24296
rect 12621 24293 12633 24296
rect 12667 24293 12679 24327
rect 17052 24324 17080 24352
rect 17052 24296 17816 24324
rect 12621 24287 12679 24293
rect 5629 24259 5687 24265
rect 5629 24225 5641 24259
rect 5675 24225 5687 24259
rect 5896 24259 5954 24265
rect 5896 24256 5908 24259
rect 5629 24219 5687 24225
rect 5736 24228 5908 24256
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24157 3111 24191
rect 4614 24188 4620 24200
rect 4575 24160 4620 24188
rect 3053 24151 3111 24157
rect 3068 24120 3096 24151
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 5166 24188 5172 24200
rect 5079 24160 5172 24188
rect 5166 24148 5172 24160
rect 5224 24188 5230 24200
rect 5736 24188 5764 24228
rect 5896 24225 5908 24228
rect 5942 24256 5954 24259
rect 6362 24256 6368 24268
rect 5942 24228 6368 24256
rect 5942 24225 5954 24228
rect 5896 24219 5954 24225
rect 6362 24216 6368 24228
rect 6420 24216 6426 24268
rect 8113 24259 8171 24265
rect 8113 24225 8125 24259
rect 8159 24256 8171 24259
rect 8202 24256 8208 24268
rect 8159 24228 8208 24256
rect 8159 24225 8171 24228
rect 8113 24219 8171 24225
rect 8202 24216 8208 24228
rect 8260 24216 8266 24268
rect 12710 24256 12716 24268
rect 12671 24228 12716 24256
rect 12710 24216 12716 24228
rect 12768 24216 12774 24268
rect 14093 24259 14151 24265
rect 14093 24225 14105 24259
rect 14139 24256 14151 24259
rect 14642 24256 14648 24268
rect 14139 24228 14648 24256
rect 14139 24225 14151 24228
rect 14093 24219 14151 24225
rect 14642 24216 14648 24228
rect 14700 24216 14706 24268
rect 15286 24216 15292 24268
rect 15344 24256 15350 24268
rect 16025 24259 16083 24265
rect 16025 24256 16037 24259
rect 15344 24228 16037 24256
rect 15344 24216 15350 24228
rect 16025 24225 16037 24228
rect 16071 24225 16083 24259
rect 17586 24256 17592 24268
rect 17547 24228 17592 24256
rect 16025 24219 16083 24225
rect 17586 24216 17592 24228
rect 17644 24216 17650 24268
rect 5224 24160 5764 24188
rect 5224 24148 5230 24160
rect 9306 24148 9312 24200
rect 9364 24188 9370 24200
rect 9677 24191 9735 24197
rect 9677 24188 9689 24191
rect 9364 24160 9689 24188
rect 9364 24148 9370 24160
rect 9677 24157 9689 24160
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 11333 24191 11391 24197
rect 11333 24157 11345 24191
rect 11379 24188 11391 24191
rect 11698 24188 11704 24200
rect 11379 24160 11704 24188
rect 11379 24157 11391 24160
rect 11333 24151 11391 24157
rect 11698 24148 11704 24160
rect 11756 24148 11762 24200
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24188 12219 24191
rect 12802 24188 12808 24200
rect 12207 24160 12808 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 12802 24148 12808 24160
rect 12860 24148 12866 24200
rect 14734 24148 14740 24200
rect 14792 24188 14798 24200
rect 16117 24191 16175 24197
rect 16117 24188 16129 24191
rect 14792 24160 16129 24188
rect 14792 24148 14798 24160
rect 16117 24157 16129 24160
rect 16163 24157 16175 24191
rect 16298 24188 16304 24200
rect 16259 24160 16304 24188
rect 16117 24151 16175 24157
rect 16298 24148 16304 24160
rect 16356 24148 16362 24200
rect 17788 24197 17816 24296
rect 20162 24284 20168 24336
rect 20220 24324 20226 24336
rect 20625 24327 20683 24333
rect 20625 24324 20637 24327
rect 20220 24296 20637 24324
rect 20220 24284 20226 24296
rect 20625 24293 20637 24296
rect 20671 24324 20683 24327
rect 22005 24327 22063 24333
rect 22005 24324 22017 24327
rect 20671 24296 22017 24324
rect 20671 24293 20683 24296
rect 20625 24287 20683 24293
rect 22005 24293 22017 24296
rect 22051 24293 22063 24327
rect 22005 24287 22063 24293
rect 19613 24259 19671 24265
rect 19613 24225 19625 24259
rect 19659 24256 19671 24259
rect 20346 24256 20352 24268
rect 19659 24228 20352 24256
rect 19659 24225 19671 24228
rect 19613 24219 19671 24225
rect 20346 24216 20352 24228
rect 20404 24216 20410 24268
rect 21818 24216 21824 24268
rect 21876 24256 21882 24268
rect 21913 24259 21971 24265
rect 21913 24256 21925 24259
rect 21876 24228 21925 24256
rect 21876 24216 21882 24228
rect 21913 24225 21925 24228
rect 21959 24225 21971 24259
rect 21913 24219 21971 24225
rect 22830 24216 22836 24268
rect 22888 24256 22894 24268
rect 23661 24259 23719 24265
rect 23661 24256 23673 24259
rect 22888 24228 23673 24256
rect 22888 24216 22894 24228
rect 23661 24225 23673 24228
rect 23707 24225 23719 24259
rect 23661 24219 23719 24225
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24157 17739 24191
rect 17681 24151 17739 24157
rect 17773 24191 17831 24197
rect 17773 24157 17785 24191
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 3510 24120 3516 24132
rect 3068 24092 3516 24120
rect 3510 24080 3516 24092
rect 3568 24120 3574 24132
rect 5184 24120 5212 24148
rect 7926 24120 7932 24132
rect 3568 24092 5212 24120
rect 7887 24092 7932 24120
rect 3568 24080 3574 24092
rect 7926 24080 7932 24092
rect 7984 24080 7990 24132
rect 14274 24120 14280 24132
rect 14235 24092 14280 24120
rect 14274 24080 14280 24092
rect 14332 24080 14338 24132
rect 15013 24123 15071 24129
rect 15013 24120 15025 24123
rect 14384 24092 15025 24120
rect 2406 24052 2412 24064
rect 2367 24024 2412 24052
rect 2406 24012 2412 24024
rect 2464 24012 2470 24064
rect 4062 24052 4068 24064
rect 4023 24024 4068 24052
rect 4062 24012 4068 24024
rect 4120 24012 4126 24064
rect 5534 24052 5540 24064
rect 5495 24024 5540 24052
rect 5534 24012 5540 24024
rect 5592 24012 5598 24064
rect 6914 24012 6920 24064
rect 6972 24052 6978 24064
rect 7009 24055 7067 24061
rect 7009 24052 7021 24055
rect 6972 24024 7021 24052
rect 6972 24012 6978 24024
rect 7009 24021 7021 24024
rect 7055 24021 7067 24055
rect 7009 24015 7067 24021
rect 7098 24012 7104 24064
rect 7156 24052 7162 24064
rect 7466 24052 7472 24064
rect 7156 24024 7472 24052
rect 7156 24012 7162 24024
rect 7466 24012 7472 24024
rect 7524 24052 7530 24064
rect 7561 24055 7619 24061
rect 7561 24052 7573 24055
rect 7524 24024 7573 24052
rect 7524 24012 7530 24024
rect 7561 24021 7573 24024
rect 7607 24021 7619 24055
rect 8294 24052 8300 24064
rect 8255 24024 8300 24052
rect 7561 24015 7619 24021
rect 8294 24012 8300 24024
rect 8352 24012 8358 24064
rect 9490 24052 9496 24064
rect 9451 24024 9496 24052
rect 9490 24012 9496 24024
rect 9548 24012 9554 24064
rect 12250 24052 12256 24064
rect 12211 24024 12256 24052
rect 12250 24012 12256 24024
rect 12308 24012 12314 24064
rect 12986 24012 12992 24064
rect 13044 24052 13050 24064
rect 13265 24055 13323 24061
rect 13265 24052 13277 24055
rect 13044 24024 13277 24052
rect 13044 24012 13050 24024
rect 13265 24021 13277 24024
rect 13311 24021 13323 24055
rect 13265 24015 13323 24021
rect 13906 24012 13912 24064
rect 13964 24052 13970 24064
rect 14384 24052 14412 24092
rect 15013 24089 15025 24092
rect 15059 24120 15071 24123
rect 15378 24120 15384 24132
rect 15059 24092 15384 24120
rect 15059 24089 15071 24092
rect 15013 24083 15071 24089
rect 15378 24080 15384 24092
rect 15436 24080 15442 24132
rect 15565 24123 15623 24129
rect 15565 24089 15577 24123
rect 15611 24120 15623 24123
rect 15746 24120 15752 24132
rect 15611 24092 15752 24120
rect 15611 24089 15623 24092
rect 15565 24083 15623 24089
rect 15746 24080 15752 24092
rect 15804 24080 15810 24132
rect 17696 24120 17724 24151
rect 19334 24148 19340 24200
rect 19392 24188 19398 24200
rect 19705 24191 19763 24197
rect 19705 24188 19717 24191
rect 19392 24160 19717 24188
rect 19392 24148 19398 24160
rect 19705 24157 19717 24160
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24188 19947 24191
rect 19978 24188 19984 24200
rect 19935 24160 19984 24188
rect 19935 24157 19947 24160
rect 19889 24151 19947 24157
rect 17862 24120 17868 24132
rect 17696 24092 17868 24120
rect 17862 24080 17868 24092
rect 17920 24080 17926 24132
rect 18782 24080 18788 24132
rect 18840 24120 18846 24132
rect 19153 24123 19211 24129
rect 19153 24120 19165 24123
rect 18840 24092 19165 24120
rect 18840 24080 18846 24092
rect 19153 24089 19165 24092
rect 19199 24120 19211 24123
rect 19904 24120 19932 24151
rect 19978 24148 19984 24160
rect 20036 24148 20042 24200
rect 21453 24191 21511 24197
rect 21453 24157 21465 24191
rect 21499 24188 21511 24191
rect 21726 24188 21732 24200
rect 21499 24160 21732 24188
rect 21499 24157 21511 24160
rect 21453 24151 21511 24157
rect 21726 24148 21732 24160
rect 21784 24188 21790 24200
rect 22097 24191 22155 24197
rect 22097 24188 22109 24191
rect 21784 24160 22109 24188
rect 21784 24148 21790 24160
rect 22097 24157 22109 24160
rect 22143 24157 22155 24191
rect 22097 24151 22155 24157
rect 22922 24148 22928 24200
rect 22980 24188 22986 24200
rect 23845 24191 23903 24197
rect 23845 24188 23857 24191
rect 22980 24160 23857 24188
rect 22980 24148 22986 24160
rect 23845 24157 23857 24160
rect 23891 24188 23903 24191
rect 24210 24188 24216 24200
rect 23891 24160 24216 24188
rect 23891 24157 23903 24160
rect 23845 24151 23903 24157
rect 24210 24148 24216 24160
rect 24268 24188 24274 24200
rect 24305 24191 24363 24197
rect 24305 24188 24317 24191
rect 24268 24160 24317 24188
rect 24268 24148 24274 24160
rect 24305 24157 24317 24160
rect 24351 24188 24363 24191
rect 25409 24191 25467 24197
rect 25409 24188 25421 24191
rect 24351 24160 25421 24188
rect 24351 24157 24363 24160
rect 24305 24151 24363 24157
rect 25409 24157 25421 24160
rect 25455 24188 25467 24191
rect 25682 24188 25688 24200
rect 25455 24160 25688 24188
rect 25455 24157 25467 24160
rect 25409 24151 25467 24157
rect 25682 24148 25688 24160
rect 25740 24148 25746 24200
rect 19199 24092 19932 24120
rect 19199 24089 19211 24092
rect 19153 24083 19211 24089
rect 21818 24080 21824 24132
rect 21876 24120 21882 24132
rect 22649 24123 22707 24129
rect 22649 24120 22661 24123
rect 21876 24092 22661 24120
rect 21876 24080 21882 24092
rect 22649 24089 22661 24092
rect 22695 24120 22707 24123
rect 23382 24120 23388 24132
rect 22695 24092 23388 24120
rect 22695 24089 22707 24092
rect 22649 24083 22707 24089
rect 23382 24080 23388 24092
rect 23440 24080 23446 24132
rect 13964 24024 14412 24052
rect 13964 24012 13970 24024
rect 14458 24012 14464 24064
rect 14516 24052 14522 24064
rect 14645 24055 14703 24061
rect 14645 24052 14657 24055
rect 14516 24024 14657 24052
rect 14516 24012 14522 24024
rect 14645 24021 14657 24024
rect 14691 24021 14703 24055
rect 14645 24015 14703 24021
rect 15657 24055 15715 24061
rect 15657 24021 15669 24055
rect 15703 24052 15715 24055
rect 16206 24052 16212 24064
rect 15703 24024 16212 24052
rect 15703 24021 15715 24024
rect 15657 24015 15715 24021
rect 16206 24012 16212 24024
rect 16264 24012 16270 24064
rect 21545 24055 21603 24061
rect 21545 24021 21557 24055
rect 21591 24052 21603 24055
rect 22002 24052 22008 24064
rect 21591 24024 22008 24052
rect 21591 24021 21603 24024
rect 21545 24015 21603 24021
rect 22002 24012 22008 24024
rect 22060 24012 22066 24064
rect 23290 24052 23296 24064
rect 23251 24024 23296 24052
rect 23290 24012 23296 24024
rect 23348 24012 23354 24064
rect 24854 24052 24860 24064
rect 24815 24024 24860 24052
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1581 23851 1639 23857
rect 1581 23817 1593 23851
rect 1627 23848 1639 23851
rect 2682 23848 2688 23860
rect 1627 23820 2688 23848
rect 1627 23817 1639 23820
rect 1581 23811 1639 23817
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 3326 23808 3332 23860
rect 3384 23848 3390 23860
rect 3421 23851 3479 23857
rect 3421 23848 3433 23851
rect 3384 23820 3433 23848
rect 3384 23808 3390 23820
rect 3421 23817 3433 23820
rect 3467 23817 3479 23851
rect 3421 23811 3479 23817
rect 4614 23808 4620 23860
rect 4672 23848 4678 23860
rect 5350 23848 5356 23860
rect 4672 23820 5356 23848
rect 4672 23808 4678 23820
rect 5350 23808 5356 23820
rect 5408 23808 5414 23860
rect 9306 23848 9312 23860
rect 9267 23820 9312 23848
rect 9306 23808 9312 23820
rect 9364 23808 9370 23860
rect 9582 23848 9588 23860
rect 9543 23820 9588 23848
rect 9582 23808 9588 23820
rect 9640 23808 9646 23860
rect 12066 23808 12072 23860
rect 12124 23848 12130 23860
rect 12161 23851 12219 23857
rect 12161 23848 12173 23851
rect 12124 23820 12173 23848
rect 12124 23808 12130 23820
rect 12161 23817 12173 23820
rect 12207 23817 12219 23851
rect 12710 23848 12716 23860
rect 12671 23820 12716 23848
rect 12161 23811 12219 23817
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 14734 23808 14740 23860
rect 14792 23848 14798 23860
rect 14921 23851 14979 23857
rect 14921 23848 14933 23851
rect 14792 23820 14933 23848
rect 14792 23808 14798 23820
rect 14921 23817 14933 23820
rect 14967 23817 14979 23851
rect 14921 23811 14979 23817
rect 18141 23851 18199 23857
rect 18141 23817 18153 23851
rect 18187 23848 18199 23851
rect 19518 23848 19524 23860
rect 18187 23820 19524 23848
rect 18187 23817 18199 23820
rect 18141 23811 18199 23817
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 19886 23848 19892 23860
rect 19847 23820 19892 23848
rect 19886 23808 19892 23820
rect 19944 23808 19950 23860
rect 25406 23848 25412 23860
rect 25367 23820 25412 23848
rect 25406 23808 25412 23820
rect 25464 23808 25470 23860
rect 25682 23808 25688 23860
rect 25740 23848 25746 23860
rect 25777 23851 25835 23857
rect 25777 23848 25789 23851
rect 25740 23820 25789 23848
rect 25740 23808 25746 23820
rect 25777 23817 25789 23820
rect 25823 23817 25835 23851
rect 25777 23811 25835 23817
rect 1949 23783 2007 23789
rect 1949 23749 1961 23783
rect 1995 23780 2007 23783
rect 2866 23780 2872 23792
rect 1995 23752 2872 23780
rect 1995 23749 2007 23752
rect 1949 23743 2007 23749
rect 2866 23740 2872 23752
rect 2924 23740 2930 23792
rect 3510 23780 3516 23792
rect 3068 23752 3516 23780
rect 1854 23672 1860 23724
rect 1912 23712 1918 23724
rect 2498 23712 2504 23724
rect 1912 23684 2504 23712
rect 1912 23672 1918 23684
rect 2498 23672 2504 23684
rect 2556 23672 2562 23724
rect 3068 23721 3096 23752
rect 3510 23740 3516 23752
rect 3568 23740 3574 23792
rect 6362 23780 6368 23792
rect 6275 23752 6368 23780
rect 6362 23740 6368 23752
rect 6420 23780 6426 23792
rect 9122 23780 9128 23792
rect 6420 23752 9128 23780
rect 6420 23740 6426 23752
rect 9122 23740 9128 23752
rect 9180 23740 9186 23792
rect 3053 23715 3111 23721
rect 3053 23681 3065 23715
rect 3099 23681 3111 23715
rect 3053 23675 3111 23681
rect 3234 23672 3240 23724
rect 3292 23712 3298 23724
rect 3973 23715 4031 23721
rect 3973 23712 3985 23715
rect 3292 23684 3985 23712
rect 3292 23672 3298 23684
rect 3973 23681 3985 23684
rect 4019 23681 4031 23715
rect 8846 23712 8852 23724
rect 8807 23684 8852 23712
rect 3973 23675 4031 23681
rect 8846 23672 8852 23684
rect 8904 23672 8910 23724
rect 9600 23712 9628 23808
rect 16850 23780 16856 23792
rect 16811 23752 16856 23780
rect 16850 23740 16856 23752
rect 16908 23740 16914 23792
rect 20346 23780 20352 23792
rect 20307 23752 20352 23780
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 24946 23780 24952 23792
rect 24859 23752 24952 23780
rect 24946 23740 24952 23752
rect 25004 23780 25010 23792
rect 25498 23780 25504 23792
rect 25004 23752 25504 23780
rect 25004 23740 25010 23752
rect 25498 23740 25504 23752
rect 25556 23740 25562 23792
rect 9769 23715 9827 23721
rect 9769 23712 9781 23715
rect 9600 23684 9781 23712
rect 9769 23681 9781 23684
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 2130 23644 2136 23656
rect 1443 23616 2136 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 2130 23604 2136 23616
rect 2188 23604 2194 23656
rect 2777 23647 2835 23653
rect 2777 23644 2789 23647
rect 2240 23616 2789 23644
rect 1302 23536 1308 23588
rect 1360 23576 1366 23588
rect 2240 23576 2268 23616
rect 2777 23613 2789 23616
rect 2823 23644 2835 23647
rect 3602 23644 3608 23656
rect 2823 23616 3608 23644
rect 2823 23613 2835 23616
rect 2777 23607 2835 23613
rect 3602 23604 3608 23616
rect 3660 23644 3666 23656
rect 3789 23647 3847 23653
rect 3789 23644 3801 23647
rect 3660 23616 3801 23644
rect 3660 23604 3666 23616
rect 3789 23613 3801 23616
rect 3835 23613 3847 23647
rect 3789 23607 3847 23613
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 8113 23647 8171 23653
rect 6871 23616 7512 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 1360 23548 2268 23576
rect 2317 23579 2375 23585
rect 1360 23536 1366 23548
rect 2317 23545 2329 23579
rect 2363 23576 2375 23579
rect 2363 23548 2912 23576
rect 2363 23545 2375 23548
rect 2317 23539 2375 23545
rect 2409 23511 2467 23517
rect 2409 23477 2421 23511
rect 2455 23508 2467 23511
rect 2682 23508 2688 23520
rect 2455 23480 2688 23508
rect 2455 23477 2467 23480
rect 2409 23471 2467 23477
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 2884 23517 2912 23548
rect 3878 23536 3884 23588
rect 3936 23576 3942 23588
rect 4218 23579 4276 23585
rect 4218 23576 4230 23579
rect 3936 23548 4230 23576
rect 3936 23536 3942 23548
rect 4218 23545 4230 23548
rect 4264 23545 4276 23579
rect 6546 23576 6552 23588
rect 4218 23539 4276 23545
rect 5368 23548 6552 23576
rect 2869 23511 2927 23517
rect 2869 23477 2881 23511
rect 2915 23508 2927 23511
rect 5368 23508 5396 23548
rect 6546 23536 6552 23548
rect 6604 23536 6610 23588
rect 2915 23480 5396 23508
rect 2915 23477 2927 23480
rect 2869 23471 2927 23477
rect 5626 23468 5632 23520
rect 5684 23508 5690 23520
rect 5905 23511 5963 23517
rect 5905 23508 5917 23511
rect 5684 23480 5917 23508
rect 5684 23468 5690 23480
rect 5905 23477 5917 23480
rect 5951 23508 5963 23511
rect 6086 23508 6092 23520
rect 5951 23480 6092 23508
rect 5951 23477 5963 23480
rect 5905 23471 5963 23477
rect 6086 23468 6092 23480
rect 6144 23468 6150 23520
rect 7006 23508 7012 23520
rect 6967 23480 7012 23508
rect 7006 23468 7012 23480
rect 7064 23468 7070 23520
rect 7484 23517 7512 23616
rect 8113 23613 8125 23647
rect 8159 23644 8171 23647
rect 8202 23644 8208 23656
rect 8159 23616 8208 23644
rect 8159 23613 8171 23616
rect 8113 23607 8171 23613
rect 8202 23604 8208 23616
rect 8260 23604 8266 23656
rect 8573 23647 8631 23653
rect 8573 23613 8585 23647
rect 8619 23644 8631 23647
rect 9306 23644 9312 23656
rect 8619 23616 9312 23644
rect 8619 23613 8631 23616
rect 8573 23607 8631 23613
rect 9306 23604 9312 23616
rect 9364 23604 9370 23656
rect 9784 23644 9812 23675
rect 15378 23672 15384 23724
rect 15436 23712 15442 23724
rect 15473 23715 15531 23721
rect 15473 23712 15485 23715
rect 15436 23684 15485 23712
rect 15436 23672 15442 23684
rect 15473 23681 15485 23684
rect 15519 23681 15531 23715
rect 18782 23712 18788 23724
rect 18743 23684 18788 23712
rect 15473 23675 15531 23681
rect 18782 23672 18788 23684
rect 18840 23672 18846 23724
rect 24210 23712 24216 23724
rect 24171 23684 24216 23712
rect 24210 23672 24216 23684
rect 24268 23672 24274 23724
rect 11514 23644 11520 23656
rect 9784 23616 11520 23644
rect 11514 23604 11520 23616
rect 11572 23644 11578 23656
rect 12986 23644 12992 23656
rect 11572 23616 12992 23644
rect 11572 23604 11578 23616
rect 12986 23604 12992 23616
rect 13044 23604 13050 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 13188 23616 17417 23644
rect 9950 23536 9956 23588
rect 10008 23585 10014 23588
rect 10008 23579 10072 23585
rect 10008 23545 10026 23579
rect 10060 23545 10072 23579
rect 13188 23576 13216 23616
rect 17405 23613 17417 23616
rect 17451 23644 17463 23647
rect 17586 23644 17592 23656
rect 17451 23616 17592 23644
rect 17451 23613 17463 23616
rect 17405 23607 17463 23613
rect 17586 23604 17592 23616
rect 17644 23604 17650 23656
rect 18138 23604 18144 23656
rect 18196 23644 18202 23656
rect 18509 23647 18567 23653
rect 18509 23644 18521 23647
rect 18196 23616 18521 23644
rect 18196 23604 18202 23616
rect 18509 23613 18521 23616
rect 18555 23613 18567 23647
rect 18509 23607 18567 23613
rect 19426 23604 19432 23656
rect 19484 23644 19490 23656
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 19484 23616 19717 23644
rect 19484 23604 19490 23616
rect 19705 23613 19717 23616
rect 19751 23613 19763 23647
rect 19705 23607 19763 23613
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23613 20959 23647
rect 20901 23607 20959 23613
rect 10008 23539 10072 23545
rect 10796 23548 13216 23576
rect 13256 23579 13314 23585
rect 10008 23536 10014 23539
rect 10796 23520 10824 23548
rect 13256 23545 13268 23579
rect 13302 23576 13314 23579
rect 13538 23576 13544 23588
rect 13302 23548 13544 23576
rect 13302 23545 13314 23548
rect 13256 23539 13314 23545
rect 13538 23536 13544 23548
rect 13596 23536 13602 23588
rect 14090 23536 14096 23588
rect 14148 23576 14154 23588
rect 15286 23576 15292 23588
rect 14148 23548 15292 23576
rect 14148 23536 14154 23548
rect 15286 23536 15292 23548
rect 15344 23536 15350 23588
rect 15746 23585 15752 23588
rect 15740 23539 15752 23585
rect 15804 23576 15810 23588
rect 17770 23576 17776 23588
rect 15804 23548 15840 23576
rect 17731 23548 17776 23576
rect 15746 23536 15752 23539
rect 15804 23536 15810 23548
rect 17770 23536 17776 23548
rect 17828 23576 17834 23588
rect 18601 23579 18659 23585
rect 18601 23576 18613 23579
rect 17828 23548 18613 23576
rect 17828 23536 17834 23548
rect 18601 23545 18613 23548
rect 18647 23545 18659 23579
rect 18601 23539 18659 23545
rect 7469 23511 7527 23517
rect 7469 23477 7481 23511
rect 7515 23508 7527 23511
rect 7926 23508 7932 23520
rect 7515 23480 7932 23508
rect 7515 23477 7527 23480
rect 7469 23471 7527 23477
rect 7926 23468 7932 23480
rect 7984 23468 7990 23520
rect 8110 23468 8116 23520
rect 8168 23508 8174 23520
rect 8205 23511 8263 23517
rect 8205 23508 8217 23511
rect 8168 23480 8217 23508
rect 8168 23468 8174 23480
rect 8205 23477 8217 23480
rect 8251 23477 8263 23511
rect 8662 23508 8668 23520
rect 8623 23480 8668 23508
rect 8205 23471 8263 23477
rect 8662 23468 8668 23480
rect 8720 23468 8726 23520
rect 9766 23468 9772 23520
rect 9824 23508 9830 23520
rect 10778 23508 10784 23520
rect 9824 23480 10784 23508
rect 9824 23468 9830 23480
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 11054 23468 11060 23520
rect 11112 23508 11118 23520
rect 11149 23511 11207 23517
rect 11149 23508 11161 23511
rect 11112 23480 11161 23508
rect 11112 23468 11118 23480
rect 11149 23477 11161 23480
rect 11195 23477 11207 23511
rect 11790 23508 11796 23520
rect 11751 23480 11796 23508
rect 11149 23471 11207 23477
rect 11790 23468 11796 23480
rect 11848 23508 11854 23520
rect 13998 23508 14004 23520
rect 11848 23480 14004 23508
rect 11848 23468 11854 23480
rect 13998 23468 14004 23480
rect 14056 23508 14062 23520
rect 14369 23511 14427 23517
rect 14369 23508 14381 23511
rect 14056 23480 14381 23508
rect 14056 23468 14062 23480
rect 14369 23477 14381 23480
rect 14415 23477 14427 23511
rect 19334 23508 19340 23520
rect 19295 23480 19340 23508
rect 14369 23471 14427 23477
rect 19334 23468 19340 23480
rect 19392 23468 19398 23520
rect 20809 23511 20867 23517
rect 20809 23477 20821 23511
rect 20855 23508 20867 23511
rect 20916 23508 20944 23607
rect 20990 23604 20996 23656
rect 21048 23644 21054 23656
rect 21157 23647 21215 23653
rect 21157 23644 21169 23647
rect 21048 23616 21169 23644
rect 21048 23604 21054 23616
rect 21157 23613 21169 23616
rect 21203 23613 21215 23647
rect 21157 23607 21215 23613
rect 25225 23647 25283 23653
rect 25225 23613 25237 23647
rect 25271 23644 25283 23647
rect 25682 23644 25688 23656
rect 25271 23616 25688 23644
rect 25271 23613 25283 23616
rect 25225 23607 25283 23613
rect 25682 23604 25688 23616
rect 25740 23644 25746 23656
rect 26145 23647 26203 23653
rect 26145 23644 26157 23647
rect 25740 23616 26157 23644
rect 25740 23604 25746 23616
rect 26145 23613 26157 23616
rect 26191 23613 26203 23647
rect 26145 23607 26203 23613
rect 24029 23579 24087 23585
rect 24029 23576 24041 23579
rect 23584 23548 24041 23576
rect 23584 23520 23612 23548
rect 24029 23545 24041 23548
rect 24075 23545 24087 23579
rect 24029 23539 24087 23545
rect 21450 23508 21456 23520
rect 20855 23480 21456 23508
rect 20855 23477 20867 23480
rect 20809 23471 20867 23477
rect 21450 23468 21456 23480
rect 21508 23468 21514 23520
rect 21726 23468 21732 23520
rect 21784 23508 21790 23520
rect 22281 23511 22339 23517
rect 22281 23508 22293 23511
rect 21784 23480 22293 23508
rect 21784 23468 21790 23480
rect 22281 23477 22293 23480
rect 22327 23477 22339 23511
rect 22281 23471 22339 23477
rect 22830 23468 22836 23520
rect 22888 23508 22894 23520
rect 23017 23511 23075 23517
rect 23017 23508 23029 23511
rect 22888 23480 23029 23508
rect 22888 23468 22894 23480
rect 23017 23477 23029 23480
rect 23063 23477 23075 23511
rect 23017 23471 23075 23477
rect 23477 23511 23535 23517
rect 23477 23477 23489 23511
rect 23523 23508 23535 23511
rect 23566 23508 23572 23520
rect 23523 23480 23572 23508
rect 23523 23477 23535 23480
rect 23477 23471 23535 23477
rect 23566 23468 23572 23480
rect 23624 23468 23630 23520
rect 23661 23511 23719 23517
rect 23661 23477 23673 23511
rect 23707 23508 23719 23511
rect 23934 23508 23940 23520
rect 23707 23480 23940 23508
rect 23707 23477 23719 23480
rect 23661 23471 23719 23477
rect 23934 23468 23940 23480
rect 23992 23468 23998 23520
rect 24118 23508 24124 23520
rect 24079 23480 24124 23508
rect 24118 23468 24124 23480
rect 24176 23468 24182 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 2832 23276 2912 23304
rect 2832 23264 2838 23276
rect 1394 23196 1400 23248
rect 1452 23236 1458 23248
rect 1762 23236 1768 23248
rect 1452 23208 1768 23236
rect 1452 23196 1458 23208
rect 1762 23196 1768 23208
rect 1820 23196 1826 23248
rect 2884 23177 2912 23276
rect 3234 23264 3240 23316
rect 3292 23304 3298 23316
rect 3789 23307 3847 23313
rect 3789 23304 3801 23307
rect 3292 23276 3801 23304
rect 3292 23264 3298 23276
rect 3789 23273 3801 23276
rect 3835 23273 3847 23307
rect 3789 23267 3847 23273
rect 3510 23236 3516 23248
rect 3471 23208 3516 23236
rect 3510 23196 3516 23208
rect 3568 23196 3574 23248
rect 2777 23171 2835 23177
rect 2777 23137 2789 23171
rect 2823 23137 2835 23171
rect 2777 23131 2835 23137
rect 2869 23171 2927 23177
rect 2869 23137 2881 23171
rect 2915 23168 2927 23171
rect 3234 23168 3240 23180
rect 2915 23140 3240 23168
rect 2915 23137 2927 23140
rect 2869 23131 2927 23137
rect 1397 23103 1455 23109
rect 1397 23069 1409 23103
rect 1443 23100 1455 23103
rect 1578 23100 1584 23112
rect 1443 23072 1584 23100
rect 1443 23069 1455 23072
rect 1397 23063 1455 23069
rect 1578 23060 1584 23072
rect 1636 23060 1642 23112
rect 2792 23100 2820 23131
rect 3234 23128 3240 23140
rect 3292 23128 3298 23180
rect 3804 23168 3832 23267
rect 4430 23264 4436 23316
rect 4488 23304 4494 23316
rect 4617 23307 4675 23313
rect 4617 23304 4629 23307
rect 4488 23276 4629 23304
rect 4488 23264 4494 23276
rect 4617 23273 4629 23276
rect 4663 23273 4675 23307
rect 4617 23267 4675 23273
rect 7561 23307 7619 23313
rect 7561 23273 7573 23307
rect 7607 23304 7619 23307
rect 8110 23304 8116 23316
rect 7607 23276 8116 23304
rect 7607 23273 7619 23276
rect 7561 23267 7619 23273
rect 8110 23264 8116 23276
rect 8168 23304 8174 23316
rect 8389 23307 8447 23313
rect 8389 23304 8401 23307
rect 8168 23276 8401 23304
rect 8168 23264 8174 23276
rect 8389 23273 8401 23276
rect 8435 23273 8447 23307
rect 8389 23267 8447 23273
rect 8481 23307 8539 23313
rect 8481 23273 8493 23307
rect 8527 23304 8539 23307
rect 8662 23304 8668 23316
rect 8527 23276 8668 23304
rect 8527 23273 8539 23276
rect 8481 23267 8539 23273
rect 8662 23264 8668 23276
rect 8720 23304 8726 23316
rect 9677 23307 9735 23313
rect 9677 23304 9689 23307
rect 8720 23276 9689 23304
rect 8720 23264 8726 23276
rect 9677 23273 9689 23276
rect 9723 23273 9735 23307
rect 9677 23267 9735 23273
rect 10781 23307 10839 23313
rect 10781 23273 10793 23307
rect 10827 23304 10839 23307
rect 10962 23304 10968 23316
rect 10827 23276 10968 23304
rect 10827 23273 10839 23276
rect 10781 23267 10839 23273
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 11146 23304 11152 23316
rect 11107 23276 11152 23304
rect 11146 23264 11152 23276
rect 11204 23264 11210 23316
rect 12894 23304 12900 23316
rect 12807 23276 12900 23304
rect 12894 23264 12900 23276
rect 12952 23304 12958 23316
rect 13170 23304 13176 23316
rect 12952 23276 13176 23304
rect 12952 23264 12958 23276
rect 13170 23264 13176 23276
rect 13228 23264 13234 23316
rect 18417 23307 18475 23313
rect 18417 23273 18429 23307
rect 18463 23304 18475 23307
rect 18782 23304 18788 23316
rect 18463 23276 18788 23304
rect 18463 23273 18475 23276
rect 18417 23267 18475 23273
rect 18782 23264 18788 23276
rect 18840 23264 18846 23316
rect 20990 23264 20996 23316
rect 21048 23304 21054 23316
rect 21085 23307 21143 23313
rect 21085 23304 21097 23307
rect 21048 23276 21097 23304
rect 21048 23264 21054 23276
rect 21085 23273 21097 23276
rect 21131 23273 21143 23307
rect 21085 23267 21143 23273
rect 23382 23264 23388 23316
rect 23440 23304 23446 23316
rect 23937 23307 23995 23313
rect 23937 23304 23949 23307
rect 23440 23276 23949 23304
rect 23440 23264 23446 23276
rect 23937 23273 23949 23276
rect 23983 23273 23995 23307
rect 23937 23267 23995 23273
rect 24305 23307 24363 23313
rect 24305 23273 24317 23307
rect 24351 23304 24363 23307
rect 24762 23304 24768 23316
rect 24351 23276 24768 23304
rect 24351 23273 24363 23276
rect 24305 23267 24363 23273
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 24946 23304 24952 23316
rect 24859 23276 24952 23304
rect 24946 23264 24952 23276
rect 25004 23304 25010 23316
rect 25222 23304 25228 23316
rect 25004 23276 25228 23304
rect 25004 23264 25010 23276
rect 25222 23264 25228 23276
rect 25280 23264 25286 23316
rect 5626 23236 5632 23248
rect 5000 23208 5632 23236
rect 5000 23180 5028 23208
rect 5626 23196 5632 23208
rect 5684 23196 5690 23248
rect 7834 23236 7840 23248
rect 7795 23208 7840 23236
rect 7834 23196 7840 23208
rect 7892 23196 7898 23248
rect 8846 23196 8852 23248
rect 8904 23236 8910 23248
rect 9125 23239 9183 23245
rect 9125 23236 9137 23239
rect 8904 23208 9137 23236
rect 8904 23196 8910 23208
rect 9125 23205 9137 23208
rect 9171 23236 9183 23239
rect 9398 23236 9404 23248
rect 9171 23208 9404 23236
rect 9171 23205 9183 23208
rect 9125 23199 9183 23205
rect 9398 23196 9404 23208
rect 9456 23236 9462 23248
rect 9950 23236 9956 23248
rect 9456 23208 9956 23236
rect 9456 23196 9462 23208
rect 9950 23196 9956 23208
rect 10008 23236 10014 23248
rect 10008 23208 10272 23236
rect 10008 23196 10014 23208
rect 4893 23171 4951 23177
rect 4893 23168 4905 23171
rect 3804 23140 4905 23168
rect 4893 23137 4905 23140
rect 4939 23168 4951 23171
rect 4982 23168 4988 23180
rect 4939 23140 4988 23168
rect 4939 23137 4951 23140
rect 4893 23131 4951 23137
rect 4982 23128 4988 23140
rect 5040 23128 5046 23180
rect 5160 23171 5218 23177
rect 5160 23137 5172 23171
rect 5206 23168 5218 23171
rect 5442 23168 5448 23180
rect 5206 23140 5448 23168
rect 5206 23137 5218 23140
rect 5160 23131 5218 23137
rect 5442 23128 5448 23140
rect 5500 23128 5506 23180
rect 6914 23168 6920 23180
rect 6875 23140 6920 23168
rect 6914 23128 6920 23140
rect 6972 23128 6978 23180
rect 10042 23168 10048 23180
rect 10003 23140 10048 23168
rect 10042 23128 10048 23140
rect 10100 23128 10106 23180
rect 3050 23100 3056 23112
rect 2792 23072 2912 23100
rect 2963 23072 3056 23100
rect 1670 22992 1676 23044
rect 1728 23032 1734 23044
rect 2884 23032 2912 23072
rect 3050 23060 3056 23072
rect 3108 23100 3114 23112
rect 3418 23100 3424 23112
rect 3108 23072 3424 23100
rect 3108 23060 3114 23072
rect 3418 23060 3424 23072
rect 3476 23060 3482 23112
rect 6546 23060 6552 23112
rect 6604 23100 6610 23112
rect 8110 23100 8116 23112
rect 6604 23072 8116 23100
rect 6604 23060 6610 23072
rect 8110 23060 8116 23072
rect 8168 23060 8174 23112
rect 8665 23103 8723 23109
rect 8665 23069 8677 23103
rect 8711 23100 8723 23103
rect 8754 23100 8760 23112
rect 8711 23072 8760 23100
rect 8711 23069 8723 23072
rect 8665 23063 8723 23069
rect 8754 23060 8760 23072
rect 8812 23060 8818 23112
rect 8938 23060 8944 23112
rect 8996 23100 9002 23112
rect 10244 23109 10272 23208
rect 11974 23196 11980 23248
rect 12032 23236 12038 23248
rect 16292 23239 16350 23245
rect 12032 23208 14863 23236
rect 12032 23196 12038 23208
rect 11514 23168 11520 23180
rect 11475 23140 11520 23168
rect 11514 23128 11520 23140
rect 11572 23128 11578 23180
rect 11790 23177 11796 23180
rect 11784 23168 11796 23177
rect 11751 23140 11796 23168
rect 11784 23131 11796 23140
rect 11790 23128 11796 23131
rect 11848 23128 11854 23180
rect 14093 23171 14151 23177
rect 14093 23137 14105 23171
rect 14139 23168 14151 23171
rect 14734 23168 14740 23180
rect 14139 23140 14740 23168
rect 14139 23137 14151 23140
rect 14093 23131 14151 23137
rect 14734 23128 14740 23140
rect 14792 23128 14798 23180
rect 14835 23168 14863 23208
rect 16292 23205 16304 23239
rect 16338 23236 16350 23239
rect 16390 23236 16396 23248
rect 16338 23208 16396 23236
rect 16338 23205 16350 23208
rect 16292 23199 16350 23205
rect 16390 23196 16396 23208
rect 16448 23196 16454 23248
rect 17954 23236 17960 23248
rect 17915 23208 17960 23236
rect 17954 23196 17960 23208
rect 18012 23196 18018 23248
rect 18322 23196 18328 23248
rect 18380 23236 18386 23248
rect 18693 23239 18751 23245
rect 18693 23236 18705 23239
rect 18380 23208 18705 23236
rect 18380 23196 18386 23208
rect 18693 23205 18705 23208
rect 18739 23236 18751 23239
rect 24394 23236 24400 23248
rect 18739 23208 19932 23236
rect 24355 23208 24400 23236
rect 18739 23205 18751 23208
rect 18693 23199 18751 23205
rect 16850 23168 16856 23180
rect 14835 23140 16856 23168
rect 16850 23128 16856 23140
rect 16908 23128 16914 23180
rect 19518 23128 19524 23180
rect 19576 23168 19582 23180
rect 19613 23171 19671 23177
rect 19613 23168 19625 23171
rect 19576 23140 19625 23168
rect 19576 23128 19582 23140
rect 19613 23137 19625 23140
rect 19659 23137 19671 23171
rect 19613 23131 19671 23137
rect 19904 23112 19932 23208
rect 24394 23196 24400 23208
rect 24452 23236 24458 23248
rect 25038 23236 25044 23248
rect 24452 23208 25044 23236
rect 24452 23196 24458 23208
rect 25038 23196 25044 23208
rect 25096 23196 25102 23248
rect 21726 23177 21732 23180
rect 21720 23168 21732 23177
rect 21687 23140 21732 23168
rect 21720 23131 21732 23140
rect 21726 23128 21732 23131
rect 21784 23128 21790 23180
rect 9401 23103 9459 23109
rect 9401 23100 9413 23103
rect 8996 23072 9413 23100
rect 8996 23060 9002 23072
rect 9401 23069 9413 23072
rect 9447 23100 9459 23103
rect 10137 23103 10195 23109
rect 10137 23100 10149 23103
rect 9447 23072 10149 23100
rect 9447 23069 9459 23072
rect 9401 23063 9459 23069
rect 10137 23069 10149 23072
rect 10183 23069 10195 23103
rect 10137 23063 10195 23069
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 12986 23060 12992 23112
rect 13044 23100 13050 23112
rect 15378 23100 15384 23112
rect 13044 23072 15384 23100
rect 13044 23060 13050 23072
rect 15378 23060 15384 23072
rect 15436 23100 15442 23112
rect 15473 23103 15531 23109
rect 15473 23100 15485 23103
rect 15436 23072 15485 23100
rect 15436 23060 15442 23072
rect 15473 23069 15485 23072
rect 15519 23100 15531 23103
rect 16022 23100 16028 23112
rect 15519 23072 16028 23100
rect 15519 23069 15531 23072
rect 15473 23063 15531 23069
rect 16022 23060 16028 23072
rect 16080 23060 16086 23112
rect 19153 23103 19211 23109
rect 19153 23069 19165 23103
rect 19199 23100 19211 23103
rect 19702 23100 19708 23112
rect 19199 23072 19708 23100
rect 19199 23069 19211 23072
rect 19153 23063 19211 23069
rect 19702 23060 19708 23072
rect 19760 23060 19766 23112
rect 19886 23100 19892 23112
rect 19847 23072 19892 23100
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 21450 23100 21456 23112
rect 21411 23072 21456 23100
rect 21450 23060 21456 23072
rect 21508 23060 21514 23112
rect 24210 23060 24216 23112
rect 24268 23100 24274 23112
rect 24489 23103 24547 23109
rect 24489 23100 24501 23103
rect 24268 23072 24501 23100
rect 24268 23060 24274 23072
rect 24489 23069 24501 23072
rect 24535 23069 24547 23103
rect 24489 23063 24547 23069
rect 3694 23032 3700 23044
rect 1728 23004 2728 23032
rect 2884 23004 3700 23032
rect 1728 22992 1734 23004
rect 1946 22964 1952 22976
rect 1907 22936 1952 22964
rect 1946 22924 1952 22936
rect 2004 22924 2010 22976
rect 2314 22964 2320 22976
rect 2275 22936 2320 22964
rect 2314 22924 2320 22936
rect 2372 22924 2378 22976
rect 2409 22967 2467 22973
rect 2409 22933 2421 22967
rect 2455 22964 2467 22967
rect 2590 22964 2596 22976
rect 2455 22936 2596 22964
rect 2455 22933 2467 22936
rect 2409 22927 2467 22933
rect 2590 22924 2596 22936
rect 2648 22924 2654 22976
rect 2700 22964 2728 23004
rect 3694 22992 3700 23004
rect 3752 22992 3758 23044
rect 8018 23032 8024 23044
rect 7979 23004 8024 23032
rect 8018 22992 8024 23004
rect 8076 22992 8082 23044
rect 13538 23032 13544 23044
rect 13499 23004 13544 23032
rect 13538 22992 13544 23004
rect 13596 22992 13602 23044
rect 14277 23035 14335 23041
rect 14277 23001 14289 23035
rect 14323 23032 14335 23035
rect 14826 23032 14832 23044
rect 14323 23004 14832 23032
rect 14323 23001 14335 23004
rect 14277 22995 14335 23001
rect 14826 22992 14832 23004
rect 14884 22992 14890 23044
rect 17402 23032 17408 23044
rect 17363 23004 17408 23032
rect 17402 22992 17408 23004
rect 17460 22992 17466 23044
rect 18966 22992 18972 23044
rect 19024 23032 19030 23044
rect 19426 23032 19432 23044
rect 19024 23004 19432 23032
rect 19024 22992 19030 23004
rect 19426 22992 19432 23004
rect 19484 23032 19490 23044
rect 20257 23035 20315 23041
rect 20257 23032 20269 23035
rect 19484 23004 20269 23032
rect 19484 22992 19490 23004
rect 20257 23001 20269 23004
rect 20303 23001 20315 23035
rect 20257 22995 20315 23001
rect 4249 22967 4307 22973
rect 4249 22964 4261 22967
rect 2700 22936 4261 22964
rect 4249 22933 4261 22936
rect 4295 22964 4307 22967
rect 4522 22964 4528 22976
rect 4295 22936 4528 22964
rect 4295 22933 4307 22936
rect 4249 22927 4307 22933
rect 4522 22924 4528 22936
rect 4580 22924 4586 22976
rect 6273 22967 6331 22973
rect 6273 22933 6285 22967
rect 6319 22964 6331 22967
rect 6362 22964 6368 22976
rect 6319 22936 6368 22964
rect 6319 22933 6331 22936
rect 6273 22927 6331 22933
rect 6362 22924 6368 22936
rect 6420 22964 6426 22976
rect 7098 22964 7104 22976
rect 6420 22936 7104 22964
rect 6420 22924 6426 22936
rect 7098 22924 7104 22936
rect 7156 22924 7162 22976
rect 13814 22964 13820 22976
rect 13775 22936 13820 22964
rect 13814 22924 13820 22936
rect 13872 22964 13878 22976
rect 13998 22964 14004 22976
rect 13872 22936 14004 22964
rect 13872 22924 13878 22936
rect 13998 22924 14004 22936
rect 14056 22924 14062 22976
rect 14642 22964 14648 22976
rect 14603 22936 14648 22964
rect 14642 22924 14648 22936
rect 14700 22924 14706 22976
rect 15933 22967 15991 22973
rect 15933 22933 15945 22967
rect 15979 22964 15991 22967
rect 16298 22964 16304 22976
rect 15979 22936 16304 22964
rect 15979 22933 15991 22936
rect 15933 22927 15991 22933
rect 16298 22924 16304 22936
rect 16356 22964 16362 22976
rect 17420 22964 17448 22992
rect 19242 22964 19248 22976
rect 16356 22936 17448 22964
rect 19203 22936 19248 22964
rect 16356 22924 16362 22936
rect 19242 22924 19248 22936
rect 19300 22924 19306 22976
rect 20714 22964 20720 22976
rect 20675 22936 20720 22964
rect 20714 22924 20720 22936
rect 20772 22924 20778 22976
rect 22554 22924 22560 22976
rect 22612 22964 22618 22976
rect 22833 22967 22891 22973
rect 22833 22964 22845 22967
rect 22612 22936 22845 22964
rect 22612 22924 22618 22936
rect 22833 22933 22845 22936
rect 22879 22933 22891 22967
rect 22833 22927 22891 22933
rect 23014 22924 23020 22976
rect 23072 22964 23078 22976
rect 23661 22967 23719 22973
rect 23661 22964 23673 22967
rect 23072 22936 23673 22964
rect 23072 22924 23078 22936
rect 23661 22933 23673 22936
rect 23707 22964 23719 22967
rect 24118 22964 24124 22976
rect 23707 22936 24124 22964
rect 23707 22933 23719 22936
rect 23661 22927 23719 22933
rect 24118 22924 24124 22936
rect 24176 22924 24182 22976
rect 25130 22924 25136 22976
rect 25188 22964 25194 22976
rect 25317 22967 25375 22973
rect 25317 22964 25329 22967
rect 25188 22936 25329 22964
rect 25188 22924 25194 22936
rect 25317 22933 25329 22936
rect 25363 22933 25375 22967
rect 25317 22927 25375 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2869 22763 2927 22769
rect 2869 22729 2881 22763
rect 2915 22760 2927 22763
rect 3510 22760 3516 22772
rect 2915 22732 3516 22760
rect 2915 22729 2927 22732
rect 2869 22723 2927 22729
rect 2314 22584 2320 22636
rect 2372 22624 2378 22636
rect 2409 22627 2467 22633
rect 2409 22624 2421 22627
rect 2372 22596 2421 22624
rect 2372 22584 2378 22596
rect 2409 22593 2421 22596
rect 2455 22624 2467 22627
rect 2884 22624 2912 22723
rect 3510 22720 3516 22732
rect 3568 22720 3574 22772
rect 4982 22760 4988 22772
rect 4943 22732 4988 22760
rect 4982 22720 4988 22732
rect 5040 22720 5046 22772
rect 5169 22763 5227 22769
rect 5169 22729 5181 22763
rect 5215 22760 5227 22763
rect 5534 22760 5540 22772
rect 5215 22732 5540 22760
rect 5215 22729 5227 22732
rect 5169 22723 5227 22729
rect 4433 22695 4491 22701
rect 4433 22661 4445 22695
rect 4479 22692 4491 22695
rect 4614 22692 4620 22704
rect 4479 22664 4620 22692
rect 4479 22661 4491 22664
rect 4433 22655 4491 22661
rect 4614 22652 4620 22664
rect 4672 22652 4678 22704
rect 3878 22624 3884 22636
rect 2455 22596 2912 22624
rect 3839 22596 3884 22624
rect 2455 22593 2467 22596
rect 2409 22587 2467 22593
rect 3878 22584 3884 22596
rect 3936 22584 3942 22636
rect 4798 22584 4804 22636
rect 4856 22624 4862 22636
rect 4982 22624 4988 22636
rect 4856 22596 4988 22624
rect 4856 22584 4862 22596
rect 4982 22584 4988 22596
rect 5040 22584 5046 22636
rect 1946 22516 1952 22568
rect 2004 22556 2010 22568
rect 2225 22559 2283 22565
rect 2225 22556 2237 22559
rect 2004 22528 2237 22556
rect 2004 22516 2010 22528
rect 2225 22525 2237 22528
rect 2271 22525 2283 22559
rect 2225 22519 2283 22525
rect 3237 22559 3295 22565
rect 3237 22525 3249 22559
rect 3283 22556 3295 22559
rect 3896 22556 3924 22584
rect 3283 22528 3924 22556
rect 3283 22525 3295 22528
rect 3237 22519 3295 22525
rect 2133 22491 2191 22497
rect 2133 22488 2145 22491
rect 1596 22460 2145 22488
rect 1394 22380 1400 22432
rect 1452 22420 1458 22432
rect 1596 22429 1624 22460
rect 2133 22457 2145 22460
rect 2179 22457 2191 22491
rect 2133 22451 2191 22457
rect 2590 22448 2596 22500
rect 2648 22488 2654 22500
rect 3789 22491 3847 22497
rect 2648 22460 3740 22488
rect 2648 22448 2654 22460
rect 1581 22423 1639 22429
rect 1581 22420 1593 22423
rect 1452 22392 1593 22420
rect 1452 22380 1458 22392
rect 1581 22389 1593 22392
rect 1627 22389 1639 22423
rect 1762 22420 1768 22432
rect 1723 22392 1768 22420
rect 1581 22383 1639 22389
rect 1762 22380 1768 22392
rect 1820 22380 1826 22432
rect 2498 22380 2504 22432
rect 2556 22420 2562 22432
rect 3712 22429 3740 22460
rect 3789 22457 3801 22491
rect 3835 22488 3847 22491
rect 5184 22488 5212 22723
rect 5534 22720 5540 22732
rect 5592 22720 5598 22772
rect 7466 22760 7472 22772
rect 7427 22732 7472 22760
rect 7466 22720 7472 22732
rect 7524 22720 7530 22772
rect 7929 22763 7987 22769
rect 7929 22729 7941 22763
rect 7975 22760 7987 22763
rect 8754 22760 8760 22772
rect 7975 22732 8760 22760
rect 7975 22729 7987 22732
rect 7929 22723 7987 22729
rect 8754 22720 8760 22732
rect 8812 22720 8818 22772
rect 9122 22720 9128 22772
rect 9180 22760 9186 22772
rect 9401 22763 9459 22769
rect 9401 22760 9413 22763
rect 9180 22732 9413 22760
rect 9180 22720 9186 22732
rect 9401 22729 9413 22732
rect 9447 22729 9459 22763
rect 11514 22760 11520 22772
rect 11475 22732 11520 22760
rect 9401 22723 9459 22729
rect 11514 22720 11520 22732
rect 11572 22720 11578 22772
rect 13081 22763 13139 22769
rect 13081 22729 13093 22763
rect 13127 22760 13139 22763
rect 14642 22760 14648 22772
rect 13127 22732 14648 22760
rect 13127 22729 13139 22732
rect 13081 22723 13139 22729
rect 14642 22720 14648 22732
rect 14700 22720 14706 22772
rect 15286 22760 15292 22772
rect 15247 22732 15292 22760
rect 15286 22720 15292 22732
rect 15344 22720 15350 22772
rect 16022 22760 16028 22772
rect 15983 22732 16028 22760
rect 16022 22720 16028 22732
rect 16080 22720 16086 22772
rect 17494 22720 17500 22772
rect 17552 22760 17558 22772
rect 17773 22763 17831 22769
rect 17773 22760 17785 22763
rect 17552 22732 17785 22760
rect 17552 22720 17558 22732
rect 17773 22729 17785 22732
rect 17819 22729 17831 22763
rect 18506 22760 18512 22772
rect 18467 22732 18512 22760
rect 17773 22723 17831 22729
rect 6822 22692 6828 22704
rect 5828 22664 6828 22692
rect 5350 22584 5356 22636
rect 5408 22624 5414 22636
rect 5828 22633 5856 22664
rect 6822 22652 6828 22664
rect 6880 22652 6886 22704
rect 5813 22627 5871 22633
rect 5813 22624 5825 22627
rect 5408 22596 5825 22624
rect 5408 22584 5414 22596
rect 5813 22593 5825 22596
rect 5859 22593 5871 22627
rect 7484 22624 7512 22720
rect 9674 22652 9680 22704
rect 9732 22692 9738 22704
rect 10042 22692 10048 22704
rect 9732 22664 10048 22692
rect 9732 22652 9738 22664
rect 10042 22652 10048 22664
rect 10100 22692 10106 22704
rect 10505 22695 10563 22701
rect 10505 22692 10517 22695
rect 10100 22664 10517 22692
rect 10100 22652 10106 22664
rect 10505 22661 10517 22664
rect 10551 22661 10563 22695
rect 10505 22655 10563 22661
rect 12986 22652 12992 22704
rect 13044 22692 13050 22704
rect 13725 22695 13783 22701
rect 13725 22692 13737 22695
rect 13044 22664 13737 22692
rect 13044 22652 13050 22664
rect 13725 22661 13737 22664
rect 13771 22692 13783 22695
rect 13771 22664 13952 22692
rect 13771 22661 13783 22664
rect 13725 22655 13783 22661
rect 8021 22627 8079 22633
rect 8021 22624 8033 22627
rect 7484 22596 8033 22624
rect 5813 22587 5871 22593
rect 8021 22593 8033 22596
rect 8067 22593 8079 22627
rect 8021 22587 8079 22593
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 10962 22624 10968 22636
rect 9999 22596 10968 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 10962 22584 10968 22596
rect 11020 22584 11026 22636
rect 13924 22633 13952 22664
rect 11057 22627 11115 22633
rect 11057 22593 11069 22627
rect 11103 22593 11115 22627
rect 11057 22587 11115 22593
rect 13909 22627 13967 22633
rect 13909 22593 13921 22627
rect 13955 22593 13967 22627
rect 16942 22624 16948 22636
rect 16903 22596 16948 22624
rect 13909 22587 13967 22593
rect 5629 22559 5687 22565
rect 5629 22525 5641 22559
rect 5675 22556 5687 22559
rect 5994 22556 6000 22568
rect 5675 22528 6000 22556
rect 5675 22525 5687 22528
rect 5629 22519 5687 22525
rect 5994 22516 6000 22528
rect 6052 22556 6058 22568
rect 6181 22559 6239 22565
rect 6181 22556 6193 22559
rect 6052 22528 6193 22556
rect 6052 22516 6058 22528
rect 6181 22525 6193 22528
rect 6227 22525 6239 22559
rect 6825 22559 6883 22565
rect 6825 22556 6837 22559
rect 6181 22519 6239 22525
rect 6564 22528 6837 22556
rect 3835 22460 5212 22488
rect 3835 22457 3847 22460
rect 3789 22451 3847 22457
rect 6564 22432 6592 22528
rect 6825 22525 6837 22528
rect 6871 22525 6883 22559
rect 6825 22519 6883 22525
rect 9858 22516 9864 22568
rect 9916 22556 9922 22568
rect 10778 22556 10784 22568
rect 9916 22528 10784 22556
rect 9916 22516 9922 22528
rect 10778 22516 10784 22528
rect 10836 22556 10842 22568
rect 11072 22556 11100 22587
rect 16942 22584 16948 22596
rect 17000 22584 17006 22636
rect 10836 22528 11100 22556
rect 10836 22516 10842 22528
rect 11790 22516 11796 22568
rect 11848 22556 11854 22568
rect 11977 22559 12035 22565
rect 11977 22556 11989 22559
rect 11848 22528 11989 22556
rect 11848 22516 11854 22528
rect 11977 22525 11989 22528
rect 12023 22556 12035 22559
rect 12710 22556 12716 22568
rect 12023 22528 12716 22556
rect 12023 22525 12035 22528
rect 11977 22519 12035 22525
rect 12710 22516 12716 22528
rect 12768 22516 12774 22568
rect 12897 22559 12955 22565
rect 12897 22525 12909 22559
rect 12943 22556 12955 22559
rect 13814 22556 13820 22568
rect 12943 22528 13820 22556
rect 12943 22525 12955 22528
rect 12897 22519 12955 22525
rect 13814 22516 13820 22528
rect 13872 22516 13878 22568
rect 17788 22556 17816 22723
rect 18506 22720 18512 22732
rect 18564 22720 18570 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 20806 22760 20812 22772
rect 19484 22732 20812 22760
rect 19484 22720 19490 22732
rect 20806 22720 20812 22732
rect 20864 22720 20870 22772
rect 20901 22763 20959 22769
rect 20901 22729 20913 22763
rect 20947 22760 20959 22763
rect 20990 22760 20996 22772
rect 20947 22732 20996 22760
rect 20947 22729 20959 22732
rect 20901 22723 20959 22729
rect 20990 22720 20996 22732
rect 21048 22760 21054 22772
rect 22186 22760 22192 22772
rect 21048 22732 22192 22760
rect 21048 22720 21054 22732
rect 22186 22720 22192 22732
rect 22244 22720 22250 22772
rect 24118 22720 24124 22772
rect 24176 22760 24182 22772
rect 24670 22760 24676 22772
rect 24176 22732 24676 22760
rect 24176 22720 24182 22732
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 25038 22760 25044 22772
rect 24999 22732 25044 22760
rect 25038 22720 25044 22732
rect 25096 22720 25102 22772
rect 25409 22763 25467 22769
rect 25409 22729 25421 22763
rect 25455 22760 25467 22763
rect 26142 22760 26148 22772
rect 25455 22732 26148 22760
rect 25455 22729 25467 22732
rect 25409 22723 25467 22729
rect 26142 22720 26148 22732
rect 26200 22720 26206 22772
rect 21818 22692 21824 22704
rect 21779 22664 21824 22692
rect 21818 22652 21824 22664
rect 21876 22692 21882 22704
rect 21876 22664 21956 22692
rect 21876 22652 21882 22664
rect 21928 22624 21956 22664
rect 22094 22652 22100 22704
rect 22152 22692 22158 22704
rect 22462 22692 22468 22704
rect 22152 22664 22468 22692
rect 22152 22652 22158 22664
rect 22462 22652 22468 22664
rect 22520 22652 22526 22704
rect 22554 22624 22560 22636
rect 21928 22596 22560 22624
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 24210 22624 24216 22636
rect 24171 22596 24216 22624
rect 24210 22584 24216 22596
rect 24268 22624 24274 22636
rect 24673 22627 24731 22633
rect 24673 22624 24685 22627
rect 24268 22596 24685 22624
rect 24268 22584 24274 22596
rect 24673 22593 24685 22596
rect 24719 22593 24731 22627
rect 24673 22587 24731 22593
rect 18325 22559 18383 22565
rect 18325 22556 18337 22559
rect 17788 22528 18337 22556
rect 18325 22525 18337 22528
rect 18371 22525 18383 22559
rect 19521 22559 19579 22565
rect 19521 22556 19533 22559
rect 18325 22519 18383 22525
rect 18892 22528 19533 22556
rect 8288 22491 8346 22497
rect 8288 22457 8300 22491
rect 8334 22488 8346 22491
rect 8386 22488 8392 22500
rect 8334 22460 8392 22488
rect 8334 22457 8346 22460
rect 8288 22451 8346 22457
rect 8386 22448 8392 22460
rect 8444 22448 8450 22500
rect 10873 22491 10931 22497
rect 10873 22488 10885 22491
rect 10336 22460 10885 22488
rect 3329 22423 3387 22429
rect 3329 22420 3341 22423
rect 2556 22392 3341 22420
rect 2556 22380 2562 22392
rect 3329 22389 3341 22392
rect 3375 22389 3387 22423
rect 3329 22383 3387 22389
rect 3697 22423 3755 22429
rect 3697 22389 3709 22423
rect 3743 22420 3755 22423
rect 4706 22420 4712 22432
rect 3743 22392 4712 22420
rect 3743 22389 3755 22392
rect 3697 22383 3755 22389
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 5534 22420 5540 22432
rect 5495 22392 5540 22420
rect 5534 22380 5540 22392
rect 5592 22380 5598 22432
rect 6546 22420 6552 22432
rect 6507 22392 6552 22420
rect 6546 22380 6552 22392
rect 6604 22380 6610 22432
rect 7009 22423 7067 22429
rect 7009 22389 7021 22423
rect 7055 22420 7067 22423
rect 7098 22420 7104 22432
rect 7055 22392 7104 22420
rect 7055 22389 7067 22392
rect 7009 22383 7067 22389
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 10134 22380 10140 22432
rect 10192 22420 10198 22432
rect 10336 22429 10364 22460
rect 10873 22457 10885 22460
rect 10919 22457 10931 22491
rect 10873 22451 10931 22457
rect 11146 22448 11152 22500
rect 11204 22488 11210 22500
rect 14182 22497 14188 22500
rect 13357 22491 13415 22497
rect 13357 22488 13369 22491
rect 11204 22460 13369 22488
rect 11204 22448 11210 22460
rect 13357 22457 13369 22460
rect 13403 22457 13415 22491
rect 14176 22488 14188 22497
rect 14143 22460 14188 22488
rect 13357 22451 13415 22457
rect 14176 22451 14188 22460
rect 14182 22448 14188 22451
rect 14240 22448 14246 22500
rect 16482 22448 16488 22500
rect 16540 22488 16546 22500
rect 16540 22460 16896 22488
rect 16540 22448 16546 22460
rect 10321 22423 10379 22429
rect 10321 22420 10333 22423
rect 10192 22392 10333 22420
rect 10192 22380 10198 22392
rect 10321 22389 10333 22392
rect 10367 22389 10379 22423
rect 12618 22420 12624 22432
rect 12579 22392 12624 22420
rect 10321 22383 10379 22389
rect 12618 22380 12624 22392
rect 12676 22380 12682 22432
rect 16390 22420 16396 22432
rect 16351 22392 16396 22420
rect 16390 22380 16396 22392
rect 16448 22380 16454 22432
rect 16758 22420 16764 22432
rect 16719 22392 16764 22420
rect 16758 22380 16764 22392
rect 16816 22380 16822 22432
rect 16868 22429 16896 22460
rect 16853 22423 16911 22429
rect 16853 22389 16865 22423
rect 16899 22420 16911 22423
rect 17405 22423 17463 22429
rect 17405 22420 17417 22423
rect 16899 22392 17417 22420
rect 16899 22389 16911 22392
rect 16853 22383 16911 22389
rect 17405 22389 17417 22392
rect 17451 22389 17463 22423
rect 17405 22383 17463 22389
rect 18322 22380 18328 22432
rect 18380 22420 18386 22432
rect 18892 22429 18920 22528
rect 19521 22525 19533 22528
rect 19567 22556 19579 22559
rect 21450 22556 21456 22568
rect 19567 22528 21456 22556
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 21450 22516 21456 22528
rect 21508 22516 21514 22568
rect 22462 22556 22468 22568
rect 22423 22528 22468 22556
rect 22462 22516 22468 22528
rect 22520 22516 22526 22568
rect 23474 22516 23480 22568
rect 23532 22556 23538 22568
rect 24029 22559 24087 22565
rect 24029 22556 24041 22559
rect 23532 22528 24041 22556
rect 23532 22516 23538 22528
rect 24029 22525 24041 22528
rect 24075 22556 24087 22559
rect 25130 22556 25136 22568
rect 24075 22528 25136 22556
rect 24075 22525 24087 22528
rect 24029 22519 24087 22525
rect 25130 22516 25136 22528
rect 25188 22516 25194 22568
rect 25225 22559 25283 22565
rect 25225 22525 25237 22559
rect 25271 22556 25283 22559
rect 25314 22556 25320 22568
rect 25271 22528 25320 22556
rect 25271 22525 25283 22528
rect 25225 22519 25283 22525
rect 25314 22516 25320 22528
rect 25372 22516 25378 22568
rect 19788 22491 19846 22497
rect 19788 22457 19800 22491
rect 19834 22488 19846 22491
rect 19978 22488 19984 22500
rect 19834 22460 19984 22488
rect 19834 22457 19846 22460
rect 19788 22451 19846 22457
rect 19978 22448 19984 22460
rect 20036 22488 20042 22500
rect 20346 22488 20352 22500
rect 20036 22460 20352 22488
rect 20036 22448 20042 22460
rect 20346 22448 20352 22460
rect 20404 22448 20410 22500
rect 23750 22448 23756 22500
rect 23808 22488 23814 22500
rect 24121 22491 24179 22497
rect 24121 22488 24133 22491
rect 23808 22460 24133 22488
rect 23808 22448 23814 22460
rect 24121 22457 24133 22460
rect 24167 22488 24179 22491
rect 25777 22491 25835 22497
rect 25777 22488 25789 22491
rect 24167 22460 25789 22488
rect 24167 22457 24179 22460
rect 24121 22451 24179 22457
rect 25777 22457 25789 22460
rect 25823 22457 25835 22491
rect 25777 22451 25835 22457
rect 18877 22423 18935 22429
rect 18877 22420 18889 22423
rect 18380 22392 18889 22420
rect 18380 22380 18386 22392
rect 18877 22389 18889 22392
rect 18923 22389 18935 22423
rect 18877 22383 18935 22389
rect 19337 22423 19395 22429
rect 19337 22389 19349 22423
rect 19383 22420 19395 22423
rect 19518 22420 19524 22432
rect 19383 22392 19524 22420
rect 19383 22389 19395 22392
rect 19337 22383 19395 22389
rect 19518 22380 19524 22392
rect 19576 22420 19582 22432
rect 20438 22420 20444 22432
rect 19576 22392 20444 22420
rect 19576 22380 19582 22392
rect 20438 22380 20444 22392
rect 20496 22380 20502 22432
rect 21818 22380 21824 22432
rect 21876 22420 21882 22432
rect 22005 22423 22063 22429
rect 22005 22420 22017 22423
rect 21876 22392 22017 22420
rect 21876 22380 21882 22392
rect 22005 22389 22017 22392
rect 22051 22389 22063 22423
rect 22370 22420 22376 22432
rect 22331 22392 22376 22420
rect 22005 22383 22063 22389
rect 22370 22380 22376 22392
rect 22428 22380 22434 22432
rect 22922 22380 22928 22432
rect 22980 22420 22986 22432
rect 23290 22420 23296 22432
rect 22980 22392 23296 22420
rect 22980 22380 22986 22392
rect 23290 22380 23296 22392
rect 23348 22380 23354 22432
rect 23474 22380 23480 22432
rect 23532 22420 23538 22432
rect 23661 22423 23719 22429
rect 23661 22420 23673 22423
rect 23532 22392 23673 22420
rect 23532 22380 23538 22392
rect 23661 22389 23673 22392
rect 23707 22389 23719 22423
rect 23661 22383 23719 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1210 22176 1216 22228
rect 1268 22216 1274 22228
rect 1949 22219 2007 22225
rect 1949 22216 1961 22219
rect 1268 22188 1961 22216
rect 1268 22176 1274 22188
rect 1949 22185 1961 22188
rect 1995 22216 2007 22219
rect 2590 22216 2596 22228
rect 1995 22188 2596 22216
rect 1995 22185 2007 22188
rect 1949 22179 2007 22185
rect 2590 22176 2596 22188
rect 2648 22176 2654 22228
rect 3050 22216 3056 22228
rect 3011 22188 3056 22216
rect 3050 22176 3056 22188
rect 3108 22216 3114 22228
rect 3881 22219 3939 22225
rect 3881 22216 3893 22219
rect 3108 22188 3893 22216
rect 3108 22176 3114 22188
rect 3881 22185 3893 22188
rect 3927 22185 3939 22219
rect 3881 22179 3939 22185
rect 5534 22176 5540 22228
rect 5592 22216 5598 22228
rect 5905 22219 5963 22225
rect 5905 22216 5917 22219
rect 5592 22188 5917 22216
rect 5592 22176 5598 22188
rect 5905 22185 5917 22188
rect 5951 22185 5963 22219
rect 8662 22216 8668 22228
rect 8623 22188 8668 22216
rect 5905 22179 5963 22185
rect 8662 22176 8668 22188
rect 8720 22176 8726 22228
rect 9398 22216 9404 22228
rect 9359 22188 9404 22216
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 10042 22176 10048 22228
rect 10100 22216 10106 22228
rect 10321 22219 10379 22225
rect 10321 22216 10333 22219
rect 10100 22188 10333 22216
rect 10100 22176 10106 22188
rect 1670 22108 1676 22160
rect 1728 22148 1734 22160
rect 2041 22151 2099 22157
rect 2041 22148 2053 22151
rect 1728 22120 2053 22148
rect 1728 22108 1734 22120
rect 2041 22117 2053 22120
rect 2087 22117 2099 22151
rect 2041 22111 2099 22117
rect 4433 22151 4491 22157
rect 4433 22117 4445 22151
rect 4479 22148 4491 22151
rect 4614 22148 4620 22160
rect 4479 22120 4620 22148
rect 4479 22117 4491 22120
rect 4433 22111 4491 22117
rect 4614 22108 4620 22120
rect 4672 22108 4678 22160
rect 5442 22080 5448 22092
rect 4724 22052 5448 22080
rect 2222 22012 2228 22024
rect 2135 21984 2228 22012
rect 2222 21972 2228 21984
rect 2280 22012 2286 22024
rect 3329 22015 3387 22021
rect 3329 22012 3341 22015
rect 2280 21984 3341 22012
rect 2280 21972 2286 21984
rect 3329 21981 3341 21984
rect 3375 21981 3387 22015
rect 4522 22012 4528 22024
rect 4483 21984 4528 22012
rect 3329 21975 3387 21981
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 4724 22021 4752 22052
rect 5442 22040 5448 22052
rect 5500 22080 5506 22092
rect 5537 22083 5595 22089
rect 5537 22080 5549 22083
rect 5500 22052 5549 22080
rect 5500 22040 5506 22052
rect 5537 22049 5549 22052
rect 5583 22049 5595 22083
rect 5537 22043 5595 22049
rect 6362 22040 6368 22092
rect 6420 22080 6426 22092
rect 6529 22083 6587 22089
rect 6529 22080 6541 22083
rect 6420 22052 6541 22080
rect 6420 22040 6426 22052
rect 6529 22049 6541 22052
rect 6575 22049 6587 22083
rect 10152 22080 10180 22188
rect 10321 22185 10333 22188
rect 10367 22185 10379 22219
rect 10321 22179 10379 22185
rect 10778 22176 10784 22228
rect 10836 22216 10842 22228
rect 10873 22219 10931 22225
rect 10873 22216 10885 22219
rect 10836 22188 10885 22216
rect 10836 22176 10842 22188
rect 10873 22185 10885 22188
rect 10919 22185 10931 22219
rect 10873 22179 10931 22185
rect 12434 22176 12440 22228
rect 12492 22216 12498 22228
rect 16298 22216 16304 22228
rect 12492 22188 14596 22216
rect 16259 22188 16304 22216
rect 12492 22176 12498 22188
rect 10229 22151 10287 22157
rect 10229 22117 10241 22151
rect 10275 22148 10287 22151
rect 10686 22148 10692 22160
rect 10275 22120 10692 22148
rect 10275 22117 10287 22120
rect 10229 22111 10287 22117
rect 10686 22108 10692 22120
rect 10744 22108 10750 22160
rect 11514 22108 11520 22160
rect 11572 22108 11578 22160
rect 11692 22151 11750 22157
rect 11692 22117 11704 22151
rect 11738 22148 11750 22151
rect 12250 22148 12256 22160
rect 11738 22120 12256 22148
rect 11738 22117 11750 22120
rect 11692 22111 11750 22117
rect 12250 22108 12256 22120
rect 12308 22148 12314 22160
rect 12894 22148 12900 22160
rect 12308 22120 12900 22148
rect 12308 22108 12314 22120
rect 12894 22108 12900 22120
rect 12952 22108 12958 22160
rect 14001 22151 14059 22157
rect 14001 22117 14013 22151
rect 14047 22148 14059 22151
rect 14182 22148 14188 22160
rect 14047 22120 14188 22148
rect 14047 22117 14059 22120
rect 14001 22111 14059 22117
rect 14182 22108 14188 22120
rect 14240 22108 14246 22160
rect 14458 22108 14464 22160
rect 14516 22108 14522 22160
rect 14568 22148 14596 22188
rect 16298 22176 16304 22188
rect 16356 22176 16362 22228
rect 18690 22216 18696 22228
rect 16408 22188 18696 22216
rect 16408 22148 16436 22188
rect 18690 22176 18696 22188
rect 18748 22176 18754 22228
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 21913 22219 21971 22225
rect 21913 22216 21925 22219
rect 20772 22188 21925 22216
rect 20772 22176 20778 22188
rect 21913 22185 21925 22188
rect 21959 22216 21971 22219
rect 22370 22216 22376 22228
rect 21959 22188 22376 22216
rect 21959 22185 21971 22188
rect 21913 22179 21971 22185
rect 22370 22176 22376 22188
rect 22428 22176 22434 22228
rect 22462 22176 22468 22228
rect 22520 22216 22526 22228
rect 22925 22219 22983 22225
rect 22925 22216 22937 22219
rect 22520 22188 22937 22216
rect 22520 22176 22526 22188
rect 22925 22185 22937 22188
rect 22971 22185 22983 22219
rect 22925 22179 22983 22185
rect 17126 22148 17132 22160
rect 14568 22120 16436 22148
rect 17087 22120 17132 22148
rect 17126 22108 17132 22120
rect 17184 22108 17190 22160
rect 20806 22108 20812 22160
rect 20864 22148 20870 22160
rect 20901 22151 20959 22157
rect 20901 22148 20913 22151
rect 20864 22120 20913 22148
rect 20864 22108 20870 22120
rect 20901 22117 20913 22120
rect 20947 22117 20959 22151
rect 23290 22148 23296 22160
rect 20901 22111 20959 22117
rect 21008 22120 23296 22148
rect 10318 22080 10324 22092
rect 10152 22052 10324 22080
rect 6529 22043 6587 22049
rect 10318 22040 10324 22052
rect 10376 22040 10382 22092
rect 11330 22080 11336 22092
rect 11291 22052 11336 22080
rect 11330 22040 11336 22052
rect 11388 22040 11394 22092
rect 4709 22015 4767 22021
rect 4709 21981 4721 22015
rect 4755 21981 4767 22015
rect 4709 21975 4767 21981
rect 6086 21972 6092 22024
rect 6144 22012 6150 22024
rect 6273 22015 6331 22021
rect 6273 22012 6285 22015
rect 6144 21984 6285 22012
rect 6144 21972 6150 21984
rect 6273 21981 6285 21984
rect 6319 21981 6331 22015
rect 6273 21975 6331 21981
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 22012 9183 22015
rect 9582 22012 9588 22024
rect 9171 21984 9588 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 9582 21972 9588 21984
rect 9640 21972 9646 22024
rect 10502 22012 10508 22024
rect 10463 21984 10508 22012
rect 10502 21972 10508 21984
rect 10560 21972 10566 22024
rect 11425 22015 11483 22021
rect 11425 21981 11437 22015
rect 11471 22012 11483 22015
rect 11532 22012 11560 22108
rect 14093 22083 14151 22089
rect 14093 22049 14105 22083
rect 14139 22080 14151 22083
rect 14139 22052 14412 22080
rect 14139 22049 14151 22052
rect 14093 22043 14151 22049
rect 11471 21984 11560 22012
rect 11471 21981 11483 21984
rect 11425 21975 11483 21981
rect 3050 21904 3056 21956
rect 3108 21944 3114 21956
rect 3881 21947 3939 21953
rect 3108 21916 3832 21944
rect 3108 21904 3114 21916
rect 1578 21876 1584 21888
rect 1539 21848 1584 21876
rect 1578 21836 1584 21848
rect 1636 21836 1642 21888
rect 1946 21836 1952 21888
rect 2004 21876 2010 21888
rect 2593 21879 2651 21885
rect 2593 21876 2605 21879
rect 2004 21848 2605 21876
rect 2004 21836 2010 21848
rect 2593 21845 2605 21848
rect 2639 21845 2651 21879
rect 2593 21839 2651 21845
rect 2866 21836 2872 21888
rect 2924 21876 2930 21888
rect 3418 21876 3424 21888
rect 2924 21848 3424 21876
rect 2924 21836 2930 21848
rect 3418 21836 3424 21848
rect 3476 21836 3482 21888
rect 3602 21836 3608 21888
rect 3660 21876 3666 21888
rect 3697 21879 3755 21885
rect 3697 21876 3709 21879
rect 3660 21848 3709 21876
rect 3660 21836 3666 21848
rect 3697 21845 3709 21848
rect 3743 21845 3755 21879
rect 3804 21876 3832 21916
rect 3881 21913 3893 21947
rect 3927 21944 3939 21947
rect 5169 21947 5227 21953
rect 5169 21944 5181 21947
rect 3927 21916 5181 21944
rect 3927 21913 3939 21916
rect 3881 21907 3939 21913
rect 5169 21913 5181 21916
rect 5215 21944 5227 21947
rect 5350 21944 5356 21956
rect 5215 21916 5356 21944
rect 5215 21913 5227 21916
rect 5169 21907 5227 21913
rect 5350 21904 5356 21916
rect 5408 21904 5414 21956
rect 9858 21944 9864 21956
rect 9819 21916 9864 21944
rect 9858 21904 9864 21916
rect 9916 21904 9922 21956
rect 14274 21944 14280 21956
rect 14235 21916 14280 21944
rect 14274 21904 14280 21916
rect 14332 21904 14338 21956
rect 14384 21944 14412 22052
rect 14476 22012 14504 22108
rect 15378 22040 15384 22092
rect 15436 22080 15442 22092
rect 15657 22083 15715 22089
rect 15657 22080 15669 22083
rect 15436 22052 15669 22080
rect 15436 22040 15442 22052
rect 15657 22049 15669 22052
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 17221 22083 17279 22089
rect 17221 22049 17233 22083
rect 17267 22080 17279 22083
rect 17310 22080 17316 22092
rect 17267 22052 17316 22080
rect 17267 22049 17279 22052
rect 17221 22043 17279 22049
rect 17310 22040 17316 22052
rect 17368 22040 17374 22092
rect 17862 22040 17868 22092
rect 17920 22080 17926 22092
rect 18581 22083 18639 22089
rect 18581 22080 18593 22083
rect 17920 22052 18593 22080
rect 17920 22040 17926 22052
rect 18581 22049 18593 22052
rect 18627 22049 18639 22083
rect 20346 22080 20352 22092
rect 20307 22052 20352 22080
rect 18581 22043 18639 22049
rect 20346 22040 20352 22052
rect 20404 22080 20410 22092
rect 21008 22080 21036 22120
rect 23290 22108 23296 22120
rect 23348 22108 23354 22160
rect 20404 22052 21036 22080
rect 22281 22083 22339 22089
rect 20404 22040 20410 22052
rect 22281 22049 22293 22083
rect 22327 22080 22339 22083
rect 22922 22080 22928 22092
rect 22327 22052 22928 22080
rect 22327 22049 22339 22052
rect 22281 22043 22339 22049
rect 22922 22040 22928 22052
rect 22980 22040 22986 22092
rect 23845 22083 23903 22089
rect 23845 22080 23857 22083
rect 23768 22052 23857 22080
rect 23768 22024 23796 22052
rect 23845 22049 23857 22052
rect 23891 22049 23903 22083
rect 24854 22080 24860 22092
rect 24815 22052 24860 22080
rect 23845 22043 23903 22049
rect 24854 22040 24860 22052
rect 24912 22040 24918 22092
rect 25038 22080 25044 22092
rect 24999 22052 25044 22080
rect 25038 22040 25044 22052
rect 25096 22040 25102 22092
rect 25314 22040 25320 22092
rect 25372 22080 25378 22092
rect 25593 22083 25651 22089
rect 25593 22080 25605 22083
rect 25372 22052 25605 22080
rect 25372 22040 25378 22052
rect 25593 22049 25605 22052
rect 25639 22049 25651 22083
rect 25593 22043 25651 22049
rect 14642 22012 14648 22024
rect 14476 21984 14648 22012
rect 14642 21972 14648 21984
rect 14700 21972 14706 22024
rect 17402 22012 17408 22024
rect 17363 21984 17408 22012
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 18322 22012 18328 22024
rect 18283 21984 18328 22012
rect 18322 21972 18328 21984
rect 18380 21972 18386 22024
rect 20717 22015 20775 22021
rect 20717 21981 20729 22015
rect 20763 22012 20775 22015
rect 21726 22012 21732 22024
rect 20763 21984 21732 22012
rect 20763 21981 20775 21984
rect 20717 21975 20775 21981
rect 21726 21972 21732 21984
rect 21784 21972 21790 22024
rect 22373 22015 22431 22021
rect 22373 21981 22385 22015
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22465 22015 22523 22021
rect 22465 21981 22477 22015
rect 22511 22012 22523 22015
rect 22511 21984 22683 22012
rect 22511 21981 22523 21984
rect 22465 21975 22523 21981
rect 14826 21944 14832 21956
rect 14384 21916 14832 21944
rect 14826 21904 14832 21916
rect 14884 21904 14890 21956
rect 15838 21944 15844 21956
rect 15799 21916 15844 21944
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 16758 21944 16764 21956
rect 16671 21916 16764 21944
rect 16758 21904 16764 21916
rect 16816 21944 16822 21956
rect 17773 21947 17831 21953
rect 17773 21944 17785 21947
rect 16816 21916 17785 21944
rect 16816 21904 16822 21916
rect 17773 21913 17785 21916
rect 17819 21913 17831 21947
rect 19702 21944 19708 21956
rect 19663 21916 19708 21944
rect 17773 21907 17831 21913
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 22388 21944 22416 21975
rect 22554 21944 22560 21956
rect 22388 21916 22560 21944
rect 22554 21904 22560 21916
rect 22612 21904 22618 21956
rect 4065 21879 4123 21885
rect 4065 21876 4077 21879
rect 3804 21848 4077 21876
rect 3697 21839 3755 21845
rect 4065 21845 4077 21848
rect 4111 21845 4123 21879
rect 7650 21876 7656 21888
rect 7611 21848 7656 21876
rect 4065 21839 4123 21845
rect 7650 21836 7656 21848
rect 7708 21836 7714 21888
rect 8297 21879 8355 21885
rect 8297 21845 8309 21879
rect 8343 21876 8355 21879
rect 8386 21876 8392 21888
rect 8343 21848 8392 21876
rect 8343 21845 8355 21848
rect 8297 21839 8355 21845
rect 8386 21836 8392 21848
rect 8444 21836 8450 21888
rect 11422 21836 11428 21888
rect 11480 21876 11486 21888
rect 12342 21876 12348 21888
rect 11480 21848 12348 21876
rect 11480 21836 11486 21848
rect 12342 21836 12348 21848
rect 12400 21876 12406 21888
rect 12805 21879 12863 21885
rect 12805 21876 12817 21879
rect 12400 21848 12817 21876
rect 12400 21836 12406 21848
rect 12805 21845 12817 21848
rect 12851 21845 12863 21879
rect 12805 21839 12863 21845
rect 12894 21836 12900 21888
rect 12952 21876 12958 21888
rect 13357 21879 13415 21885
rect 13357 21876 13369 21879
rect 12952 21848 13369 21876
rect 12952 21836 12958 21848
rect 13357 21845 13369 21848
rect 13403 21845 13415 21879
rect 14734 21876 14740 21888
rect 14695 21848 14740 21876
rect 13357 21839 13415 21845
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 15562 21876 15568 21888
rect 15523 21848 15568 21876
rect 15562 21836 15568 21848
rect 15620 21836 15626 21888
rect 16022 21836 16028 21888
rect 16080 21876 16086 21888
rect 16577 21879 16635 21885
rect 16577 21876 16589 21879
rect 16080 21848 16589 21876
rect 16080 21836 16086 21848
rect 16577 21845 16589 21848
rect 16623 21876 16635 21879
rect 16942 21876 16948 21888
rect 16623 21848 16948 21876
rect 16623 21845 16635 21848
rect 16577 21839 16635 21845
rect 16942 21836 16948 21848
rect 17000 21836 17006 21888
rect 18233 21879 18291 21885
rect 18233 21845 18245 21879
rect 18279 21876 18291 21879
rect 18598 21876 18604 21888
rect 18279 21848 18604 21876
rect 18279 21845 18291 21848
rect 18233 21839 18291 21845
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 21542 21876 21548 21888
rect 21503 21848 21548 21876
rect 21542 21836 21548 21848
rect 21600 21836 21606 21888
rect 21726 21836 21732 21888
rect 21784 21876 21790 21888
rect 22186 21876 22192 21888
rect 21784 21848 22192 21876
rect 21784 21836 21790 21848
rect 22186 21836 22192 21848
rect 22244 21876 22250 21888
rect 22655 21876 22683 21984
rect 23750 21972 23756 22024
rect 23808 21972 23814 22024
rect 23934 22012 23940 22024
rect 23895 21984 23940 22012
rect 23934 21972 23940 21984
rect 23992 21972 23998 22024
rect 24026 21972 24032 22024
rect 24084 22012 24090 22024
rect 24210 22012 24216 22024
rect 24084 21984 24216 22012
rect 24084 21972 24090 21984
rect 24210 21972 24216 21984
rect 24268 22012 24274 22024
rect 24489 22015 24547 22021
rect 24489 22012 24501 22015
rect 24268 21984 24501 22012
rect 24268 21972 24274 21984
rect 24489 21981 24501 21984
rect 24535 21981 24547 22015
rect 24489 21975 24547 21981
rect 22922 21904 22928 21956
rect 22980 21944 22986 21956
rect 23477 21947 23535 21953
rect 23477 21944 23489 21947
rect 22980 21916 23489 21944
rect 22980 21904 22986 21916
rect 23477 21913 23489 21916
rect 23523 21913 23535 21947
rect 23477 21907 23535 21913
rect 22244 21848 22683 21876
rect 22244 21836 22250 21848
rect 23198 21836 23204 21888
rect 23256 21876 23262 21888
rect 23385 21879 23443 21885
rect 23385 21876 23397 21879
rect 23256 21848 23397 21876
rect 23256 21836 23262 21848
rect 23385 21845 23397 21848
rect 23431 21876 23443 21879
rect 24210 21876 24216 21888
rect 23431 21848 24216 21876
rect 23431 21845 23443 21848
rect 23385 21839 23443 21845
rect 24210 21836 24216 21848
rect 24268 21836 24274 21888
rect 25222 21876 25228 21888
rect 25183 21848 25228 21876
rect 25222 21836 25228 21848
rect 25280 21836 25286 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 2038 21672 2044 21684
rect 1636 21644 2044 21672
rect 1636 21632 1642 21644
rect 2038 21632 2044 21644
rect 2096 21632 2102 21684
rect 2590 21672 2596 21684
rect 2551 21644 2596 21672
rect 2590 21632 2596 21644
rect 2648 21672 2654 21684
rect 2866 21672 2872 21684
rect 2648 21644 2872 21672
rect 2648 21632 2654 21644
rect 2866 21632 2872 21644
rect 2924 21632 2930 21684
rect 4709 21675 4767 21681
rect 4709 21641 4721 21675
rect 4755 21672 4767 21675
rect 5353 21675 5411 21681
rect 5353 21672 5365 21675
rect 4755 21644 5365 21672
rect 4755 21641 4767 21644
rect 4709 21635 4767 21641
rect 5353 21641 5365 21644
rect 5399 21672 5411 21675
rect 5442 21672 5448 21684
rect 5399 21644 5448 21672
rect 5399 21641 5411 21644
rect 5353 21635 5411 21641
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 5905 21675 5963 21681
rect 5905 21641 5917 21675
rect 5951 21672 5963 21675
rect 6362 21672 6368 21684
rect 5951 21644 6368 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 6362 21632 6368 21644
rect 6420 21632 6426 21684
rect 10318 21672 10324 21684
rect 10279 21644 10324 21672
rect 10318 21632 10324 21644
rect 10376 21632 10382 21684
rect 10686 21672 10692 21684
rect 10647 21644 10692 21672
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 11422 21632 11428 21684
rect 11480 21672 11486 21684
rect 11606 21672 11612 21684
rect 11480 21644 11612 21672
rect 11480 21632 11486 21644
rect 11606 21632 11612 21644
rect 11664 21672 11670 21684
rect 11793 21675 11851 21681
rect 11793 21672 11805 21675
rect 11664 21644 11805 21672
rect 11664 21632 11670 21644
rect 11793 21641 11805 21644
rect 11839 21641 11851 21675
rect 12250 21672 12256 21684
rect 12211 21644 12256 21672
rect 11793 21635 11851 21641
rect 10042 21564 10048 21616
rect 10100 21604 10106 21616
rect 10502 21604 10508 21616
rect 10100 21576 10508 21604
rect 10100 21564 10106 21576
rect 10502 21564 10508 21576
rect 10560 21604 10566 21616
rect 11808 21604 11836 21635
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 14182 21632 14188 21684
rect 14240 21672 14246 21684
rect 14645 21675 14703 21681
rect 14645 21672 14657 21675
rect 14240 21644 14657 21672
rect 14240 21632 14246 21644
rect 14645 21641 14657 21644
rect 14691 21641 14703 21675
rect 14645 21635 14703 21641
rect 16393 21675 16451 21681
rect 16393 21641 16405 21675
rect 16439 21672 16451 21675
rect 16482 21672 16488 21684
rect 16439 21644 16488 21672
rect 16439 21641 16451 21644
rect 16393 21635 16451 21641
rect 16482 21632 16488 21644
rect 16540 21632 16546 21684
rect 17862 21672 17868 21684
rect 17823 21644 17868 21672
rect 17862 21632 17868 21644
rect 17920 21632 17926 21684
rect 22278 21632 22284 21684
rect 22336 21672 22342 21684
rect 22649 21675 22707 21681
rect 22649 21672 22661 21675
rect 22336 21644 22661 21672
rect 22336 21632 22342 21644
rect 22649 21641 22661 21644
rect 22695 21672 22707 21675
rect 24026 21672 24032 21684
rect 22695 21644 24032 21672
rect 22695 21641 22707 21644
rect 22649 21635 22707 21641
rect 24026 21632 24032 21644
rect 24084 21632 24090 21684
rect 25590 21672 25596 21684
rect 25551 21644 25596 21672
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 13081 21607 13139 21613
rect 13081 21604 13093 21607
rect 10560 21576 11468 21604
rect 11808 21576 13093 21604
rect 10560 21564 10566 21576
rect 2222 21536 2228 21548
rect 2183 21508 2228 21536
rect 2222 21496 2228 21508
rect 2280 21496 2286 21548
rect 7190 21496 7196 21548
rect 7248 21536 7254 21548
rect 7285 21539 7343 21545
rect 7285 21536 7297 21539
rect 7248 21508 7297 21536
rect 7248 21496 7254 21508
rect 7285 21505 7297 21508
rect 7331 21505 7343 21539
rect 7285 21499 7343 21505
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21536 7527 21539
rect 7650 21536 7656 21548
rect 7515 21508 7656 21536
rect 7515 21505 7527 21508
rect 7469 21499 7527 21505
rect 7650 21496 7656 21508
rect 7708 21536 7714 21548
rect 7837 21539 7895 21545
rect 7837 21536 7849 21539
rect 7708 21508 7849 21536
rect 7708 21496 7714 21508
rect 7837 21505 7849 21508
rect 7883 21536 7895 21539
rect 7926 21536 7932 21548
rect 7883 21508 7932 21536
rect 7883 21505 7895 21508
rect 7837 21499 7895 21505
rect 7926 21496 7932 21508
rect 7984 21496 7990 21548
rect 8294 21536 8300 21548
rect 8255 21508 8300 21536
rect 8294 21496 8300 21508
rect 8352 21496 8358 21548
rect 9125 21539 9183 21545
rect 9125 21505 9137 21539
rect 9171 21536 9183 21539
rect 9769 21539 9827 21545
rect 9769 21536 9781 21539
rect 9171 21508 9781 21536
rect 9171 21505 9183 21508
rect 9125 21499 9183 21505
rect 9769 21505 9781 21508
rect 9815 21536 9827 21539
rect 10870 21536 10876 21548
rect 9815 21508 10876 21536
rect 9815 21505 9827 21508
rect 9769 21499 9827 21505
rect 10870 21496 10876 21508
rect 10928 21496 10934 21548
rect 11330 21536 11336 21548
rect 11291 21508 11336 21536
rect 11330 21496 11336 21508
rect 11388 21496 11394 21548
rect 11440 21536 11468 21576
rect 13081 21573 13093 21576
rect 13127 21604 13139 21607
rect 13127 21576 13308 21604
rect 13127 21573 13139 21576
rect 13081 21567 13139 21573
rect 13280 21545 13308 21576
rect 20898 21564 20904 21616
rect 20956 21604 20962 21616
rect 22370 21604 22376 21616
rect 20956 21576 22376 21604
rect 20956 21564 20962 21576
rect 22370 21564 22376 21576
rect 22428 21564 22434 21616
rect 23566 21564 23572 21616
rect 23624 21564 23630 21616
rect 23845 21607 23903 21613
rect 23845 21573 23857 21607
rect 23891 21604 23903 21607
rect 24854 21604 24860 21616
rect 23891 21576 24860 21604
rect 23891 21573 23903 21576
rect 23845 21567 23903 21573
rect 24854 21564 24860 21576
rect 24912 21564 24918 21616
rect 13265 21539 13323 21545
rect 11440 21508 13032 21536
rect 3237 21471 3295 21477
rect 3237 21437 3249 21471
rect 3283 21468 3295 21471
rect 3326 21468 3332 21480
rect 3283 21440 3332 21468
rect 3283 21437 3295 21440
rect 3237 21431 3295 21437
rect 3326 21428 3332 21440
rect 3384 21468 3390 21480
rect 6086 21468 6092 21480
rect 3384 21440 6092 21468
rect 3384 21428 3390 21440
rect 6086 21428 6092 21440
rect 6144 21468 6150 21480
rect 6181 21471 6239 21477
rect 6181 21468 6193 21471
rect 6144 21440 6193 21468
rect 6144 21428 6150 21440
rect 6181 21437 6193 21440
rect 6227 21437 6239 21471
rect 6181 21431 6239 21437
rect 9585 21471 9643 21477
rect 9585 21437 9597 21471
rect 9631 21468 9643 21471
rect 9858 21468 9864 21480
rect 9631 21440 9864 21468
rect 9631 21437 9643 21440
rect 9585 21431 9643 21437
rect 9858 21428 9864 21440
rect 9916 21428 9922 21480
rect 11146 21468 11152 21480
rect 11107 21440 11152 21468
rect 11146 21428 11152 21440
rect 11204 21428 11210 21480
rect 12618 21468 12624 21480
rect 12579 21440 12624 21468
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 13004 21468 13032 21508
rect 13265 21505 13277 21539
rect 13311 21505 13323 21539
rect 15562 21536 15568 21548
rect 15475 21508 15568 21536
rect 13265 21499 13323 21505
rect 15562 21496 15568 21508
rect 15620 21536 15626 21548
rect 17037 21539 17095 21545
rect 17037 21536 17049 21539
rect 15620 21508 17049 21536
rect 15620 21496 15626 21508
rect 17037 21505 17049 21508
rect 17083 21536 17095 21539
rect 17402 21536 17408 21548
rect 17083 21508 17408 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 17402 21496 17408 21508
rect 17460 21496 17466 21548
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 20916 21508 22017 21536
rect 13354 21468 13360 21480
rect 13004 21440 13360 21468
rect 13354 21428 13360 21440
rect 13412 21468 13418 21480
rect 13532 21471 13590 21477
rect 13532 21468 13544 21471
rect 13412 21440 13544 21468
rect 13412 21428 13418 21440
rect 13532 21437 13544 21440
rect 13578 21468 13590 21471
rect 14366 21468 14372 21480
rect 13578 21440 14372 21468
rect 13578 21437 13590 21440
rect 13532 21431 13590 21437
rect 14366 21428 14372 21440
rect 14424 21428 14430 21480
rect 16298 21428 16304 21480
rect 16356 21468 16362 21480
rect 16853 21471 16911 21477
rect 16853 21468 16865 21471
rect 16356 21440 16865 21468
rect 16356 21428 16362 21440
rect 16853 21437 16865 21440
rect 16899 21437 16911 21471
rect 18969 21471 19027 21477
rect 18969 21468 18981 21471
rect 16853 21431 16911 21437
rect 18524 21440 18981 21468
rect 2041 21403 2099 21409
rect 2041 21369 2053 21403
rect 2087 21400 2099 21403
rect 2590 21400 2596 21412
rect 2087 21372 2596 21400
rect 2087 21369 2099 21372
rect 2041 21363 2099 21369
rect 2590 21360 2596 21372
rect 2648 21400 2654 21412
rect 3602 21409 3608 21412
rect 3596 21400 3608 21409
rect 2648 21372 2912 21400
rect 3563 21372 3608 21400
rect 2648 21360 2654 21372
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 1946 21332 1952 21344
rect 1907 21304 1952 21332
rect 1946 21292 1952 21304
rect 2004 21292 2010 21344
rect 2884 21332 2912 21372
rect 3596 21363 3608 21372
rect 3602 21360 3608 21363
rect 3660 21360 3666 21412
rect 6641 21403 6699 21409
rect 6641 21369 6653 21403
rect 6687 21400 6699 21403
rect 11241 21403 11299 21409
rect 11241 21400 11253 21403
rect 6687 21372 7236 21400
rect 6687 21369 6699 21372
rect 6641 21363 6699 21369
rect 7208 21344 7236 21372
rect 9232 21372 11253 21400
rect 3970 21332 3976 21344
rect 2884 21304 3976 21332
rect 3970 21292 3976 21304
rect 4028 21332 4034 21344
rect 4430 21332 4436 21344
rect 4028 21304 4436 21332
rect 4028 21292 4034 21304
rect 4430 21292 4436 21304
rect 4488 21292 4494 21344
rect 6454 21292 6460 21344
rect 6512 21332 6518 21344
rect 6825 21335 6883 21341
rect 6825 21332 6837 21335
rect 6512 21304 6837 21332
rect 6512 21292 6518 21304
rect 6825 21301 6837 21304
rect 6871 21301 6883 21335
rect 7190 21332 7196 21344
rect 7151 21304 7196 21332
rect 6825 21295 6883 21301
rect 7190 21292 7196 21304
rect 7248 21292 7254 21344
rect 8570 21332 8576 21344
rect 8531 21304 8576 21332
rect 8570 21292 8576 21304
rect 8628 21292 8634 21344
rect 9232 21341 9260 21372
rect 11241 21369 11253 21372
rect 11287 21400 11299 21403
rect 12894 21400 12900 21412
rect 11287 21372 12900 21400
rect 11287 21369 11299 21372
rect 11241 21363 11299 21369
rect 12894 21360 12900 21372
rect 12952 21360 12958 21412
rect 15933 21403 15991 21409
rect 15933 21369 15945 21403
rect 15979 21400 15991 21403
rect 16482 21400 16488 21412
rect 15979 21372 16488 21400
rect 15979 21369 15991 21372
rect 15933 21363 15991 21369
rect 16482 21360 16488 21372
rect 16540 21400 16546 21412
rect 17126 21400 17132 21412
rect 16540 21372 17132 21400
rect 16540 21360 16546 21372
rect 17126 21360 17132 21372
rect 17184 21360 17190 21412
rect 9217 21335 9275 21341
rect 9217 21301 9229 21335
rect 9263 21301 9275 21335
rect 9674 21332 9680 21344
rect 9635 21304 9680 21332
rect 9217 21295 9275 21301
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 9858 21292 9864 21344
rect 9916 21332 9922 21344
rect 10134 21332 10140 21344
rect 9916 21304 10140 21332
rect 9916 21292 9922 21304
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 10686 21292 10692 21344
rect 10744 21332 10750 21344
rect 10781 21335 10839 21341
rect 10781 21332 10793 21335
rect 10744 21304 10793 21332
rect 10744 21292 10750 21304
rect 10781 21301 10793 21304
rect 10827 21301 10839 21335
rect 10781 21295 10839 21301
rect 15286 21292 15292 21344
rect 15344 21332 15350 21344
rect 16301 21335 16359 21341
rect 16301 21332 16313 21335
rect 15344 21304 16313 21332
rect 15344 21292 15350 21304
rect 16301 21301 16313 21304
rect 16347 21332 16359 21335
rect 16758 21332 16764 21344
rect 16347 21304 16764 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 16758 21292 16764 21304
rect 16816 21292 16822 21344
rect 17310 21292 17316 21344
rect 17368 21332 17374 21344
rect 17405 21335 17463 21341
rect 17405 21332 17417 21335
rect 17368 21304 17417 21332
rect 17368 21292 17374 21304
rect 17405 21301 17417 21304
rect 17451 21301 17463 21335
rect 17405 21295 17463 21301
rect 17678 21292 17684 21344
rect 17736 21332 17742 21344
rect 18322 21332 18328 21344
rect 17736 21304 18328 21332
rect 17736 21292 17742 21304
rect 18322 21292 18328 21304
rect 18380 21332 18386 21344
rect 18524 21332 18552 21440
rect 18969 21437 18981 21440
rect 19015 21437 19027 21471
rect 18969 21431 19027 21437
rect 18598 21360 18604 21412
rect 18656 21400 18662 21412
rect 19150 21400 19156 21412
rect 18656 21372 19156 21400
rect 18656 21360 18662 21372
rect 19150 21360 19156 21372
rect 19208 21409 19214 21412
rect 19208 21403 19272 21409
rect 19208 21369 19226 21403
rect 19260 21369 19272 21403
rect 19208 21363 19272 21369
rect 19208 21360 19214 21363
rect 18785 21335 18843 21341
rect 18785 21332 18797 21335
rect 18380 21304 18797 21332
rect 18380 21292 18386 21304
rect 18785 21301 18797 21304
rect 18831 21301 18843 21335
rect 20346 21332 20352 21344
rect 20307 21304 20352 21332
rect 18785 21295 18843 21301
rect 20346 21292 20352 21304
rect 20404 21292 20410 21344
rect 20714 21292 20720 21344
rect 20772 21332 20778 21344
rect 20916 21341 20944 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 23584 21536 23612 21564
rect 24026 21536 24032 21548
rect 23584 21508 24032 21536
rect 22005 21499 22063 21505
rect 24026 21496 24032 21508
rect 24084 21496 24090 21548
rect 24486 21536 24492 21548
rect 24447 21508 24492 21536
rect 24486 21496 24492 21508
rect 24544 21496 24550 21548
rect 21542 21428 21548 21480
rect 21600 21468 21606 21480
rect 21821 21471 21879 21477
rect 21821 21468 21833 21471
rect 21600 21440 21833 21468
rect 21600 21428 21606 21440
rect 21821 21437 21833 21440
rect 21867 21437 21879 21471
rect 21821 21431 21879 21437
rect 23109 21471 23167 21477
rect 23109 21437 23121 21471
rect 23155 21468 23167 21471
rect 23566 21468 23572 21480
rect 23155 21440 23572 21468
rect 23155 21437 23167 21440
rect 23109 21431 23167 21437
rect 23566 21428 23572 21440
rect 23624 21468 23630 21480
rect 24213 21471 24271 21477
rect 24213 21468 24225 21471
rect 23624 21440 24225 21468
rect 23624 21428 23630 21440
rect 24213 21437 24225 21440
rect 24259 21468 24271 21471
rect 24762 21468 24768 21480
rect 24259 21440 24768 21468
rect 24259 21437 24271 21440
rect 24213 21431 24271 21437
rect 24762 21428 24768 21440
rect 24820 21428 24826 21480
rect 25314 21428 25320 21480
rect 25372 21468 25378 21480
rect 25409 21471 25467 21477
rect 25409 21468 25421 21471
rect 25372 21440 25421 21468
rect 25372 21428 25378 21440
rect 25409 21437 25421 21440
rect 25455 21468 25467 21471
rect 25961 21471 26019 21477
rect 25961 21468 25973 21471
rect 25455 21440 25973 21468
rect 25455 21437 25467 21440
rect 25409 21431 25467 21437
rect 25961 21437 25973 21440
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 21913 21403 21971 21409
rect 21913 21400 21925 21403
rect 21284 21372 21925 21400
rect 21284 21344 21312 21372
rect 21913 21369 21925 21372
rect 21959 21369 21971 21403
rect 24118 21400 24124 21412
rect 21913 21363 21971 21369
rect 23492 21372 24124 21400
rect 23492 21344 23520 21372
rect 24118 21360 24124 21372
rect 24176 21400 24182 21412
rect 24305 21403 24363 21409
rect 24305 21400 24317 21403
rect 24176 21372 24317 21400
rect 24176 21360 24182 21372
rect 24305 21369 24317 21372
rect 24351 21369 24363 21403
rect 24305 21363 24363 21369
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20772 21304 20913 21332
rect 20772 21292 20778 21304
rect 20901 21301 20913 21304
rect 20947 21301 20959 21335
rect 21266 21332 21272 21344
rect 21227 21304 21272 21332
rect 20901 21295 20959 21301
rect 21266 21292 21272 21304
rect 21324 21292 21330 21344
rect 21453 21335 21511 21341
rect 21453 21301 21465 21335
rect 21499 21332 21511 21335
rect 21726 21332 21732 21344
rect 21499 21304 21732 21332
rect 21499 21301 21511 21304
rect 21453 21295 21511 21301
rect 21726 21292 21732 21304
rect 21784 21292 21790 21344
rect 23474 21332 23480 21344
rect 23435 21304 23480 21332
rect 23474 21292 23480 21304
rect 23532 21292 23538 21344
rect 25038 21332 25044 21344
rect 24999 21304 25044 21332
rect 25038 21292 25044 21304
rect 25096 21292 25102 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1486 21088 1492 21140
rect 1544 21088 1550 21140
rect 1762 21088 1768 21140
rect 1820 21128 1826 21140
rect 1857 21131 1915 21137
rect 1857 21128 1869 21131
rect 1820 21100 1869 21128
rect 1820 21088 1826 21100
rect 1857 21097 1869 21100
rect 1903 21097 1915 21131
rect 2406 21128 2412 21140
rect 2367 21100 2412 21128
rect 1857 21091 1915 21097
rect 1504 21060 1532 21088
rect 1504 21032 1808 21060
rect 1394 20924 1400 20936
rect 1355 20896 1400 20924
rect 1394 20884 1400 20896
rect 1452 20884 1458 20936
rect 1780 20924 1808 21032
rect 1872 20992 1900 21091
rect 2406 21088 2412 21100
rect 2464 21088 2470 21140
rect 3326 21088 3332 21140
rect 3384 21128 3390 21140
rect 3697 21131 3755 21137
rect 3697 21128 3709 21131
rect 3384 21100 3709 21128
rect 3384 21088 3390 21100
rect 3697 21097 3709 21100
rect 3743 21097 3755 21131
rect 3697 21091 3755 21097
rect 3881 21131 3939 21137
rect 3881 21097 3893 21131
rect 3927 21128 3939 21131
rect 4430 21128 4436 21140
rect 3927 21100 4436 21128
rect 3927 21097 3939 21100
rect 3881 21091 3939 21097
rect 4430 21088 4436 21100
rect 4488 21088 4494 21140
rect 4706 21088 4712 21140
rect 4764 21128 4770 21140
rect 5997 21131 6055 21137
rect 5997 21128 6009 21131
rect 4764 21100 6009 21128
rect 4764 21088 4770 21100
rect 5997 21097 6009 21100
rect 6043 21097 6055 21131
rect 6362 21128 6368 21140
rect 6323 21100 6368 21128
rect 5997 21091 6055 21097
rect 6362 21088 6368 21100
rect 6420 21088 6426 21140
rect 7377 21131 7435 21137
rect 7377 21097 7389 21131
rect 7423 21128 7435 21131
rect 7650 21128 7656 21140
rect 7423 21100 7656 21128
rect 7423 21097 7435 21100
rect 7377 21091 7435 21097
rect 7650 21088 7656 21100
rect 7708 21088 7714 21140
rect 9953 21131 10011 21137
rect 9953 21097 9965 21131
rect 9999 21128 10011 21131
rect 10042 21128 10048 21140
rect 9999 21100 10048 21128
rect 9999 21097 10011 21100
rect 9953 21091 10011 21097
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 10505 21131 10563 21137
rect 10505 21097 10517 21131
rect 10551 21128 10563 21131
rect 11146 21128 11152 21140
rect 10551 21100 11152 21128
rect 10551 21097 10563 21100
rect 10505 21091 10563 21097
rect 11146 21088 11152 21100
rect 11204 21088 11210 21140
rect 11514 21128 11520 21140
rect 11475 21100 11520 21128
rect 11514 21088 11520 21100
rect 11572 21088 11578 21140
rect 12069 21131 12127 21137
rect 12069 21097 12081 21131
rect 12115 21128 12127 21131
rect 12158 21128 12164 21140
rect 12115 21100 12164 21128
rect 12115 21097 12127 21100
rect 12069 21091 12127 21097
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 12342 21088 12348 21140
rect 12400 21128 12406 21140
rect 12526 21128 12532 21140
rect 12400 21100 12532 21128
rect 12400 21088 12406 21100
rect 12526 21088 12532 21100
rect 12584 21088 12590 21140
rect 13354 21128 13360 21140
rect 13315 21100 13360 21128
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 13633 21131 13691 21137
rect 13633 21097 13645 21131
rect 13679 21128 13691 21131
rect 15654 21128 15660 21140
rect 13679 21100 15516 21128
rect 15615 21100 15660 21128
rect 13679 21097 13691 21100
rect 13633 21091 13691 21097
rect 2317 21063 2375 21069
rect 2317 21029 2329 21063
rect 2363 21060 2375 21063
rect 2590 21060 2596 21072
rect 2363 21032 2596 21060
rect 2363 21029 2375 21032
rect 2317 21023 2375 21029
rect 2590 21020 2596 21032
rect 2648 21020 2654 21072
rect 2777 21063 2835 21069
rect 2777 21029 2789 21063
rect 2823 21060 2835 21063
rect 4062 21060 4068 21072
rect 2823 21032 4068 21060
rect 2823 21029 2835 21032
rect 2777 21023 2835 21029
rect 4062 21020 4068 21032
rect 4120 21020 4126 21072
rect 8021 21063 8079 21069
rect 8021 21060 8033 21063
rect 7024 21032 8033 21060
rect 7024 21004 7052 21032
rect 8021 21029 8033 21032
rect 8067 21029 8079 21063
rect 10962 21060 10968 21072
rect 10923 21032 10968 21060
rect 8021 21023 8079 21029
rect 10962 21020 10968 21032
rect 11020 21020 11026 21072
rect 11977 21063 12035 21069
rect 11977 21029 11989 21063
rect 12023 21060 12035 21063
rect 12360 21060 12388 21088
rect 12023 21032 12388 21060
rect 14001 21063 14059 21069
rect 12023 21029 12035 21032
rect 11977 21023 12035 21029
rect 14001 21029 14013 21063
rect 14047 21060 14059 21063
rect 14274 21060 14280 21072
rect 14047 21032 14280 21060
rect 14047 21029 14059 21032
rect 14001 21023 14059 21029
rect 14274 21020 14280 21032
rect 14332 21020 14338 21072
rect 15488 21060 15516 21100
rect 15654 21088 15660 21100
rect 15712 21088 15718 21140
rect 15930 21088 15936 21140
rect 15988 21088 15994 21140
rect 16298 21088 16304 21140
rect 16356 21128 16362 21140
rect 16393 21131 16451 21137
rect 16393 21128 16405 21131
rect 16356 21100 16405 21128
rect 16356 21088 16362 21100
rect 16393 21097 16405 21100
rect 16439 21097 16451 21131
rect 16393 21091 16451 21097
rect 17862 21088 17868 21140
rect 17920 21128 17926 21140
rect 18969 21131 19027 21137
rect 18969 21128 18981 21131
rect 17920 21100 18981 21128
rect 17920 21088 17926 21100
rect 18969 21097 18981 21100
rect 19015 21097 19027 21131
rect 18969 21091 19027 21097
rect 15948 21060 15976 21088
rect 16942 21069 16948 21072
rect 16936 21060 16948 21069
rect 15488 21032 15976 21060
rect 16855 21032 16948 21060
rect 16936 21023 16948 21032
rect 17000 21060 17006 21072
rect 17402 21060 17408 21072
rect 17000 21032 17408 21060
rect 16942 21020 16948 21023
rect 17000 21020 17006 21032
rect 17402 21020 17408 21032
rect 17460 21020 17466 21072
rect 18598 21060 18604 21072
rect 18559 21032 18604 21060
rect 18598 21020 18604 21032
rect 18656 21020 18662 21072
rect 2869 20995 2927 21001
rect 1872 20964 2820 20992
rect 2792 20936 2820 20964
rect 2869 20961 2881 20995
rect 2915 20992 2927 20995
rect 3326 20992 3332 21004
rect 2915 20964 3332 20992
rect 2915 20961 2927 20964
rect 2869 20955 2927 20961
rect 3326 20952 3332 20964
rect 3384 20952 3390 21004
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4321 20995 4379 21001
rect 4321 20992 4333 20995
rect 4212 20964 4333 20992
rect 4212 20952 4218 20964
rect 4321 20961 4333 20964
rect 4367 20961 4379 20995
rect 4321 20955 4379 20961
rect 7006 20952 7012 21004
rect 7064 20952 7070 21004
rect 7466 20952 7472 21004
rect 7524 20992 7530 21004
rect 7742 20992 7748 21004
rect 7524 20964 7748 20992
rect 7524 20952 7530 20964
rect 7742 20952 7748 20964
rect 7800 20952 7806 21004
rect 8294 20952 8300 21004
rect 8352 20992 8358 21004
rect 9582 20992 9588 21004
rect 8352 20964 9588 20992
rect 8352 20952 8358 20964
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 10870 20992 10876 21004
rect 10831 20964 10876 20992
rect 10870 20952 10876 20964
rect 10928 20952 10934 21004
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 14093 20995 14151 21001
rect 12492 20964 12537 20992
rect 12492 20952 12498 20964
rect 14093 20961 14105 20995
rect 14139 20992 14151 20995
rect 14826 20992 14832 21004
rect 14139 20964 14832 20992
rect 14139 20961 14151 20964
rect 14093 20955 14151 20961
rect 14826 20952 14832 20964
rect 14884 20952 14890 21004
rect 15473 20995 15531 21001
rect 15473 20961 15485 20995
rect 15519 20992 15531 20995
rect 15838 20992 15844 21004
rect 15519 20964 15844 20992
rect 15519 20961 15531 20964
rect 15473 20955 15531 20961
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 16114 20952 16120 21004
rect 16172 20992 16178 21004
rect 16669 20995 16727 21001
rect 16669 20992 16681 20995
rect 16172 20964 16681 20992
rect 16172 20952 16178 20964
rect 16669 20961 16681 20964
rect 16715 20961 16727 20995
rect 16669 20955 16727 20961
rect 1780 20896 2452 20924
rect 2424 20800 2452 20896
rect 2774 20884 2780 20936
rect 2832 20884 2838 20936
rect 3053 20927 3111 20933
rect 3053 20893 3065 20927
rect 3099 20924 3111 20927
rect 3237 20927 3295 20933
rect 3237 20924 3249 20927
rect 3099 20896 3249 20924
rect 3099 20893 3111 20896
rect 3053 20887 3111 20893
rect 3237 20893 3249 20896
rect 3283 20893 3295 20927
rect 3237 20887 3295 20893
rect 3510 20884 3516 20936
rect 3568 20924 3574 20936
rect 3697 20927 3755 20933
rect 3697 20924 3709 20927
rect 3568 20896 3709 20924
rect 3568 20884 3574 20896
rect 3697 20893 3709 20896
rect 3743 20924 3755 20927
rect 4065 20927 4123 20933
rect 4065 20924 4077 20927
rect 3743 20896 4077 20924
rect 3743 20893 3755 20896
rect 3697 20887 3755 20893
rect 4065 20893 4077 20896
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 5350 20884 5356 20936
rect 5408 20924 5414 20936
rect 7558 20924 7564 20936
rect 5408 20896 7144 20924
rect 7519 20896 7564 20924
rect 5408 20884 5414 20896
rect 6914 20856 6920 20868
rect 6875 20828 6920 20856
rect 6914 20816 6920 20828
rect 6972 20816 6978 20868
rect 7116 20856 7144 20896
rect 7558 20884 7564 20896
rect 7616 20884 7622 20936
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20924 8631 20927
rect 8938 20924 8944 20936
rect 8619 20896 8944 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 11054 20924 11060 20936
rect 11015 20896 11060 20924
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 12342 20884 12348 20936
rect 12400 20924 12406 20936
rect 12529 20927 12587 20933
rect 12529 20924 12541 20927
rect 12400 20896 12541 20924
rect 12400 20884 12406 20896
rect 12529 20893 12541 20896
rect 12575 20893 12587 20927
rect 12710 20924 12716 20936
rect 12671 20896 12716 20924
rect 12529 20887 12587 20893
rect 9401 20859 9459 20865
rect 9401 20856 9413 20859
rect 7116 20828 9413 20856
rect 9401 20825 9413 20828
rect 9447 20825 9459 20859
rect 12544 20856 12572 20887
rect 12710 20884 12716 20896
rect 12768 20924 12774 20936
rect 14185 20927 14243 20933
rect 14185 20924 14197 20927
rect 12768 20896 14197 20924
rect 12768 20884 12774 20896
rect 14185 20893 14197 20896
rect 14231 20893 14243 20927
rect 14185 20887 14243 20893
rect 13446 20856 13452 20868
rect 12544 20828 13452 20856
rect 9401 20819 9459 20825
rect 13446 20816 13452 20828
rect 13504 20816 13510 20868
rect 14918 20816 14924 20868
rect 14976 20816 14982 20868
rect 18984 20856 19012 21091
rect 19058 21088 19064 21140
rect 19116 21128 19122 21140
rect 19153 21131 19211 21137
rect 19153 21128 19165 21131
rect 19116 21100 19165 21128
rect 19116 21088 19122 21100
rect 19153 21097 19165 21100
rect 19199 21097 19211 21131
rect 22738 21128 22744 21140
rect 22699 21100 22744 21128
rect 19153 21091 19211 21097
rect 22738 21088 22744 21100
rect 22796 21088 22802 21140
rect 23201 21131 23259 21137
rect 23201 21097 23213 21131
rect 23247 21128 23259 21131
rect 23934 21128 23940 21140
rect 23247 21100 23940 21128
rect 23247 21097 23259 21100
rect 23201 21091 23259 21097
rect 23934 21088 23940 21100
rect 23992 21088 23998 21140
rect 22005 21063 22063 21069
rect 22005 21029 22017 21063
rect 22051 21060 22063 21063
rect 22186 21060 22192 21072
rect 22051 21032 22192 21060
rect 22051 21029 22063 21032
rect 22005 21023 22063 21029
rect 22186 21020 22192 21032
rect 22244 21020 22250 21072
rect 22373 21063 22431 21069
rect 22373 21029 22385 21063
rect 22419 21060 22431 21063
rect 22922 21060 22928 21072
rect 22419 21032 22928 21060
rect 22419 21029 22431 21032
rect 22373 21023 22431 21029
rect 22922 21020 22928 21032
rect 22980 21020 22986 21072
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 19521 20995 19579 21001
rect 19521 20992 19533 20995
rect 19392 20964 19533 20992
rect 19392 20952 19398 20964
rect 19521 20961 19533 20964
rect 19567 20992 19579 20995
rect 20165 20995 20223 21001
rect 20165 20992 20177 20995
rect 19567 20964 20177 20992
rect 19567 20961 19579 20964
rect 19521 20955 19579 20961
rect 20165 20961 20177 20964
rect 20211 20961 20223 20995
rect 20165 20955 20223 20961
rect 21174 20952 21180 21004
rect 21232 20992 21238 21004
rect 21269 20995 21327 21001
rect 21269 20992 21281 20995
rect 21232 20964 21281 20992
rect 21232 20952 21238 20964
rect 21269 20961 21281 20964
rect 21315 20961 21327 20995
rect 22554 20992 22560 21004
rect 22515 20964 22560 20992
rect 21269 20955 21327 20961
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 23934 20952 23940 21004
rect 23992 20992 23998 21004
rect 24305 20995 24363 21001
rect 24305 20992 24317 20995
rect 23992 20964 24317 20992
rect 23992 20952 23998 20964
rect 24305 20961 24317 20964
rect 24351 20961 24363 20995
rect 24305 20955 24363 20961
rect 24397 20995 24455 21001
rect 24397 20961 24409 20995
rect 24443 20992 24455 20995
rect 24670 20992 24676 21004
rect 24443 20964 24676 20992
rect 24443 20961 24455 20964
rect 24397 20955 24455 20961
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 19610 20924 19616 20936
rect 19571 20896 19616 20924
rect 19610 20884 19616 20896
rect 19668 20884 19674 20936
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20924 19763 20927
rect 20346 20924 20352 20936
rect 19751 20896 20352 20924
rect 19751 20893 19763 20896
rect 19705 20887 19763 20893
rect 19720 20856 19748 20887
rect 20346 20884 20352 20896
rect 20404 20884 20410 20936
rect 20714 20924 20720 20936
rect 20675 20896 20720 20924
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 21358 20924 21364 20936
rect 21319 20896 21364 20924
rect 21358 20884 21364 20896
rect 21416 20884 21422 20936
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 18984 20828 19748 20856
rect 20732 20856 20760 20884
rect 21468 20856 21496 20887
rect 24210 20884 24216 20936
rect 24268 20924 24274 20936
rect 24486 20924 24492 20936
rect 24268 20896 24492 20924
rect 24268 20884 24274 20896
rect 24486 20884 24492 20896
rect 24544 20884 24550 20936
rect 20732 20828 21496 20856
rect 2406 20748 2412 20800
rect 2464 20748 2470 20800
rect 3237 20791 3295 20797
rect 3237 20757 3249 20791
rect 3283 20788 3295 20791
rect 3513 20791 3571 20797
rect 3513 20788 3525 20791
rect 3283 20760 3525 20788
rect 3283 20757 3295 20760
rect 3237 20751 3295 20757
rect 3513 20757 3525 20760
rect 3559 20788 3571 20791
rect 3602 20788 3608 20800
rect 3559 20760 3608 20788
rect 3559 20757 3571 20760
rect 3513 20751 3571 20757
rect 3602 20748 3608 20760
rect 3660 20788 3666 20800
rect 5442 20788 5448 20800
rect 3660 20760 5448 20788
rect 3660 20748 3666 20760
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 7006 20788 7012 20800
rect 6967 20760 7012 20788
rect 7006 20748 7012 20760
rect 7064 20748 7070 20800
rect 8386 20788 8392 20800
rect 8347 20760 8392 20788
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 9030 20788 9036 20800
rect 8991 20760 9036 20788
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 10226 20788 10232 20800
rect 10187 20760 10232 20788
rect 10226 20748 10232 20760
rect 10284 20748 10290 20800
rect 14366 20748 14372 20800
rect 14424 20788 14430 20800
rect 14645 20791 14703 20797
rect 14645 20788 14657 20791
rect 14424 20760 14657 20788
rect 14424 20748 14430 20760
rect 14645 20757 14657 20760
rect 14691 20788 14703 20791
rect 14936 20788 14964 20816
rect 14691 20760 14964 20788
rect 15105 20791 15163 20797
rect 14691 20757 14703 20760
rect 14645 20751 14703 20757
rect 15105 20757 15117 20791
rect 15151 20788 15163 20791
rect 15378 20788 15384 20800
rect 15151 20760 15384 20788
rect 15151 20757 15163 20760
rect 15105 20751 15163 20757
rect 15378 20748 15384 20760
rect 15436 20748 15442 20800
rect 16022 20788 16028 20800
rect 15983 20760 16028 20788
rect 16022 20748 16028 20760
rect 16080 20788 16086 20800
rect 18049 20791 18107 20797
rect 18049 20788 18061 20791
rect 16080 20760 18061 20788
rect 16080 20748 16086 20760
rect 18049 20757 18061 20760
rect 18095 20757 18107 20791
rect 18049 20751 18107 20757
rect 20714 20748 20720 20800
rect 20772 20788 20778 20800
rect 20901 20791 20959 20797
rect 20901 20788 20913 20791
rect 20772 20760 20913 20788
rect 20772 20748 20778 20760
rect 20901 20757 20913 20760
rect 20947 20757 20959 20791
rect 20901 20751 20959 20757
rect 21818 20748 21824 20800
rect 21876 20788 21882 20800
rect 22094 20788 22100 20800
rect 21876 20760 22100 20788
rect 21876 20748 21882 20760
rect 22094 20748 22100 20760
rect 22152 20748 22158 20800
rect 23569 20791 23627 20797
rect 23569 20757 23581 20791
rect 23615 20788 23627 20791
rect 23750 20788 23756 20800
rect 23615 20760 23756 20788
rect 23615 20757 23627 20760
rect 23569 20751 23627 20757
rect 23750 20748 23756 20760
rect 23808 20748 23814 20800
rect 23937 20791 23995 20797
rect 23937 20757 23949 20791
rect 23983 20788 23995 20791
rect 24026 20788 24032 20800
rect 23983 20760 24032 20788
rect 23983 20757 23995 20760
rect 23937 20751 23995 20757
rect 24026 20748 24032 20760
rect 24084 20788 24090 20800
rect 24949 20791 25007 20797
rect 24949 20788 24961 20791
rect 24084 20760 24961 20788
rect 24084 20748 24090 20760
rect 24949 20757 24961 20760
rect 24995 20757 25007 20791
rect 24949 20751 25007 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1854 20544 1860 20596
rect 1912 20584 1918 20596
rect 1949 20587 2007 20593
rect 1949 20584 1961 20587
rect 1912 20556 1961 20584
rect 1912 20544 1918 20556
rect 1949 20553 1961 20556
rect 1995 20553 2007 20587
rect 1949 20547 2007 20553
rect 2222 20544 2228 20596
rect 2280 20584 2286 20596
rect 2317 20587 2375 20593
rect 2317 20584 2329 20587
rect 2280 20556 2329 20584
rect 2280 20544 2286 20556
rect 2317 20553 2329 20556
rect 2363 20553 2375 20587
rect 2317 20547 2375 20553
rect 2869 20587 2927 20593
rect 2869 20553 2881 20587
rect 2915 20584 2927 20587
rect 3326 20584 3332 20596
rect 2915 20556 3332 20584
rect 2915 20553 2927 20556
rect 2869 20547 2927 20553
rect 3326 20544 3332 20556
rect 3384 20544 3390 20596
rect 3510 20544 3516 20596
rect 3568 20584 3574 20596
rect 4157 20587 4215 20593
rect 4157 20584 4169 20587
rect 3568 20556 4169 20584
rect 3568 20544 3574 20556
rect 4157 20553 4169 20556
rect 4203 20553 4215 20587
rect 4157 20547 4215 20553
rect 4433 20587 4491 20593
rect 4433 20553 4445 20587
rect 4479 20584 4491 20587
rect 4522 20584 4528 20596
rect 4479 20556 4528 20584
rect 4479 20553 4491 20556
rect 4433 20547 4491 20553
rect 4522 20544 4528 20556
rect 4580 20544 4586 20596
rect 6822 20584 6828 20596
rect 4908 20556 6828 20584
rect 2314 20408 2320 20460
rect 2372 20448 2378 20460
rect 2682 20448 2688 20460
rect 2372 20420 2688 20448
rect 2372 20408 2378 20420
rect 2682 20408 2688 20420
rect 2740 20408 2746 20460
rect 3326 20448 3332 20460
rect 3287 20420 3332 20448
rect 3326 20408 3332 20420
rect 3384 20408 3390 20460
rect 3421 20451 3479 20457
rect 3421 20417 3433 20451
rect 3467 20448 3479 20451
rect 4154 20448 4160 20460
rect 3467 20420 4160 20448
rect 3467 20417 3479 20420
rect 3421 20411 3479 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1854 20380 1860 20392
rect 1443 20352 1860 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1854 20340 1860 20352
rect 1912 20340 1918 20392
rect 2777 20383 2835 20389
rect 2777 20349 2789 20383
rect 2823 20380 2835 20383
rect 3436 20380 3464 20411
rect 4154 20408 4160 20420
rect 4212 20408 4218 20460
rect 4908 20457 4936 20556
rect 6822 20544 6828 20556
rect 6880 20544 6886 20596
rect 9582 20544 9588 20596
rect 9640 20584 9646 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 9640 20556 9965 20584
rect 9640 20544 9646 20556
rect 9953 20553 9965 20556
rect 9999 20553 10011 20587
rect 9953 20547 10011 20553
rect 10597 20587 10655 20593
rect 10597 20553 10609 20587
rect 10643 20584 10655 20587
rect 10962 20584 10968 20596
rect 10643 20556 10968 20584
rect 10643 20553 10655 20556
rect 10597 20547 10655 20553
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 14274 20544 14280 20596
rect 14332 20584 14338 20596
rect 14369 20587 14427 20593
rect 14369 20584 14381 20587
rect 14332 20556 14381 20584
rect 14332 20544 14338 20556
rect 14369 20553 14381 20556
rect 14415 20553 14427 20587
rect 14826 20584 14832 20596
rect 14787 20556 14832 20584
rect 14369 20547 14427 20553
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 15289 20587 15347 20593
rect 15289 20553 15301 20587
rect 15335 20584 15347 20587
rect 16114 20584 16120 20596
rect 15335 20556 16120 20584
rect 15335 20553 15347 20556
rect 15289 20547 15347 20553
rect 5442 20516 5448 20528
rect 5092 20488 5448 20516
rect 5092 20457 5120 20488
rect 5442 20476 5448 20488
rect 5500 20516 5506 20528
rect 5813 20519 5871 20525
rect 5813 20516 5825 20519
rect 5500 20488 5825 20516
rect 5500 20476 5506 20488
rect 5813 20485 5825 20488
rect 5859 20485 5871 20519
rect 6270 20516 6276 20528
rect 6183 20488 6276 20516
rect 5813 20479 5871 20485
rect 6270 20476 6276 20488
rect 6328 20516 6334 20528
rect 7558 20516 7564 20528
rect 6328 20488 7564 20516
rect 6328 20476 6334 20488
rect 7558 20476 7564 20488
rect 7616 20476 7622 20528
rect 4893 20451 4951 20457
rect 4893 20417 4905 20451
rect 4939 20417 4951 20451
rect 4893 20411 4951 20417
rect 5077 20451 5135 20457
rect 5077 20417 5089 20451
rect 5123 20417 5135 20451
rect 5077 20411 5135 20417
rect 7006 20408 7012 20460
rect 7064 20448 7070 20460
rect 15396 20457 15424 20556
rect 16114 20544 16120 20556
rect 16172 20584 16178 20596
rect 17313 20587 17371 20593
rect 17313 20584 17325 20587
rect 16172 20556 17325 20584
rect 16172 20544 16178 20556
rect 17313 20553 17325 20556
rect 17359 20584 17371 20587
rect 17678 20584 17684 20596
rect 17359 20556 17684 20584
rect 17359 20553 17371 20556
rect 17313 20547 17371 20553
rect 17678 20544 17684 20556
rect 17736 20544 17742 20596
rect 17862 20584 17868 20596
rect 17823 20556 17868 20584
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 18233 20587 18291 20593
rect 18233 20553 18245 20587
rect 18279 20584 18291 20587
rect 18966 20584 18972 20596
rect 18279 20556 18972 20584
rect 18279 20553 18291 20556
rect 18233 20547 18291 20553
rect 18966 20544 18972 20556
rect 19024 20544 19030 20596
rect 19153 20587 19211 20593
rect 19153 20553 19165 20587
rect 19199 20584 19211 20587
rect 19242 20584 19248 20596
rect 19199 20556 19248 20584
rect 19199 20553 19211 20556
rect 19153 20547 19211 20553
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 22186 20544 22192 20596
rect 22244 20584 22250 20596
rect 22281 20587 22339 20593
rect 22281 20584 22293 20587
rect 22244 20556 22293 20584
rect 22244 20544 22250 20556
rect 22281 20553 22293 20556
rect 22327 20553 22339 20587
rect 22281 20547 22339 20553
rect 22554 20544 22560 20596
rect 22612 20584 22618 20596
rect 22833 20587 22891 20593
rect 22833 20584 22845 20587
rect 22612 20556 22845 20584
rect 22612 20544 22618 20556
rect 22833 20553 22845 20556
rect 22879 20553 22891 20587
rect 25406 20584 25412 20596
rect 25367 20556 25412 20584
rect 22833 20547 22891 20553
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 7285 20451 7343 20457
rect 7285 20448 7297 20451
rect 7064 20420 7297 20448
rect 7064 20408 7070 20420
rect 7285 20417 7297 20420
rect 7331 20417 7343 20451
rect 7285 20411 7343 20417
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 15381 20451 15439 20457
rect 15381 20417 15393 20451
rect 15427 20417 15439 20451
rect 15381 20411 15439 20417
rect 7392 20380 7420 20411
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 19392 20420 19717 20448
rect 19392 20408 19398 20420
rect 19705 20417 19717 20420
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 20346 20408 20352 20460
rect 20404 20448 20410 20460
rect 20901 20451 20959 20457
rect 20901 20448 20913 20451
rect 20404 20420 20913 20448
rect 20404 20408 20410 20420
rect 20901 20417 20913 20420
rect 20947 20417 20959 20451
rect 20901 20411 20959 20417
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20448 24363 20451
rect 24670 20448 24676 20460
rect 24351 20420 24532 20448
rect 24631 20420 24676 20448
rect 24351 20417 24363 20420
rect 24305 20411 24363 20417
rect 2823 20352 3464 20380
rect 6932 20352 7420 20380
rect 8573 20383 8631 20389
rect 2823 20349 2835 20352
rect 2777 20343 2835 20349
rect 6932 20324 6960 20352
rect 8573 20349 8585 20383
rect 8619 20349 8631 20383
rect 8573 20343 8631 20349
rect 11057 20383 11115 20389
rect 11057 20349 11069 20383
rect 11103 20380 11115 20383
rect 11606 20380 11612 20392
rect 11103 20352 11612 20380
rect 11103 20349 11115 20352
rect 11057 20343 11115 20349
rect 3234 20312 3240 20324
rect 3195 20284 3240 20312
rect 3234 20272 3240 20284
rect 3292 20272 3298 20324
rect 6914 20312 6920 20324
rect 5460 20284 6920 20312
rect 5460 20256 5488 20284
rect 6914 20272 6920 20284
rect 6972 20272 6978 20324
rect 7466 20312 7472 20324
rect 7024 20284 7472 20312
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 2590 20204 2596 20256
rect 2648 20244 2654 20256
rect 4430 20244 4436 20256
rect 2648 20216 4436 20244
rect 2648 20204 2654 20216
rect 4430 20204 4436 20216
rect 4488 20204 4494 20256
rect 4798 20244 4804 20256
rect 4759 20216 4804 20244
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 5442 20244 5448 20256
rect 5403 20216 5448 20244
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 6641 20247 6699 20253
rect 6641 20213 6653 20247
rect 6687 20244 6699 20247
rect 7024 20244 7052 20284
rect 7466 20272 7472 20284
rect 7524 20272 7530 20324
rect 7190 20244 7196 20256
rect 6687 20216 7052 20244
rect 7151 20216 7196 20244
rect 6687 20213 6699 20216
rect 6641 20207 6699 20213
rect 7190 20204 7196 20216
rect 7248 20204 7254 20256
rect 7650 20204 7656 20256
rect 7708 20244 7714 20256
rect 7929 20247 7987 20253
rect 7929 20244 7941 20247
rect 7708 20216 7941 20244
rect 7708 20204 7714 20216
rect 7929 20213 7941 20216
rect 7975 20244 7987 20247
rect 8018 20244 8024 20256
rect 7975 20216 8024 20244
rect 7975 20213 7987 20216
rect 7929 20207 7987 20213
rect 8018 20204 8024 20216
rect 8076 20204 8082 20256
rect 8481 20247 8539 20253
rect 8481 20213 8493 20247
rect 8527 20244 8539 20247
rect 8588 20244 8616 20343
rect 11606 20340 11612 20352
rect 11664 20340 11670 20392
rect 12250 20340 12256 20392
rect 12308 20380 12314 20392
rect 12437 20383 12495 20389
rect 12437 20380 12449 20383
rect 12308 20352 12449 20380
rect 12308 20340 12314 20352
rect 12437 20349 12449 20352
rect 12483 20349 12495 20383
rect 12437 20343 12495 20349
rect 12526 20340 12532 20392
rect 12584 20380 12590 20392
rect 12693 20383 12751 20389
rect 12693 20380 12705 20383
rect 12584 20352 12705 20380
rect 12584 20340 12590 20352
rect 12693 20349 12705 20352
rect 12739 20349 12751 20383
rect 12693 20343 12751 20349
rect 15648 20383 15706 20389
rect 15648 20349 15660 20383
rect 15694 20380 15706 20383
rect 16022 20380 16028 20392
rect 15694 20352 16028 20380
rect 15694 20349 15706 20352
rect 15648 20343 15706 20349
rect 16022 20340 16028 20352
rect 16080 20340 16086 20392
rect 18046 20380 18052 20392
rect 18007 20352 18052 20380
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 18693 20383 18751 20389
rect 18693 20349 18705 20383
rect 18739 20380 18751 20383
rect 19521 20383 19579 20389
rect 19521 20380 19533 20383
rect 18739 20352 19533 20380
rect 18739 20349 18751 20352
rect 18693 20343 18751 20349
rect 19521 20349 19533 20352
rect 19567 20380 19579 20383
rect 20806 20380 20812 20392
rect 19567 20352 20812 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 20806 20340 20812 20352
rect 20864 20340 20870 20392
rect 24026 20380 24032 20392
rect 23987 20352 24032 20380
rect 24026 20340 24032 20352
rect 24084 20340 24090 20392
rect 8846 20321 8852 20324
rect 8840 20312 8852 20321
rect 8807 20284 8852 20312
rect 8840 20275 8852 20284
rect 8846 20272 8852 20275
rect 8904 20272 8910 20324
rect 9122 20272 9128 20324
rect 9180 20312 9186 20324
rect 12069 20315 12127 20321
rect 12069 20312 12081 20315
rect 9180 20284 12081 20312
rect 9180 20272 9186 20284
rect 12069 20281 12081 20284
rect 12115 20312 12127 20315
rect 12342 20312 12348 20324
rect 12115 20284 12348 20312
rect 12115 20281 12127 20284
rect 12069 20275 12127 20281
rect 12342 20272 12348 20284
rect 12400 20272 12406 20324
rect 17678 20272 17684 20324
rect 17736 20312 17742 20324
rect 20346 20312 20352 20324
rect 17736 20284 20352 20312
rect 17736 20272 17742 20284
rect 20346 20272 20352 20284
rect 20404 20272 20410 20324
rect 21146 20315 21204 20321
rect 21146 20312 21158 20315
rect 20916 20284 21158 20312
rect 20916 20256 20944 20284
rect 21146 20281 21158 20284
rect 21192 20281 21204 20315
rect 21146 20275 21204 20281
rect 23477 20315 23535 20321
rect 23477 20281 23489 20315
rect 23523 20312 23535 20315
rect 23934 20312 23940 20324
rect 23523 20284 23940 20312
rect 23523 20281 23535 20284
rect 23477 20275 23535 20281
rect 23934 20272 23940 20284
rect 23992 20272 23998 20324
rect 24504 20312 24532 20420
rect 24670 20408 24676 20420
rect 24728 20408 24734 20460
rect 24688 20380 24716 20408
rect 25225 20383 25283 20389
rect 25225 20380 25237 20383
rect 24688 20352 25237 20380
rect 25225 20349 25237 20352
rect 25271 20380 25283 20383
rect 25777 20383 25835 20389
rect 25777 20380 25789 20383
rect 25271 20352 25789 20380
rect 25271 20349 25283 20352
rect 25225 20343 25283 20349
rect 25777 20349 25789 20352
rect 25823 20349 25835 20383
rect 25777 20343 25835 20349
rect 24504 20284 25176 20312
rect 8754 20244 8760 20256
rect 8527 20216 8760 20244
rect 8527 20213 8539 20216
rect 8481 20207 8539 20213
rect 8754 20204 8760 20216
rect 8812 20244 8818 20256
rect 9582 20244 9588 20256
rect 8812 20216 9588 20244
rect 8812 20204 8818 20216
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 10042 20204 10048 20256
rect 10100 20244 10106 20256
rect 10873 20247 10931 20253
rect 10873 20244 10885 20247
rect 10100 20216 10885 20244
rect 10100 20204 10106 20216
rect 10873 20213 10885 20216
rect 10919 20213 10931 20247
rect 10873 20207 10931 20213
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 11241 20247 11299 20253
rect 11241 20244 11253 20247
rect 11112 20216 11253 20244
rect 11112 20204 11118 20216
rect 11241 20213 11253 20216
rect 11287 20213 11299 20247
rect 11606 20244 11612 20256
rect 11567 20216 11612 20244
rect 11241 20207 11299 20213
rect 11606 20204 11612 20216
rect 11664 20204 11670 20256
rect 13814 20244 13820 20256
rect 13775 20216 13820 20244
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 16758 20244 16764 20256
rect 16719 20216 16764 20244
rect 16758 20204 16764 20216
rect 16816 20204 16822 20256
rect 18782 20204 18788 20256
rect 18840 20244 18846 20256
rect 18969 20247 19027 20253
rect 18969 20244 18981 20247
rect 18840 20216 18981 20244
rect 18840 20204 18846 20216
rect 18969 20213 18981 20216
rect 19015 20244 19027 20247
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19015 20216 19625 20244
rect 19015 20213 19027 20216
rect 18969 20207 19027 20213
rect 19613 20213 19625 20216
rect 19659 20244 19671 20247
rect 20070 20244 20076 20256
rect 19659 20216 20076 20244
rect 19659 20213 19671 20216
rect 19613 20207 19671 20213
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 20806 20244 20812 20256
rect 20767 20216 20812 20244
rect 20806 20204 20812 20216
rect 20864 20204 20870 20256
rect 20898 20204 20904 20256
rect 20956 20204 20962 20256
rect 23658 20244 23664 20256
rect 23619 20216 23664 20244
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 24118 20244 24124 20256
rect 24079 20216 24124 20244
rect 24118 20204 24124 20216
rect 24176 20204 24182 20256
rect 25148 20253 25176 20284
rect 25133 20247 25191 20253
rect 25133 20213 25145 20247
rect 25179 20244 25191 20247
rect 25590 20244 25596 20256
rect 25179 20216 25596 20244
rect 25179 20213 25191 20216
rect 25133 20207 25191 20213
rect 25590 20204 25596 20216
rect 25648 20204 25654 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 1854 20040 1860 20052
rect 1627 20012 1860 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 1854 20000 1860 20012
rect 1912 20000 1918 20052
rect 2314 20000 2320 20052
rect 2372 20040 2378 20052
rect 2409 20043 2467 20049
rect 2409 20040 2421 20043
rect 2372 20012 2421 20040
rect 2372 20000 2378 20012
rect 2409 20009 2421 20012
rect 2455 20009 2467 20043
rect 2409 20003 2467 20009
rect 2774 20000 2780 20052
rect 2832 20040 2838 20052
rect 2866 20040 2872 20052
rect 2832 20012 2872 20040
rect 2832 20000 2838 20012
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 4062 20040 4068 20052
rect 4023 20012 4068 20040
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 4430 20040 4436 20052
rect 4391 20012 4436 20040
rect 4430 20000 4436 20012
rect 4488 20000 4494 20052
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 7837 20043 7895 20049
rect 7837 20040 7849 20043
rect 7064 20012 7849 20040
rect 7064 20000 7070 20012
rect 7837 20009 7849 20012
rect 7883 20009 7895 20043
rect 7837 20003 7895 20009
rect 8846 20000 8852 20052
rect 8904 20040 8910 20052
rect 8941 20043 8999 20049
rect 8941 20040 8953 20043
rect 8904 20012 8953 20040
rect 8904 20000 8910 20012
rect 8941 20009 8953 20012
rect 8987 20040 8999 20043
rect 11057 20043 11115 20049
rect 11057 20040 11069 20043
rect 8987 20012 11069 20040
rect 8987 20009 8999 20012
rect 8941 20003 8999 20009
rect 11057 20009 11069 20012
rect 11103 20009 11115 20043
rect 11057 20003 11115 20009
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 12345 20043 12403 20049
rect 12345 20040 12357 20043
rect 11204 20012 12357 20040
rect 11204 20000 11210 20012
rect 12345 20009 12357 20012
rect 12391 20009 12403 20043
rect 12345 20003 12403 20009
rect 13633 20043 13691 20049
rect 13633 20009 13645 20043
rect 13679 20040 13691 20043
rect 13722 20040 13728 20052
rect 13679 20012 13728 20040
rect 13679 20009 13691 20012
rect 13633 20003 13691 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 14645 20043 14703 20049
rect 14645 20040 14657 20043
rect 14608 20012 14657 20040
rect 14608 20000 14614 20012
rect 14645 20009 14657 20012
rect 14691 20009 14703 20043
rect 14645 20003 14703 20009
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 16301 20043 16359 20049
rect 16301 20040 16313 20043
rect 15896 20012 16313 20040
rect 15896 20000 15902 20012
rect 16301 20009 16313 20012
rect 16347 20009 16359 20043
rect 16301 20003 16359 20009
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 17221 20043 17279 20049
rect 17221 20040 17233 20043
rect 16632 20012 17233 20040
rect 16632 20000 16638 20012
rect 17221 20009 17233 20012
rect 17267 20009 17279 20043
rect 17221 20003 17279 20009
rect 17678 20000 17684 20052
rect 17736 20040 17742 20052
rect 18049 20043 18107 20049
rect 18049 20040 18061 20043
rect 17736 20012 18061 20040
rect 17736 20000 17742 20012
rect 18049 20009 18061 20012
rect 18095 20009 18107 20043
rect 18049 20003 18107 20009
rect 842 19932 848 19984
rect 900 19972 906 19984
rect 3326 19972 3332 19984
rect 900 19944 3332 19972
rect 900 19932 906 19944
rect 3326 19932 3332 19944
rect 3384 19932 3390 19984
rect 6172 19975 6230 19981
rect 6172 19941 6184 19975
rect 6218 19972 6230 19975
rect 6270 19972 6276 19984
rect 6218 19944 6276 19972
rect 6218 19941 6230 19944
rect 6172 19935 6230 19941
rect 6270 19932 6276 19944
rect 6328 19932 6334 19984
rect 7190 19932 7196 19984
rect 7248 19972 7254 19984
rect 8205 19975 8263 19981
rect 8205 19972 8217 19975
rect 7248 19944 8217 19972
rect 7248 19932 7254 19944
rect 8205 19941 8217 19944
rect 8251 19941 8263 19975
rect 8205 19935 8263 19941
rect 11701 19975 11759 19981
rect 11701 19941 11713 19975
rect 11747 19972 11759 19975
rect 12710 19972 12716 19984
rect 11747 19944 12716 19972
rect 11747 19941 11759 19944
rect 11701 19935 11759 19941
rect 12710 19932 12716 19944
rect 12768 19972 12774 19984
rect 13449 19975 13507 19981
rect 13449 19972 13461 19975
rect 12768 19944 13461 19972
rect 12768 19932 12774 19944
rect 13449 19941 13461 19944
rect 13495 19941 13507 19975
rect 13449 19935 13507 19941
rect 16761 19975 16819 19981
rect 16761 19941 16773 19975
rect 16807 19972 16819 19975
rect 16942 19972 16948 19984
rect 16807 19944 16948 19972
rect 16807 19941 16819 19944
rect 16761 19935 16819 19941
rect 16942 19932 16948 19944
rect 17000 19932 17006 19984
rect 18064 19972 18092 20003
rect 19334 20000 19340 20052
rect 19392 20040 19398 20052
rect 19705 20043 19763 20049
rect 19705 20040 19717 20043
rect 19392 20012 19717 20040
rect 19392 20000 19398 20012
rect 19705 20009 19717 20012
rect 19751 20009 19763 20043
rect 19705 20003 19763 20009
rect 20806 20000 20812 20052
rect 20864 20040 20870 20052
rect 21358 20040 21364 20052
rect 20864 20012 21364 20040
rect 20864 20000 20870 20012
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 21910 20040 21916 20052
rect 21871 20012 21916 20040
rect 21910 20000 21916 20012
rect 21968 20000 21974 20052
rect 24118 20000 24124 20052
rect 24176 20040 24182 20052
rect 24673 20043 24731 20049
rect 24673 20040 24685 20043
rect 24176 20012 24685 20040
rect 24176 20000 24182 20012
rect 24673 20009 24685 20012
rect 24719 20009 24731 20043
rect 24673 20003 24731 20009
rect 24854 20000 24860 20052
rect 24912 20040 24918 20052
rect 25225 20043 25283 20049
rect 25225 20040 25237 20043
rect 24912 20012 25237 20040
rect 24912 20000 24918 20012
rect 25225 20009 25237 20012
rect 25271 20040 25283 20043
rect 25406 20040 25412 20052
rect 25271 20012 25412 20040
rect 25271 20009 25283 20012
rect 25225 20003 25283 20009
rect 25406 20000 25412 20012
rect 25464 20000 25470 20052
rect 18064 19944 18368 19972
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2590 19904 2596 19916
rect 1443 19876 2596 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2590 19864 2596 19876
rect 2648 19864 2654 19916
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 3142 19904 3148 19916
rect 2832 19876 3148 19904
rect 2832 19864 2838 19876
rect 3142 19864 3148 19876
rect 3200 19864 3206 19916
rect 4154 19864 4160 19916
rect 4212 19904 4218 19916
rect 5077 19907 5135 19913
rect 5077 19904 5089 19907
rect 4212 19876 5089 19904
rect 4212 19864 4218 19876
rect 2314 19836 2320 19848
rect 2275 19808 2320 19836
rect 2314 19796 2320 19808
rect 2372 19796 2378 19848
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19805 3019 19839
rect 4522 19836 4528 19848
rect 4483 19808 4528 19836
rect 2961 19799 3019 19805
rect 1854 19700 1860 19712
rect 1815 19672 1860 19700
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 2976 19700 3004 19799
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 4632 19845 4660 19876
rect 5077 19873 5089 19876
rect 5123 19904 5135 19907
rect 5442 19904 5448 19916
rect 5123 19876 5448 19904
rect 5123 19873 5135 19876
rect 5077 19867 5135 19873
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 5905 19907 5963 19913
rect 5905 19873 5917 19907
rect 5951 19904 5963 19907
rect 5994 19904 6000 19916
rect 5951 19876 6000 19904
rect 5951 19873 5963 19876
rect 5905 19867 5963 19873
rect 5994 19864 6000 19876
rect 6052 19864 6058 19916
rect 8389 19907 8447 19913
rect 8389 19873 8401 19907
rect 8435 19904 8447 19907
rect 8478 19904 8484 19916
rect 8435 19876 8484 19904
rect 8435 19873 8447 19876
rect 8389 19867 8447 19873
rect 8478 19864 8484 19876
rect 8536 19864 8542 19916
rect 9306 19864 9312 19916
rect 9364 19904 9370 19916
rect 9933 19907 9991 19913
rect 9933 19904 9945 19907
rect 9364 19876 9945 19904
rect 9364 19864 9370 19876
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 6914 19728 6920 19780
rect 6972 19768 6978 19780
rect 7285 19771 7343 19777
rect 7285 19768 7297 19771
rect 6972 19740 7297 19768
rect 6972 19728 6978 19740
rect 7285 19737 7297 19740
rect 7331 19737 7343 19771
rect 7285 19731 7343 19737
rect 3697 19703 3755 19709
rect 3697 19700 3709 19703
rect 2976 19672 3709 19700
rect 3697 19669 3709 19672
rect 3743 19700 3755 19703
rect 3786 19700 3792 19712
rect 3743 19672 3792 19700
rect 3743 19669 3755 19672
rect 3697 19663 3755 19669
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 4338 19660 4344 19712
rect 4396 19700 4402 19712
rect 8573 19703 8631 19709
rect 8573 19700 8585 19703
rect 4396 19672 8585 19700
rect 4396 19660 4402 19672
rect 8573 19669 8585 19672
rect 8619 19669 8631 19703
rect 8573 19663 8631 19669
rect 9214 19660 9220 19712
rect 9272 19700 9278 19712
rect 9416 19709 9444 19876
rect 9933 19873 9945 19876
rect 9979 19873 9991 19907
rect 9933 19867 9991 19873
rect 12161 19907 12219 19913
rect 12161 19873 12173 19907
rect 12207 19904 12219 19907
rect 12250 19904 12256 19916
rect 12207 19876 12256 19904
rect 12207 19873 12219 19876
rect 12161 19867 12219 19873
rect 12250 19864 12256 19876
rect 12308 19864 12314 19916
rect 14001 19907 14059 19913
rect 14001 19873 14013 19907
rect 14047 19904 14059 19907
rect 15013 19907 15071 19913
rect 15013 19904 15025 19907
rect 14047 19876 15025 19904
rect 14047 19873 14059 19876
rect 14001 19867 14059 19873
rect 15013 19873 15025 19876
rect 15059 19873 15071 19907
rect 15013 19867 15071 19873
rect 9582 19796 9588 19848
rect 9640 19836 9646 19848
rect 9677 19839 9735 19845
rect 9677 19836 9689 19839
rect 9640 19808 9689 19836
rect 9640 19796 9646 19808
rect 9677 19805 9689 19808
rect 9723 19805 9735 19839
rect 14090 19836 14096 19848
rect 14051 19808 14096 19836
rect 9677 19799 9735 19805
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14274 19836 14280 19848
rect 14235 19808 14280 19836
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 11698 19768 11704 19780
rect 10612 19740 11704 19768
rect 9401 19703 9459 19709
rect 9401 19700 9413 19703
rect 9272 19672 9413 19700
rect 9272 19660 9278 19672
rect 9401 19669 9413 19672
rect 9447 19669 9459 19703
rect 9401 19663 9459 19669
rect 10042 19660 10048 19712
rect 10100 19700 10106 19712
rect 10612 19700 10640 19740
rect 11698 19728 11704 19740
rect 11756 19728 11762 19780
rect 12434 19768 12440 19780
rect 11992 19740 12440 19768
rect 10100 19672 10640 19700
rect 10100 19660 10106 19672
rect 11514 19660 11520 19712
rect 11572 19700 11578 19712
rect 11992 19709 12020 19740
rect 12434 19728 12440 19740
rect 12492 19728 12498 19780
rect 15028 19768 15056 19867
rect 15286 19864 15292 19916
rect 15344 19904 15350 19916
rect 15657 19907 15715 19913
rect 15657 19904 15669 19907
rect 15344 19876 15669 19904
rect 15344 19864 15350 19876
rect 15657 19873 15669 19876
rect 15703 19873 15715 19907
rect 15657 19867 15715 19873
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 17681 19907 17739 19913
rect 17681 19904 17693 19907
rect 16632 19876 17693 19904
rect 16632 19864 16638 19876
rect 17681 19873 17693 19876
rect 17727 19904 17739 19907
rect 18046 19904 18052 19916
rect 17727 19876 18052 19904
rect 17727 19873 17739 19876
rect 17681 19867 17739 19873
rect 18046 19864 18052 19876
rect 18104 19864 18110 19916
rect 18340 19913 18368 19944
rect 18598 19913 18604 19916
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19873 18383 19907
rect 18592 19904 18604 19913
rect 18559 19876 18604 19904
rect 18325 19867 18383 19873
rect 18592 19867 18604 19876
rect 18598 19864 18604 19867
rect 18656 19864 18662 19916
rect 21269 19907 21327 19913
rect 21269 19873 21281 19907
rect 21315 19904 21327 19907
rect 21542 19904 21548 19916
rect 21315 19876 21548 19904
rect 21315 19873 21327 19876
rect 21269 19867 21327 19873
rect 21542 19864 21548 19876
rect 21600 19864 21606 19916
rect 22646 19913 22652 19916
rect 22640 19904 22652 19913
rect 22607 19876 22652 19904
rect 22640 19867 22652 19876
rect 22704 19904 22710 19916
rect 24210 19904 24216 19916
rect 22704 19876 24216 19904
rect 22646 19864 22652 19867
rect 22704 19864 22710 19876
rect 24210 19864 24216 19876
rect 24268 19904 24274 19916
rect 24305 19907 24363 19913
rect 24305 19904 24317 19907
rect 24268 19876 24317 19904
rect 24268 19864 24274 19876
rect 24305 19873 24317 19876
rect 24351 19873 24363 19907
rect 24305 19867 24363 19873
rect 15470 19796 15476 19848
rect 15528 19836 15534 19848
rect 15746 19836 15752 19848
rect 15528 19808 15752 19836
rect 15528 19796 15534 19808
rect 15746 19796 15752 19808
rect 15804 19796 15810 19848
rect 15933 19839 15991 19845
rect 15933 19805 15945 19839
rect 15979 19836 15991 19839
rect 16758 19836 16764 19848
rect 15979 19808 16764 19836
rect 15979 19805 15991 19808
rect 15933 19799 15991 19805
rect 15289 19771 15347 19777
rect 15289 19768 15301 19771
rect 15028 19740 15301 19768
rect 15289 19737 15301 19740
rect 15335 19737 15347 19771
rect 15289 19731 15347 19737
rect 11977 19703 12035 19709
rect 11977 19700 11989 19703
rect 11572 19672 11989 19700
rect 11572 19660 11578 19672
rect 11977 19669 11989 19672
rect 12023 19669 12035 19703
rect 11977 19663 12035 19669
rect 12342 19660 12348 19712
rect 12400 19700 12406 19712
rect 12713 19703 12771 19709
rect 12713 19700 12725 19703
rect 12400 19672 12725 19700
rect 12400 19660 12406 19672
rect 12713 19669 12725 19672
rect 12759 19669 12771 19703
rect 12713 19663 12771 19669
rect 13173 19703 13231 19709
rect 13173 19669 13185 19703
rect 13219 19700 13231 19703
rect 13354 19700 13360 19712
rect 13219 19672 13360 19700
rect 13219 19669 13231 19672
rect 13173 19663 13231 19669
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 14826 19660 14832 19712
rect 14884 19700 14890 19712
rect 15948 19700 15976 19799
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 22278 19796 22284 19848
rect 22336 19836 22342 19848
rect 22373 19839 22431 19845
rect 22373 19836 22385 19839
rect 22336 19808 22385 19836
rect 22336 19796 22342 19808
rect 22373 19805 22385 19808
rect 22419 19805 22431 19839
rect 22373 19799 22431 19805
rect 23750 19796 23756 19848
rect 23808 19836 23814 19848
rect 24118 19836 24124 19848
rect 23808 19808 24124 19836
rect 23808 19796 23814 19808
rect 24118 19796 24124 19808
rect 24176 19796 24182 19848
rect 25314 19836 25320 19848
rect 25275 19808 25320 19836
rect 25314 19796 25320 19808
rect 25372 19796 25378 19848
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19836 25559 19839
rect 25590 19836 25596 19848
rect 25547 19808 25596 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 14884 19672 15976 19700
rect 20717 19703 20775 19709
rect 14884 19660 14890 19672
rect 20717 19669 20729 19703
rect 20763 19700 20775 19703
rect 20898 19700 20904 19712
rect 20763 19672 20904 19700
rect 20763 19669 20775 19672
rect 20717 19663 20775 19669
rect 20898 19660 20904 19672
rect 20956 19660 20962 19712
rect 21174 19700 21180 19712
rect 21135 19672 21180 19700
rect 21174 19660 21180 19672
rect 21232 19660 21238 19712
rect 21450 19700 21456 19712
rect 21411 19672 21456 19700
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 23750 19700 23756 19712
rect 23711 19672 23756 19700
rect 23750 19660 23756 19672
rect 23808 19660 23814 19712
rect 24854 19700 24860 19712
rect 24815 19672 24860 19700
rect 24854 19660 24860 19672
rect 24912 19660 24918 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 4062 19496 4068 19508
rect 2832 19468 4068 19496
rect 2832 19456 2838 19468
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 4430 19456 4436 19508
rect 4488 19496 4494 19508
rect 4617 19499 4675 19505
rect 4617 19496 4629 19499
rect 4488 19468 4629 19496
rect 4488 19456 4494 19468
rect 4617 19465 4629 19468
rect 4663 19465 4675 19499
rect 4617 19459 4675 19465
rect 4798 19456 4804 19508
rect 4856 19496 4862 19508
rect 5169 19499 5227 19505
rect 5169 19496 5181 19499
rect 4856 19468 5181 19496
rect 4856 19456 4862 19468
rect 5169 19465 5181 19468
rect 5215 19465 5227 19499
rect 5169 19459 5227 19465
rect 6086 19456 6092 19508
rect 6144 19496 6150 19508
rect 6181 19499 6239 19505
rect 6181 19496 6193 19499
rect 6144 19468 6193 19496
rect 6144 19456 6150 19468
rect 6181 19465 6193 19468
rect 6227 19465 6239 19499
rect 6181 19459 6239 19465
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10413 19499 10471 19505
rect 10413 19496 10425 19499
rect 9732 19468 10425 19496
rect 9732 19456 9738 19468
rect 10413 19465 10425 19468
rect 10459 19465 10471 19499
rect 10413 19459 10471 19465
rect 15286 19456 15292 19508
rect 15344 19496 15350 19508
rect 16485 19499 16543 19505
rect 16485 19496 16497 19499
rect 15344 19468 16497 19496
rect 15344 19456 15350 19468
rect 16485 19465 16497 19468
rect 16531 19465 16543 19499
rect 16485 19459 16543 19465
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 16853 19499 16911 19505
rect 16853 19496 16865 19499
rect 16816 19468 16865 19496
rect 16816 19456 16822 19468
rect 16853 19465 16865 19468
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 17678 19456 17684 19508
rect 17736 19496 17742 19508
rect 17773 19499 17831 19505
rect 17773 19496 17785 19499
rect 17736 19468 17785 19496
rect 17736 19456 17742 19468
rect 17773 19465 17785 19468
rect 17819 19465 17831 19499
rect 17773 19459 17831 19465
rect 2314 19388 2320 19440
rect 2372 19428 2378 19440
rect 2372 19400 3832 19428
rect 2372 19388 2378 19400
rect 3804 19372 3832 19400
rect 3878 19388 3884 19440
rect 3936 19428 3942 19440
rect 3936 19400 5212 19428
rect 3936 19388 3942 19400
rect 1854 19320 1860 19372
rect 1912 19360 1918 19372
rect 1949 19363 2007 19369
rect 1949 19360 1961 19363
rect 1912 19332 1961 19360
rect 1912 19320 1918 19332
rect 1949 19329 1961 19332
rect 1995 19329 2007 19363
rect 1949 19323 2007 19329
rect 3602 19320 3608 19372
rect 3660 19320 3666 19372
rect 3786 19320 3792 19372
rect 3844 19360 3850 19372
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 3844 19332 4261 19360
rect 3844 19320 3850 19332
rect 4249 19329 4261 19332
rect 4295 19360 4307 19363
rect 4295 19332 5120 19360
rect 4295 19329 4307 19332
rect 4249 19323 4307 19329
rect 1670 19252 1676 19304
rect 1728 19292 1734 19304
rect 1765 19295 1823 19301
rect 1765 19292 1777 19295
rect 1728 19264 1777 19292
rect 1728 19252 1734 19264
rect 1765 19261 1777 19264
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 2501 19295 2559 19301
rect 2501 19261 2513 19295
rect 2547 19292 2559 19295
rect 2774 19292 2780 19304
rect 2547 19264 2780 19292
rect 2547 19261 2559 19264
rect 2501 19255 2559 19261
rect 2774 19252 2780 19264
rect 2832 19252 2838 19304
rect 3620 19292 3648 19320
rect 3878 19292 3884 19304
rect 3620 19264 3884 19292
rect 3878 19252 3884 19264
rect 3936 19252 3942 19304
rect 3970 19252 3976 19304
rect 4028 19292 4034 19304
rect 4065 19295 4123 19301
rect 4065 19292 4077 19295
rect 4028 19264 4077 19292
rect 4028 19252 4034 19264
rect 4065 19261 4077 19264
rect 4111 19261 4123 19295
rect 4065 19255 4123 19261
rect 3513 19227 3571 19233
rect 3513 19193 3525 19227
rect 3559 19224 3571 19227
rect 3559 19196 3740 19224
rect 3559 19193 3571 19196
rect 3513 19187 3571 19193
rect 1397 19159 1455 19165
rect 1397 19125 1409 19159
rect 1443 19156 1455 19159
rect 1670 19156 1676 19168
rect 1443 19128 1676 19156
rect 1443 19125 1455 19128
rect 1397 19119 1455 19125
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 1857 19159 1915 19165
rect 1857 19125 1869 19159
rect 1903 19156 1915 19159
rect 2038 19156 2044 19168
rect 1903 19128 2044 19156
rect 1903 19125 1915 19128
rect 1857 19119 1915 19125
rect 2038 19116 2044 19128
rect 2096 19116 2102 19168
rect 3602 19156 3608 19168
rect 3563 19128 3608 19156
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 3712 19156 3740 19196
rect 3973 19159 4031 19165
rect 3973 19156 3985 19159
rect 3712 19128 3985 19156
rect 3973 19125 3985 19128
rect 4019 19156 4031 19159
rect 4614 19156 4620 19168
rect 4019 19128 4620 19156
rect 4019 19125 4031 19128
rect 3973 19119 4031 19125
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 5092 19165 5120 19332
rect 5184 19224 5212 19400
rect 11422 19388 11428 19440
rect 11480 19428 11486 19440
rect 11480 19400 13768 19428
rect 11480 19388 11486 19400
rect 5442 19320 5448 19372
rect 5500 19360 5506 19372
rect 5721 19363 5779 19369
rect 5721 19360 5733 19363
rect 5500 19332 5733 19360
rect 5500 19320 5506 19332
rect 5721 19329 5733 19332
rect 5767 19329 5779 19363
rect 5721 19323 5779 19329
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19360 7527 19363
rect 7558 19360 7564 19372
rect 7515 19332 7564 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 9030 19320 9036 19372
rect 9088 19360 9094 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 9088 19332 9413 19360
rect 9088 19320 9094 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 10134 19320 10140 19372
rect 10192 19360 10198 19372
rect 10870 19360 10876 19372
rect 10192 19332 10876 19360
rect 10192 19320 10198 19332
rect 10870 19320 10876 19332
rect 10928 19360 10934 19372
rect 10965 19363 11023 19369
rect 10965 19360 10977 19363
rect 10928 19332 10977 19360
rect 10928 19320 10934 19332
rect 10965 19329 10977 19332
rect 11011 19329 11023 19363
rect 13538 19360 13544 19372
rect 13499 19332 13544 19360
rect 10965 19323 11023 19329
rect 13538 19320 13544 19332
rect 13596 19320 13602 19372
rect 5537 19295 5595 19301
rect 5537 19261 5549 19295
rect 5583 19292 5595 19295
rect 6178 19292 6184 19304
rect 5583 19264 6184 19292
rect 5583 19261 5595 19264
rect 5537 19255 5595 19261
rect 6178 19252 6184 19264
rect 6236 19252 6242 19304
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 9309 19295 9367 19301
rect 6687 19264 7328 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 5629 19227 5687 19233
rect 5184 19196 5580 19224
rect 5077 19159 5135 19165
rect 5077 19125 5089 19159
rect 5123 19156 5135 19159
rect 5166 19156 5172 19168
rect 5123 19128 5172 19156
rect 5123 19125 5135 19128
rect 5077 19119 5135 19125
rect 5166 19116 5172 19128
rect 5224 19116 5230 19168
rect 5552 19156 5580 19196
rect 5629 19193 5641 19227
rect 5675 19224 5687 19227
rect 5675 19196 6776 19224
rect 5675 19193 5687 19196
rect 5629 19187 5687 19193
rect 6748 19168 6776 19196
rect 7300 19168 7328 19264
rect 9309 19261 9321 19295
rect 9355 19292 9367 19295
rect 9582 19292 9588 19304
rect 9355 19264 9588 19292
rect 9355 19261 9367 19264
rect 9309 19255 9367 19261
rect 9582 19252 9588 19264
rect 9640 19252 9646 19304
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 10229 19295 10287 19301
rect 10229 19292 10241 19295
rect 9824 19264 10241 19292
rect 9824 19252 9830 19264
rect 10229 19261 10241 19264
rect 10275 19292 10287 19295
rect 10781 19295 10839 19301
rect 10781 19292 10793 19295
rect 10275 19264 10793 19292
rect 10275 19261 10287 19264
rect 10229 19255 10287 19261
rect 10781 19261 10793 19264
rect 10827 19261 10839 19295
rect 11790 19292 11796 19304
rect 11751 19264 11796 19292
rect 10781 19255 10839 19261
rect 11790 19252 11796 19264
rect 11848 19252 11854 19304
rect 13357 19295 13415 19301
rect 13357 19292 13369 19295
rect 12820 19264 13369 19292
rect 12342 19224 12348 19236
rect 11440 19196 12348 19224
rect 11440 19168 11468 19196
rect 12342 19184 12348 19196
rect 12400 19184 12406 19236
rect 6086 19156 6092 19168
rect 5552 19128 6092 19156
rect 6086 19116 6092 19128
rect 6144 19116 6150 19168
rect 6730 19116 6736 19168
rect 6788 19156 6794 19168
rect 6825 19159 6883 19165
rect 6825 19156 6837 19159
rect 6788 19128 6837 19156
rect 6788 19116 6794 19128
rect 6825 19125 6837 19128
rect 6871 19125 6883 19159
rect 6825 19119 6883 19125
rect 6914 19116 6920 19168
rect 6972 19156 6978 19168
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 6972 19128 7205 19156
rect 6972 19116 6978 19128
rect 7193 19125 7205 19128
rect 7239 19125 7251 19159
rect 7193 19119 7251 19125
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 7834 19156 7840 19168
rect 7340 19128 7385 19156
rect 7795 19128 7840 19156
rect 7340 19116 7346 19128
rect 7834 19116 7840 19128
rect 7892 19116 7898 19168
rect 8481 19159 8539 19165
rect 8481 19125 8493 19159
rect 8527 19156 8539 19159
rect 8570 19156 8576 19168
rect 8527 19128 8576 19156
rect 8527 19125 8539 19128
rect 8481 19119 8539 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 8846 19156 8852 19168
rect 8807 19128 8852 19156
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 9217 19159 9275 19165
rect 9217 19125 9229 19159
rect 9263 19156 9275 19159
rect 9490 19156 9496 19168
rect 9263 19128 9496 19156
rect 9263 19125 9275 19128
rect 9217 19119 9275 19125
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 9950 19156 9956 19168
rect 9911 19128 9956 19156
rect 9950 19116 9956 19128
rect 10008 19156 10014 19168
rect 10873 19159 10931 19165
rect 10873 19156 10885 19159
rect 10008 19128 10885 19156
rect 10008 19116 10014 19128
rect 10873 19125 10885 19128
rect 10919 19125 10931 19159
rect 11422 19156 11428 19168
rect 11383 19128 11428 19156
rect 10873 19119 10931 19125
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 12250 19156 12256 19168
rect 12211 19128 12256 19156
rect 12250 19116 12256 19128
rect 12308 19116 12314 19168
rect 12526 19116 12532 19168
rect 12584 19156 12590 19168
rect 12820 19165 12848 19264
rect 13357 19261 13369 19264
rect 13403 19261 13415 19295
rect 13740 19292 13768 19400
rect 15838 19320 15844 19372
rect 15896 19320 15902 19372
rect 17034 19320 17040 19372
rect 17092 19360 17098 19372
rect 17788 19360 17816 19459
rect 20346 19456 20352 19508
rect 20404 19496 20410 19508
rect 20809 19499 20867 19505
rect 20809 19496 20821 19499
rect 20404 19468 20821 19496
rect 20404 19456 20410 19468
rect 20809 19465 20821 19468
rect 20855 19465 20867 19499
rect 20809 19459 20867 19465
rect 18049 19363 18107 19369
rect 18049 19360 18061 19363
rect 17092 19332 18061 19360
rect 17092 19320 17098 19332
rect 18049 19329 18061 19332
rect 18095 19329 18107 19363
rect 20824 19360 20852 19459
rect 25314 19456 25320 19508
rect 25372 19496 25378 19508
rect 25961 19499 26019 19505
rect 25961 19496 25973 19499
rect 25372 19468 25973 19496
rect 25372 19456 25378 19468
rect 25961 19465 25973 19468
rect 26007 19465 26019 19499
rect 25961 19459 26019 19465
rect 25590 19428 25596 19440
rect 25551 19400 25596 19428
rect 25590 19388 25596 19400
rect 25648 19388 25654 19440
rect 20990 19360 20996 19372
rect 20824 19332 20996 19360
rect 18049 19323 18107 19329
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 14182 19292 14188 19304
rect 13740 19264 14188 19292
rect 13357 19255 13415 19261
rect 14182 19252 14188 19264
rect 14240 19292 14246 19304
rect 14826 19301 14832 19304
rect 14369 19295 14427 19301
rect 14369 19292 14381 19295
rect 14240 19264 14381 19292
rect 14240 19252 14246 19264
rect 14369 19261 14381 19264
rect 14415 19292 14427 19295
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 14415 19264 14565 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 14553 19261 14565 19264
rect 14599 19261 14611 19295
rect 14820 19292 14832 19301
rect 14787 19264 14832 19292
rect 14553 19255 14611 19261
rect 14820 19255 14832 19264
rect 14826 19252 14832 19255
rect 14884 19252 14890 19304
rect 15856 19292 15884 19320
rect 15930 19292 15936 19304
rect 15856 19264 15936 19292
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 23661 19295 23719 19301
rect 23661 19261 23673 19295
rect 23707 19261 23719 19295
rect 23661 19255 23719 19261
rect 14090 19224 14096 19236
rect 13004 19196 14096 19224
rect 13004 19165 13032 19196
rect 14090 19184 14096 19196
rect 14148 19184 14154 19236
rect 14274 19224 14280 19236
rect 14187 19196 14280 19224
rect 14274 19184 14280 19196
rect 14332 19224 14338 19236
rect 18294 19227 18352 19233
rect 18294 19224 18306 19227
rect 14332 19196 14688 19224
rect 14332 19184 14338 19196
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 12584 19128 12817 19156
rect 12584 19116 12590 19128
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 12805 19119 12863 19125
rect 12989 19159 13047 19165
rect 12989 19125 13001 19159
rect 13035 19125 13047 19159
rect 12989 19119 13047 19125
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 13412 19128 13461 19156
rect 13412 19116 13418 19128
rect 13449 19125 13461 19128
rect 13495 19156 13507 19159
rect 13722 19156 13728 19168
rect 13495 19128 13728 19156
rect 13495 19125 13507 19128
rect 13449 19119 13507 19125
rect 13722 19116 13728 19128
rect 13780 19116 13786 19168
rect 14001 19159 14059 19165
rect 14001 19125 14013 19159
rect 14047 19156 14059 19159
rect 14292 19156 14320 19184
rect 14047 19128 14320 19156
rect 14047 19125 14059 19128
rect 14001 19119 14059 19125
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 14660 19156 14688 19196
rect 17420 19196 18306 19224
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 14608 19128 15945 19156
rect 14608 19116 14614 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 17420 19165 17448 19196
rect 18294 19193 18306 19196
rect 18340 19193 18352 19227
rect 18294 19187 18352 19193
rect 20533 19227 20591 19233
rect 20533 19193 20545 19227
rect 20579 19224 20591 19227
rect 21238 19227 21296 19233
rect 21238 19224 21250 19227
rect 20579 19196 21250 19224
rect 20579 19193 20591 19196
rect 20533 19187 20591 19193
rect 21238 19193 21250 19196
rect 21284 19224 21296 19227
rect 22002 19224 22008 19236
rect 21284 19196 22008 19224
rect 21284 19193 21296 19196
rect 21238 19187 21296 19193
rect 22002 19184 22008 19196
rect 22060 19184 22066 19236
rect 22278 19224 22284 19236
rect 22191 19196 22284 19224
rect 22278 19184 22284 19196
rect 22336 19224 22342 19236
rect 22925 19227 22983 19233
rect 22925 19224 22937 19227
rect 22336 19196 22937 19224
rect 22336 19184 22342 19196
rect 22925 19193 22937 19196
rect 22971 19224 22983 19227
rect 23385 19227 23443 19233
rect 23385 19224 23397 19227
rect 22971 19196 23397 19224
rect 22971 19193 22983 19196
rect 22925 19187 22983 19193
rect 23385 19193 23397 19196
rect 23431 19224 23443 19227
rect 23676 19224 23704 19255
rect 23431 19196 23704 19224
rect 23431 19193 23443 19196
rect 23385 19187 23443 19193
rect 23750 19184 23756 19236
rect 23808 19224 23814 19236
rect 23928 19227 23986 19233
rect 23928 19224 23940 19227
rect 23808 19196 23940 19224
rect 23808 19184 23814 19196
rect 23928 19193 23940 19196
rect 23974 19224 23986 19227
rect 24486 19224 24492 19236
rect 23974 19196 24492 19224
rect 23974 19193 23986 19196
rect 23928 19187 23986 19193
rect 24486 19184 24492 19196
rect 24544 19184 24550 19236
rect 17405 19159 17463 19165
rect 17405 19156 17417 19159
rect 17000 19128 17417 19156
rect 17000 19116 17006 19128
rect 17405 19125 17417 19128
rect 17451 19125 17463 19159
rect 17405 19119 17463 19125
rect 18598 19116 18604 19168
rect 18656 19156 18662 19168
rect 19429 19159 19487 19165
rect 19429 19156 19441 19159
rect 18656 19128 19441 19156
rect 18656 19116 18662 19128
rect 19429 19125 19441 19128
rect 19475 19125 19487 19159
rect 19429 19119 19487 19125
rect 20990 19116 20996 19168
rect 21048 19156 21054 19168
rect 22296 19156 22324 19184
rect 21048 19128 22324 19156
rect 22373 19159 22431 19165
rect 21048 19116 21054 19128
rect 22373 19125 22385 19159
rect 22419 19156 22431 19159
rect 23290 19156 23296 19168
rect 22419 19128 23296 19156
rect 22419 19125 22431 19128
rect 22373 19119 22431 19125
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 24026 19116 24032 19168
rect 24084 19156 24090 19168
rect 25038 19156 25044 19168
rect 24084 19128 25044 19156
rect 24084 19116 24090 19128
rect 25038 19116 25044 19128
rect 25096 19116 25102 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1397 18955 1455 18961
rect 1397 18921 1409 18955
rect 1443 18952 1455 18955
rect 1946 18952 1952 18964
rect 1443 18924 1952 18952
rect 1443 18921 1455 18924
rect 1397 18915 1455 18921
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 3697 18955 3755 18961
rect 3697 18921 3709 18955
rect 3743 18952 3755 18955
rect 3970 18952 3976 18964
rect 3743 18924 3976 18952
rect 3743 18921 3755 18924
rect 3697 18915 3755 18921
rect 3970 18912 3976 18924
rect 4028 18912 4034 18964
rect 4433 18955 4491 18961
rect 4433 18921 4445 18955
rect 4479 18952 4491 18955
rect 4982 18952 4988 18964
rect 4479 18924 4988 18952
rect 4479 18921 4491 18924
rect 4433 18915 4491 18921
rect 4982 18912 4988 18924
rect 5040 18912 5046 18964
rect 7190 18912 7196 18964
rect 7248 18952 7254 18964
rect 7377 18955 7435 18961
rect 7377 18952 7389 18955
rect 7248 18924 7389 18952
rect 7248 18912 7254 18924
rect 7377 18921 7389 18924
rect 7423 18921 7435 18955
rect 10870 18952 10876 18964
rect 10831 18924 10876 18952
rect 7377 18915 7435 18921
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 11241 18955 11299 18961
rect 11241 18952 11253 18955
rect 11112 18924 11253 18952
rect 11112 18912 11118 18924
rect 11241 18921 11253 18924
rect 11287 18921 11299 18955
rect 13814 18952 13820 18964
rect 13775 18924 13820 18952
rect 11241 18915 11299 18921
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 14185 18955 14243 18961
rect 14185 18921 14197 18955
rect 14231 18952 14243 18955
rect 15286 18952 15292 18964
rect 14231 18924 15292 18952
rect 14231 18921 14243 18924
rect 14185 18915 14243 18921
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 16850 18912 16856 18964
rect 16908 18952 16914 18964
rect 17497 18955 17555 18961
rect 17497 18952 17509 18955
rect 16908 18924 17509 18952
rect 16908 18912 16914 18924
rect 17497 18921 17509 18924
rect 17543 18921 17555 18955
rect 19058 18952 19064 18964
rect 19019 18924 19064 18952
rect 17497 18915 17555 18921
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 21818 18952 21824 18964
rect 21779 18924 21824 18952
rect 21818 18912 21824 18924
rect 21876 18912 21882 18964
rect 22278 18912 22284 18964
rect 22336 18952 22342 18964
rect 22830 18952 22836 18964
rect 22336 18924 22836 18952
rect 22336 18912 22342 18924
rect 22830 18912 22836 18924
rect 22888 18912 22894 18964
rect 23845 18955 23903 18961
rect 23845 18921 23857 18955
rect 23891 18952 23903 18955
rect 24854 18952 24860 18964
rect 23891 18924 24860 18952
rect 23891 18921 23903 18924
rect 23845 18915 23903 18921
rect 24854 18912 24860 18924
rect 24912 18912 24918 18964
rect 25133 18955 25191 18961
rect 25133 18921 25145 18955
rect 25179 18952 25191 18955
rect 25498 18952 25504 18964
rect 25179 18924 25504 18952
rect 25179 18921 25191 18924
rect 25133 18915 25191 18921
rect 25498 18912 25504 18924
rect 25556 18912 25562 18964
rect 2777 18887 2835 18893
rect 2777 18853 2789 18887
rect 2823 18884 2835 18887
rect 2958 18884 2964 18896
rect 2823 18856 2964 18884
rect 2823 18853 2835 18856
rect 2777 18847 2835 18853
rect 2958 18844 2964 18856
rect 3016 18844 3022 18896
rect 3418 18844 3424 18896
rect 3476 18884 3482 18896
rect 4798 18884 4804 18896
rect 3476 18856 4804 18884
rect 3476 18844 3482 18856
rect 4798 18844 4804 18856
rect 4856 18884 4862 18896
rect 6914 18884 6920 18896
rect 4856 18856 6920 18884
rect 4856 18844 4862 18856
rect 6914 18844 6920 18856
rect 6972 18844 6978 18896
rect 7285 18887 7343 18893
rect 7285 18853 7297 18887
rect 7331 18884 7343 18887
rect 7558 18884 7564 18896
rect 7331 18856 7564 18884
rect 7331 18853 7343 18856
rect 7285 18847 7343 18853
rect 1486 18776 1492 18828
rect 1544 18816 1550 18828
rect 4706 18816 4712 18828
rect 1544 18788 4712 18816
rect 1544 18776 1550 18788
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 5074 18776 5080 18828
rect 5132 18816 5138 18828
rect 6181 18819 6239 18825
rect 6181 18816 6193 18819
rect 5132 18788 6193 18816
rect 5132 18776 5138 18788
rect 6181 18785 6193 18788
rect 6227 18785 6239 18819
rect 6181 18779 6239 18785
rect 2866 18748 2872 18760
rect 2827 18720 2872 18748
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 2961 18751 3019 18757
rect 2961 18717 2973 18751
rect 3007 18748 3019 18751
rect 3602 18748 3608 18760
rect 3007 18720 3608 18748
rect 3007 18717 3019 18720
rect 2961 18711 3019 18717
rect 2317 18683 2375 18689
rect 2317 18649 2329 18683
rect 2363 18680 2375 18683
rect 2976 18680 3004 18711
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 4430 18708 4436 18760
rect 4488 18748 4494 18760
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 4488 18720 4537 18748
rect 4488 18708 4494 18720
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4617 18751 4675 18757
rect 4617 18717 4629 18751
rect 4663 18717 4675 18751
rect 4617 18711 4675 18717
rect 2363 18652 3004 18680
rect 2363 18649 2375 18652
rect 2317 18643 2375 18649
rect 3234 18640 3240 18692
rect 3292 18680 3298 18692
rect 4065 18683 4123 18689
rect 4065 18680 4077 18683
rect 3292 18652 4077 18680
rect 3292 18640 3298 18652
rect 4065 18649 4077 18652
rect 4111 18649 4123 18683
rect 4065 18643 4123 18649
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 3418 18612 3424 18624
rect 2455 18584 3424 18612
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 3418 18572 3424 18584
rect 3476 18572 3482 18624
rect 4522 18572 4528 18624
rect 4580 18612 4586 18624
rect 4632 18612 4660 18711
rect 6086 18708 6092 18760
rect 6144 18748 6150 18760
rect 6273 18751 6331 18757
rect 6273 18748 6285 18751
rect 6144 18720 6285 18748
rect 6144 18708 6150 18720
rect 6273 18717 6285 18720
rect 6319 18717 6331 18751
rect 6273 18711 6331 18717
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18748 6515 18751
rect 7098 18748 7104 18760
rect 6503 18720 7104 18748
rect 6503 18717 6515 18720
rect 6457 18711 6515 18717
rect 5166 18680 5172 18692
rect 5079 18652 5172 18680
rect 5166 18640 5172 18652
rect 5224 18680 5230 18692
rect 5721 18683 5779 18689
rect 5721 18680 5733 18683
rect 5224 18652 5733 18680
rect 5224 18640 5230 18652
rect 5721 18649 5733 18652
rect 5767 18680 5779 18683
rect 6472 18680 6500 18711
rect 7098 18708 7104 18720
rect 7156 18748 7162 18760
rect 7300 18748 7328 18847
rect 7558 18844 7564 18856
rect 7616 18884 7622 18896
rect 13630 18884 13636 18896
rect 7616 18856 7972 18884
rect 7616 18844 7622 18856
rect 7745 18819 7803 18825
rect 7745 18816 7757 18819
rect 7156 18720 7328 18748
rect 7392 18788 7757 18816
rect 7156 18708 7162 18720
rect 5767 18652 6500 18680
rect 5767 18649 5779 18652
rect 5721 18643 5779 18649
rect 7282 18640 7288 18692
rect 7340 18680 7346 18692
rect 7392 18680 7420 18788
rect 7745 18785 7757 18788
rect 7791 18785 7803 18819
rect 7745 18779 7803 18785
rect 7834 18748 7840 18760
rect 7795 18720 7840 18748
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 7944 18757 7972 18856
rect 12443 18856 13636 18884
rect 10226 18816 10232 18828
rect 10187 18788 10232 18816
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 11330 18776 11336 18828
rect 11388 18816 11394 18828
rect 11692 18819 11750 18825
rect 11692 18816 11704 18819
rect 11388 18788 11704 18816
rect 11388 18776 11394 18788
rect 11692 18785 11704 18788
rect 11738 18816 11750 18819
rect 12443 18816 12471 18856
rect 13630 18844 13636 18856
rect 13688 18844 13694 18896
rect 14090 18844 14096 18896
rect 14148 18884 14154 18896
rect 15013 18887 15071 18893
rect 15013 18884 15025 18887
rect 14148 18856 15025 18884
rect 14148 18844 14154 18856
rect 15013 18853 15025 18856
rect 15059 18853 15071 18887
rect 15013 18847 15071 18853
rect 17221 18887 17279 18893
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 17957 18887 18015 18893
rect 17957 18884 17969 18887
rect 17267 18856 17969 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 17957 18853 17969 18856
rect 18003 18853 18015 18887
rect 17957 18847 18015 18853
rect 18690 18844 18696 18896
rect 18748 18884 18754 18896
rect 19150 18884 19156 18896
rect 18748 18856 19156 18884
rect 18748 18844 18754 18856
rect 19150 18844 19156 18856
rect 19208 18884 19214 18896
rect 19521 18887 19579 18893
rect 19521 18884 19533 18887
rect 19208 18856 19533 18884
rect 19208 18844 19214 18856
rect 19521 18853 19533 18856
rect 19567 18853 19579 18887
rect 19521 18847 19579 18853
rect 21729 18887 21787 18893
rect 21729 18853 21741 18887
rect 21775 18884 21787 18887
rect 22646 18884 22652 18896
rect 21775 18856 22652 18884
rect 21775 18853 21787 18856
rect 21729 18847 21787 18853
rect 11738 18788 12471 18816
rect 13449 18819 13507 18825
rect 11738 18785 11750 18788
rect 11692 18779 11750 18785
rect 13449 18785 13461 18819
rect 13495 18816 13507 18819
rect 13538 18816 13544 18828
rect 13495 18788 13544 18816
rect 13495 18785 13507 18788
rect 13449 18779 13507 18785
rect 13538 18776 13544 18788
rect 13596 18816 13602 18828
rect 14737 18819 14795 18825
rect 14737 18816 14749 18819
rect 13596 18788 14749 18816
rect 13596 18776 13602 18788
rect 14737 18785 14749 18788
rect 14783 18816 14795 18819
rect 14826 18816 14832 18828
rect 14783 18788 14832 18816
rect 14783 18785 14795 18788
rect 14737 18779 14795 18785
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 16298 18816 16304 18828
rect 16259 18788 16304 18816
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 17865 18819 17923 18825
rect 17865 18785 17877 18819
rect 17911 18785 17923 18819
rect 17865 18779 17923 18785
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18717 7987 18751
rect 7929 18711 7987 18717
rect 8846 18708 8852 18760
rect 8904 18748 8910 18760
rect 10318 18748 10324 18760
rect 8904 18720 10324 18748
rect 8904 18708 8910 18720
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 10502 18748 10508 18760
rect 10463 18720 10508 18748
rect 10502 18708 10508 18720
rect 10560 18708 10566 18760
rect 11422 18748 11428 18760
rect 11383 18720 11428 18748
rect 11422 18708 11428 18720
rect 11480 18708 11486 18760
rect 16390 18748 16396 18760
rect 16351 18720 16396 18748
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 16850 18748 16856 18760
rect 16623 18720 16856 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 7340 18652 7420 18680
rect 9493 18683 9551 18689
rect 7340 18640 7346 18652
rect 9493 18649 9505 18683
rect 9539 18680 9551 18683
rect 9674 18680 9680 18692
rect 9539 18652 9680 18680
rect 9539 18649 9551 18652
rect 9493 18643 9551 18649
rect 9674 18640 9680 18652
rect 9732 18680 9738 18692
rect 10520 18680 10548 18708
rect 9732 18652 10548 18680
rect 15933 18683 15991 18689
rect 9732 18640 9738 18652
rect 15933 18649 15945 18683
rect 15979 18680 15991 18683
rect 16945 18683 17003 18689
rect 16945 18680 16957 18683
rect 15979 18652 16957 18680
rect 15979 18649 15991 18652
rect 15933 18643 15991 18649
rect 16945 18649 16957 18652
rect 16991 18680 17003 18683
rect 17880 18680 17908 18779
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 19116 18788 19441 18816
rect 19116 18776 19122 18788
rect 19429 18785 19441 18788
rect 19475 18785 19487 18819
rect 19429 18779 19487 18785
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 22189 18819 22247 18825
rect 22189 18816 22201 18819
rect 21876 18788 22201 18816
rect 21876 18776 21882 18788
rect 22189 18785 22201 18788
rect 22235 18785 22247 18819
rect 22189 18779 22247 18785
rect 18046 18748 18052 18760
rect 18007 18720 18052 18748
rect 18046 18708 18052 18720
rect 18104 18748 18110 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 18104 18720 18521 18748
rect 18104 18708 18110 18720
rect 18509 18717 18521 18720
rect 18555 18748 18567 18751
rect 18598 18748 18604 18760
rect 18555 18720 18604 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 22278 18748 22284 18760
rect 22239 18720 22284 18748
rect 19613 18711 19671 18717
rect 16991 18652 17908 18680
rect 16991 18649 17003 18652
rect 16945 18643 17003 18649
rect 19334 18640 19340 18692
rect 19392 18680 19398 18692
rect 19628 18680 19656 18711
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 22388 18757 22416 18856
rect 22646 18844 22652 18856
rect 22704 18884 22710 18896
rect 23201 18887 23259 18893
rect 23201 18884 23213 18887
rect 22704 18856 23213 18884
rect 22704 18844 22710 18856
rect 23201 18853 23213 18856
rect 23247 18853 23259 18887
rect 24486 18884 24492 18896
rect 24399 18856 24492 18884
rect 23201 18847 23259 18853
rect 24486 18844 24492 18856
rect 24544 18884 24550 18896
rect 25590 18884 25596 18896
rect 24544 18856 25596 18884
rect 24544 18844 24550 18856
rect 25590 18844 25596 18856
rect 25648 18844 25654 18896
rect 23750 18816 23756 18828
rect 23711 18788 23756 18816
rect 23750 18776 23756 18788
rect 23808 18776 23814 18828
rect 24949 18819 25007 18825
rect 24949 18785 24961 18819
rect 24995 18785 25007 18819
rect 24949 18779 25007 18785
rect 22373 18751 22431 18757
rect 22373 18717 22385 18751
rect 22419 18717 22431 18751
rect 23934 18748 23940 18760
rect 23895 18720 23940 18748
rect 22373 18711 22431 18717
rect 23934 18708 23940 18720
rect 23992 18708 23998 18760
rect 24964 18748 24992 18779
rect 25406 18776 25412 18828
rect 25464 18816 25470 18828
rect 25501 18819 25559 18825
rect 25501 18816 25513 18819
rect 25464 18788 25513 18816
rect 25464 18776 25470 18788
rect 25501 18785 25513 18788
rect 25547 18785 25559 18819
rect 25501 18779 25559 18785
rect 25590 18748 25596 18760
rect 24964 18720 25596 18748
rect 25590 18708 25596 18720
rect 25648 18708 25654 18760
rect 19392 18652 19656 18680
rect 19392 18640 19398 18652
rect 5184 18612 5212 18640
rect 4580 18584 5212 18612
rect 5813 18615 5871 18621
rect 4580 18572 4586 18584
rect 5813 18581 5825 18615
rect 5859 18612 5871 18615
rect 6178 18612 6184 18624
rect 5859 18584 6184 18612
rect 5859 18581 5871 18584
rect 5813 18575 5871 18581
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 8478 18612 8484 18624
rect 8391 18584 8484 18612
rect 8478 18572 8484 18584
rect 8536 18612 8542 18624
rect 8941 18615 8999 18621
rect 8941 18612 8953 18615
rect 8536 18584 8953 18612
rect 8536 18572 8542 18584
rect 8941 18581 8953 18584
rect 8987 18612 8999 18615
rect 9030 18612 9036 18624
rect 8987 18584 9036 18612
rect 8987 18581 8999 18584
rect 8941 18575 8999 18581
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 9858 18612 9864 18624
rect 9819 18584 9864 18612
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 12158 18572 12164 18624
rect 12216 18612 12222 18624
rect 12805 18615 12863 18621
rect 12805 18612 12817 18615
rect 12216 18584 12817 18612
rect 12216 18572 12222 18584
rect 12805 18581 12817 18584
rect 12851 18581 12863 18615
rect 15470 18612 15476 18624
rect 15431 18584 15476 18612
rect 12805 18575 12863 18581
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 17221 18615 17279 18621
rect 17221 18612 17233 18615
rect 16632 18584 17233 18612
rect 16632 18572 16638 18584
rect 17221 18581 17233 18584
rect 17267 18612 17279 18615
rect 17313 18615 17371 18621
rect 17313 18612 17325 18615
rect 17267 18584 17325 18612
rect 17267 18581 17279 18584
rect 17221 18575 17279 18581
rect 17313 18581 17325 18584
rect 17359 18581 17371 18615
rect 17313 18575 17371 18581
rect 19518 18572 19524 18624
rect 19576 18612 19582 18624
rect 20073 18615 20131 18621
rect 20073 18612 20085 18615
rect 19576 18584 20085 18612
rect 19576 18572 19582 18584
rect 20073 18581 20085 18584
rect 20119 18612 20131 18615
rect 20622 18612 20628 18624
rect 20119 18584 20628 18612
rect 20119 18581 20131 18584
rect 20073 18575 20131 18581
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 21361 18615 21419 18621
rect 21361 18581 21373 18615
rect 21407 18612 21419 18615
rect 21542 18612 21548 18624
rect 21407 18584 21548 18612
rect 21407 18581 21419 18584
rect 21361 18575 21419 18581
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 22830 18612 22836 18624
rect 22791 18584 22836 18612
rect 22830 18572 22836 18584
rect 22888 18572 22894 18624
rect 23385 18615 23443 18621
rect 23385 18581 23397 18615
rect 23431 18612 23443 18615
rect 23566 18612 23572 18624
rect 23431 18584 23572 18612
rect 23431 18581 23443 18584
rect 23385 18575 23443 18581
rect 23566 18572 23572 18584
rect 23624 18572 23630 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2958 18408 2964 18420
rect 2919 18380 2964 18408
rect 2958 18368 2964 18380
rect 3016 18368 3022 18420
rect 3786 18368 3792 18420
rect 3844 18408 3850 18420
rect 5074 18408 5080 18420
rect 3844 18380 5080 18408
rect 3844 18368 3850 18380
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 6641 18411 6699 18417
rect 6641 18377 6653 18411
rect 6687 18408 6699 18411
rect 7742 18408 7748 18420
rect 6687 18380 7748 18408
rect 6687 18377 6699 18380
rect 6641 18371 6699 18377
rect 7742 18368 7748 18380
rect 7800 18368 7806 18420
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 11793 18411 11851 18417
rect 11793 18408 11805 18411
rect 8444 18380 11805 18408
rect 8444 18368 8450 18380
rect 11793 18377 11805 18380
rect 11839 18408 11851 18411
rect 11977 18411 12035 18417
rect 11977 18408 11989 18411
rect 11839 18380 11989 18408
rect 11839 18377 11851 18380
rect 11793 18371 11851 18377
rect 11977 18377 11989 18380
rect 12023 18377 12035 18411
rect 12618 18408 12624 18420
rect 11977 18371 12035 18377
rect 12176 18380 12624 18408
rect 4522 18340 4528 18352
rect 4483 18312 4528 18340
rect 4522 18300 4528 18312
rect 4580 18300 4586 18352
rect 5537 18343 5595 18349
rect 5537 18309 5549 18343
rect 5583 18340 5595 18343
rect 6086 18340 6092 18352
rect 5583 18312 6092 18340
rect 5583 18309 5595 18312
rect 5537 18303 5595 18309
rect 6086 18300 6092 18312
rect 6144 18300 6150 18352
rect 7834 18340 7840 18352
rect 7795 18312 7840 18340
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 1946 18232 1952 18284
rect 2004 18272 2010 18284
rect 2041 18275 2099 18281
rect 2041 18272 2053 18275
rect 2004 18244 2053 18272
rect 2004 18232 2010 18244
rect 2041 18241 2053 18244
rect 2087 18272 2099 18275
rect 8478 18272 8484 18284
rect 2087 18244 3280 18272
rect 8439 18244 8484 18272
rect 2087 18241 2099 18244
rect 2041 18235 2099 18241
rect 2958 18164 2964 18216
rect 3016 18204 3022 18216
rect 3145 18207 3203 18213
rect 3145 18204 3157 18207
rect 3016 18176 3157 18204
rect 3016 18164 3022 18176
rect 3145 18173 3157 18176
rect 3191 18173 3203 18207
rect 3252 18204 3280 18244
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 3401 18207 3459 18213
rect 3401 18204 3413 18207
rect 3252 18176 3413 18204
rect 3145 18167 3203 18173
rect 3401 18173 3413 18176
rect 3447 18204 3459 18207
rect 3786 18204 3792 18216
rect 3447 18176 3792 18204
rect 3447 18173 3459 18176
rect 3401 18167 3459 18173
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 4706 18164 4712 18216
rect 4764 18204 4770 18216
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 4764 18176 5641 18204
rect 4764 18164 4770 18176
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 1670 18096 1676 18148
rect 1728 18136 1734 18148
rect 1857 18139 1915 18145
rect 1857 18136 1869 18139
rect 1728 18108 1869 18136
rect 1728 18096 1734 18108
rect 1857 18105 1869 18108
rect 1903 18136 1915 18139
rect 2593 18139 2651 18145
rect 1903 18108 2544 18136
rect 1903 18105 1915 18108
rect 1857 18099 1915 18105
rect 1394 18028 1400 18080
rect 1452 18068 1458 18080
rect 1489 18071 1547 18077
rect 1489 18068 1501 18071
rect 1452 18040 1501 18068
rect 1452 18028 1458 18040
rect 1489 18037 1501 18040
rect 1535 18037 1547 18071
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1489 18031 1547 18037
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2516 18068 2544 18108
rect 2593 18105 2605 18139
rect 2639 18136 2651 18139
rect 2866 18136 2872 18148
rect 2639 18108 2872 18136
rect 2639 18105 2651 18108
rect 2593 18099 2651 18105
rect 2866 18096 2872 18108
rect 2924 18136 2930 18148
rect 4246 18136 4252 18148
rect 2924 18108 4252 18136
rect 2924 18096 2930 18108
rect 4246 18096 4252 18108
rect 4304 18096 4310 18148
rect 5644 18136 5672 18167
rect 8202 18164 8208 18216
rect 8260 18204 8266 18216
rect 8297 18207 8355 18213
rect 8297 18204 8309 18207
rect 8260 18176 8309 18204
rect 8260 18164 8266 18176
rect 8297 18173 8309 18176
rect 8343 18173 8355 18207
rect 8297 18167 8355 18173
rect 8754 18164 8760 18216
rect 8812 18164 8818 18216
rect 9674 18213 9680 18216
rect 9401 18207 9459 18213
rect 9401 18173 9413 18207
rect 9447 18173 9459 18207
rect 9668 18204 9680 18213
rect 9635 18176 9680 18204
rect 9401 18167 9459 18173
rect 9668 18167 9680 18176
rect 6273 18139 6331 18145
rect 6273 18136 6285 18139
rect 5644 18108 6285 18136
rect 6273 18105 6285 18108
rect 6319 18136 6331 18139
rect 7190 18136 7196 18148
rect 6319 18108 7196 18136
rect 6319 18105 6331 18108
rect 6273 18099 6331 18105
rect 7190 18096 7196 18108
rect 7248 18096 7254 18148
rect 7742 18096 7748 18148
rect 7800 18136 7806 18148
rect 8772 18136 8800 18164
rect 9217 18139 9275 18145
rect 9217 18136 9229 18139
rect 7800 18108 9229 18136
rect 7800 18096 7806 18108
rect 9217 18105 9229 18108
rect 9263 18136 9275 18139
rect 9416 18136 9444 18167
rect 9674 18164 9680 18167
rect 9732 18164 9738 18216
rect 9263 18108 9444 18136
rect 9263 18105 9275 18108
rect 9217 18099 9275 18105
rect 11054 18096 11060 18148
rect 11112 18136 11118 18148
rect 12176 18145 12204 18380
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 14182 18408 14188 18420
rect 14143 18380 14188 18408
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 16298 18368 16304 18420
rect 16356 18408 16362 18420
rect 16577 18411 16635 18417
rect 16577 18408 16589 18411
rect 16356 18380 16589 18408
rect 16356 18368 16362 18380
rect 16577 18377 16589 18380
rect 16623 18377 16635 18411
rect 16577 18371 16635 18377
rect 17589 18411 17647 18417
rect 17589 18377 17601 18411
rect 17635 18408 17647 18411
rect 18046 18408 18052 18420
rect 17635 18380 18052 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 12897 18275 12955 18281
rect 12897 18272 12909 18275
rect 12268 18244 12909 18272
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 11112 18108 12173 18136
rect 11112 18096 11118 18108
rect 12161 18105 12173 18108
rect 12207 18105 12219 18139
rect 12161 18099 12219 18105
rect 5166 18068 5172 18080
rect 2516 18040 5172 18068
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 5810 18068 5816 18080
rect 5771 18040 5816 18068
rect 5810 18028 5816 18040
rect 5868 18028 5874 18080
rect 6638 18028 6644 18080
rect 6696 18068 6702 18080
rect 6825 18071 6883 18077
rect 6825 18068 6837 18071
rect 6696 18040 6837 18068
rect 6696 18028 6702 18040
rect 6825 18037 6837 18040
rect 6871 18037 6883 18071
rect 6825 18031 6883 18037
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 7377 18071 7435 18077
rect 7377 18068 7389 18071
rect 7340 18040 7389 18068
rect 7340 18028 7346 18040
rect 7377 18037 7389 18040
rect 7423 18037 7435 18071
rect 7377 18031 7435 18037
rect 8205 18071 8263 18077
rect 8205 18037 8217 18071
rect 8251 18068 8263 18071
rect 8754 18068 8760 18080
rect 8251 18040 8760 18068
rect 8251 18037 8263 18040
rect 8205 18031 8263 18037
rect 8754 18028 8760 18040
rect 8812 18068 8818 18080
rect 8849 18071 8907 18077
rect 8849 18068 8861 18071
rect 8812 18040 8861 18068
rect 8812 18028 8818 18040
rect 8849 18037 8861 18040
rect 8895 18037 8907 18071
rect 8849 18031 8907 18037
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 10781 18071 10839 18077
rect 10781 18068 10793 18071
rect 9732 18040 10793 18068
rect 9732 18028 9738 18040
rect 10781 18037 10793 18040
rect 10827 18037 10839 18071
rect 10781 18031 10839 18037
rect 11422 18028 11428 18080
rect 11480 18068 11486 18080
rect 11517 18071 11575 18077
rect 11517 18068 11529 18071
rect 11480 18040 11529 18068
rect 11480 18028 11486 18040
rect 11517 18037 11529 18040
rect 11563 18068 11575 18071
rect 11790 18068 11796 18080
rect 11563 18040 11796 18068
rect 11563 18037 11575 18040
rect 11517 18031 11575 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 11977 18071 12035 18077
rect 11977 18037 11989 18071
rect 12023 18068 12035 18071
rect 12268 18068 12296 18244
rect 12897 18241 12909 18244
rect 12943 18241 12955 18275
rect 12897 18235 12955 18241
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18272 13139 18275
rect 13446 18272 13452 18284
rect 13127 18244 13452 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 13446 18232 13452 18244
rect 13504 18232 13510 18284
rect 13630 18232 13636 18284
rect 13688 18272 13694 18284
rect 14200 18272 14228 18368
rect 14277 18275 14335 18281
rect 14277 18272 14289 18275
rect 13688 18244 14289 18272
rect 13688 18232 13694 18244
rect 14277 18241 14289 18244
rect 14323 18241 14335 18275
rect 16592 18272 16620 18371
rect 18046 18368 18052 18380
rect 18104 18368 18110 18420
rect 18417 18411 18475 18417
rect 18417 18377 18429 18411
rect 18463 18408 18475 18411
rect 19334 18408 19340 18420
rect 18463 18380 19340 18408
rect 18463 18377 18475 18380
rect 18417 18371 18475 18377
rect 19334 18368 19340 18380
rect 19392 18368 19398 18420
rect 23474 18408 23480 18420
rect 23435 18380 23480 18408
rect 23474 18368 23480 18380
rect 23532 18408 23538 18420
rect 23532 18380 24164 18408
rect 23532 18368 23538 18380
rect 16945 18275 17003 18281
rect 16945 18272 16957 18275
rect 16592 18244 16957 18272
rect 14277 18235 14335 18241
rect 16945 18241 16957 18244
rect 16991 18241 17003 18275
rect 16945 18235 17003 18241
rect 22649 18275 22707 18281
rect 22649 18241 22661 18275
rect 22695 18272 22707 18275
rect 22830 18272 22836 18284
rect 22695 18244 22836 18272
rect 22695 18241 22707 18244
rect 22649 18235 22707 18241
rect 22830 18232 22836 18244
rect 22888 18232 22894 18284
rect 24136 18281 24164 18380
rect 24854 18368 24860 18420
rect 24912 18408 24918 18420
rect 25409 18411 25467 18417
rect 25409 18408 25421 18411
rect 24912 18380 25421 18408
rect 24912 18368 24918 18380
rect 25409 18377 25421 18380
rect 25455 18377 25467 18411
rect 26234 18408 26240 18420
rect 26195 18380 26240 18408
rect 25409 18371 25467 18377
rect 26234 18368 26240 18380
rect 26292 18368 26298 18420
rect 25038 18340 25044 18352
rect 24999 18312 25044 18340
rect 25038 18300 25044 18312
rect 25096 18300 25102 18352
rect 24121 18275 24179 18281
rect 24121 18241 24133 18275
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 24210 18232 24216 18284
rect 24268 18272 24274 18284
rect 24268 18244 24313 18272
rect 24268 18232 24274 18244
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 14550 18213 14556 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12676 18176 12817 18204
rect 12676 18164 12682 18176
rect 12805 18173 12817 18176
rect 12851 18173 12863 18207
rect 14544 18204 14556 18213
rect 14511 18176 14556 18204
rect 12805 18167 12863 18173
rect 14544 18167 14556 18176
rect 14550 18164 14556 18167
rect 14608 18164 14614 18216
rect 19242 18164 19248 18216
rect 19300 18204 19306 18216
rect 19521 18207 19579 18213
rect 19521 18204 19533 18207
rect 19300 18176 19533 18204
rect 19300 18164 19306 18176
rect 19521 18173 19533 18176
rect 19567 18173 19579 18207
rect 19521 18167 19579 18173
rect 22373 18207 22431 18213
rect 22373 18173 22385 18207
rect 22419 18204 22431 18207
rect 22462 18204 22468 18216
rect 22419 18176 22468 18204
rect 22419 18173 22431 18176
rect 22373 18167 22431 18173
rect 22462 18164 22468 18176
rect 22520 18164 22526 18216
rect 23658 18164 23664 18216
rect 23716 18204 23722 18216
rect 24029 18207 24087 18213
rect 24029 18204 24041 18207
rect 23716 18176 24041 18204
rect 23716 18164 23722 18176
rect 24029 18173 24041 18176
rect 24075 18204 24087 18207
rect 24673 18207 24731 18213
rect 24673 18204 24685 18207
rect 24075 18176 24685 18204
rect 24075 18173 24087 18176
rect 24029 18167 24087 18173
rect 24673 18173 24685 18176
rect 24719 18173 24731 18207
rect 25222 18204 25228 18216
rect 25135 18176 25228 18204
rect 24673 18167 24731 18173
rect 25222 18164 25228 18176
rect 25280 18204 25286 18216
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25280 18176 25789 18204
rect 25280 18164 25286 18176
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 15562 18096 15568 18148
rect 15620 18136 15626 18148
rect 16209 18139 16267 18145
rect 16209 18136 16221 18139
rect 15620 18108 16221 18136
rect 15620 18096 15626 18108
rect 16209 18105 16221 18108
rect 16255 18136 16267 18139
rect 16390 18136 16396 18148
rect 16255 18108 16396 18136
rect 16255 18105 16267 18108
rect 16209 18099 16267 18105
rect 16390 18096 16396 18108
rect 16448 18096 16454 18148
rect 19766 18139 19824 18145
rect 19766 18136 19778 18139
rect 19536 18108 19778 18136
rect 19536 18080 19564 18108
rect 19766 18105 19778 18108
rect 19812 18105 19824 18139
rect 19766 18099 19824 18105
rect 21545 18139 21603 18145
rect 21545 18105 21557 18139
rect 21591 18136 21603 18139
rect 22278 18136 22284 18148
rect 21591 18108 22284 18136
rect 21591 18105 21603 18108
rect 21545 18099 21603 18105
rect 22278 18096 22284 18108
rect 22336 18096 22342 18148
rect 12023 18040 12296 18068
rect 12023 18037 12035 18040
rect 11977 18031 12035 18037
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12492 18040 12537 18068
rect 12492 18028 12498 18040
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 15657 18071 15715 18077
rect 15657 18068 15669 18071
rect 15344 18040 15669 18068
rect 15344 18028 15350 18040
rect 15657 18037 15669 18040
rect 15703 18037 15715 18071
rect 18506 18068 18512 18080
rect 18467 18040 18512 18068
rect 15657 18031 15715 18037
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 19058 18068 19064 18080
rect 19019 18040 19064 18068
rect 19058 18028 19064 18040
rect 19116 18028 19122 18080
rect 19518 18028 19524 18080
rect 19576 18028 19582 18080
rect 20901 18071 20959 18077
rect 20901 18037 20913 18071
rect 20947 18068 20959 18071
rect 21450 18068 21456 18080
rect 20947 18040 21456 18068
rect 20947 18037 20959 18040
rect 20901 18031 20959 18037
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 21818 18068 21824 18080
rect 21779 18040 21824 18068
rect 21818 18028 21824 18040
rect 21876 18028 21882 18080
rect 22002 18068 22008 18080
rect 21963 18040 22008 18068
rect 22002 18028 22008 18040
rect 22060 18028 22066 18080
rect 22465 18071 22523 18077
rect 22465 18037 22477 18071
rect 22511 18068 22523 18071
rect 23017 18071 23075 18077
rect 23017 18068 23029 18071
rect 22511 18040 23029 18068
rect 22511 18037 22523 18040
rect 22465 18031 22523 18037
rect 23017 18037 23029 18040
rect 23063 18068 23075 18071
rect 23290 18068 23296 18080
rect 23063 18040 23296 18068
rect 23063 18037 23075 18040
rect 23017 18031 23075 18037
rect 23290 18028 23296 18040
rect 23348 18028 23354 18080
rect 23658 18068 23664 18080
rect 23619 18040 23664 18068
rect 23658 18028 23664 18040
rect 23716 18028 23722 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1854 17824 1860 17876
rect 1912 17864 1918 17876
rect 2314 17864 2320 17876
rect 1912 17836 2320 17864
rect 1912 17824 1918 17836
rect 2314 17824 2320 17836
rect 2372 17864 2378 17876
rect 2869 17867 2927 17873
rect 2869 17864 2881 17867
rect 2372 17836 2881 17864
rect 2372 17824 2378 17836
rect 2869 17833 2881 17836
rect 2915 17833 2927 17867
rect 3786 17864 3792 17876
rect 3747 17836 3792 17864
rect 2869 17827 2927 17833
rect 3786 17824 3792 17836
rect 3844 17824 3850 17876
rect 4709 17867 4767 17873
rect 4709 17833 4721 17867
rect 4755 17864 4767 17867
rect 4982 17864 4988 17876
rect 4755 17836 4988 17864
rect 4755 17833 4767 17836
rect 4709 17827 4767 17833
rect 4982 17824 4988 17836
rect 5040 17824 5046 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6733 17867 6791 17873
rect 6733 17864 6745 17867
rect 5592 17836 6745 17864
rect 5592 17824 5598 17836
rect 6733 17833 6745 17836
rect 6779 17833 6791 17867
rect 7098 17864 7104 17876
rect 7059 17836 7104 17864
rect 6733 17827 6791 17833
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 9493 17867 9551 17873
rect 9493 17833 9505 17867
rect 9539 17864 9551 17867
rect 9582 17864 9588 17876
rect 9539 17836 9588 17864
rect 9539 17833 9551 17836
rect 9493 17827 9551 17833
rect 9582 17824 9588 17836
rect 9640 17824 9646 17876
rect 10778 17864 10784 17876
rect 10739 17836 10784 17864
rect 10778 17824 10784 17836
rect 10836 17824 10842 17876
rect 10870 17824 10876 17876
rect 10928 17864 10934 17876
rect 11330 17864 11336 17876
rect 10928 17836 11336 17864
rect 10928 17824 10934 17836
rect 11330 17824 11336 17836
rect 11388 17824 11394 17876
rect 12802 17864 12808 17876
rect 12763 17836 12808 17864
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 13814 17864 13820 17876
rect 13775 17836 13820 17864
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 14550 17824 14556 17876
rect 14608 17864 14614 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14608 17836 14657 17864
rect 14608 17824 14614 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 19150 17864 19156 17876
rect 19111 17836 19156 17864
rect 14645 17827 14703 17833
rect 19150 17824 19156 17836
rect 19208 17824 19214 17876
rect 19889 17867 19947 17873
rect 19889 17833 19901 17867
rect 19935 17864 19947 17867
rect 19978 17864 19984 17876
rect 19935 17836 19984 17864
rect 19935 17833 19947 17836
rect 19889 17827 19947 17833
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22281 17867 22339 17873
rect 22281 17864 22293 17867
rect 22152 17836 22293 17864
rect 22152 17824 22158 17836
rect 22281 17833 22293 17836
rect 22327 17833 22339 17867
rect 22281 17827 22339 17833
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 22833 17867 22891 17873
rect 22833 17864 22845 17867
rect 22520 17836 22845 17864
rect 22520 17824 22526 17836
rect 22833 17833 22845 17836
rect 22879 17833 22891 17867
rect 22833 17827 22891 17833
rect 1756 17799 1814 17805
rect 1756 17765 1768 17799
rect 1802 17796 1814 17799
rect 2222 17796 2228 17808
rect 1802 17768 2228 17796
rect 1802 17765 1814 17768
rect 1756 17759 1814 17765
rect 2222 17756 2228 17768
rect 2280 17756 2286 17808
rect 6914 17756 6920 17808
rect 6972 17796 6978 17808
rect 7745 17799 7803 17805
rect 7745 17796 7757 17799
rect 6972 17768 7757 17796
rect 6972 17756 6978 17768
rect 7745 17765 7757 17768
rect 7791 17796 7803 17799
rect 7834 17796 7840 17808
rect 7791 17768 7840 17796
rect 7791 17765 7803 17768
rect 7745 17759 7803 17765
rect 7834 17756 7840 17768
rect 7892 17756 7898 17808
rect 9306 17756 9312 17808
rect 9364 17796 9370 17808
rect 10045 17799 10103 17805
rect 10045 17796 10057 17799
rect 9364 17768 10057 17796
rect 9364 17756 9370 17768
rect 10045 17765 10057 17768
rect 10091 17765 10103 17799
rect 13354 17796 13360 17808
rect 13315 17768 13360 17796
rect 10045 17759 10103 17765
rect 13354 17756 13360 17768
rect 13412 17756 13418 17808
rect 17212 17799 17270 17805
rect 17212 17796 17224 17799
rect 16040 17768 17224 17796
rect 2958 17728 2964 17740
rect 1504 17700 2964 17728
rect 1504 17672 1532 17700
rect 2958 17688 2964 17700
rect 3016 17728 3022 17740
rect 3421 17731 3479 17737
rect 3421 17728 3433 17731
rect 3016 17700 3433 17728
rect 3016 17688 3022 17700
rect 3421 17697 3433 17700
rect 3467 17728 3479 17731
rect 3970 17728 3976 17740
rect 3467 17700 3976 17728
rect 3467 17697 3479 17700
rect 3421 17691 3479 17697
rect 3970 17688 3976 17700
rect 4028 17688 4034 17740
rect 4062 17688 4068 17740
rect 4120 17728 4126 17740
rect 5068 17731 5126 17737
rect 5068 17728 5080 17731
rect 4120 17700 5080 17728
rect 4120 17688 4126 17700
rect 5068 17697 5080 17700
rect 5114 17728 5126 17731
rect 6822 17728 6828 17740
rect 5114 17700 6828 17728
rect 5114 17697 5126 17700
rect 5068 17691 5126 17697
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 7558 17688 7564 17740
rect 7616 17728 7622 17740
rect 7653 17731 7711 17737
rect 7653 17728 7665 17731
rect 7616 17700 7665 17728
rect 7616 17688 7622 17700
rect 7653 17697 7665 17700
rect 7699 17697 7711 17731
rect 9030 17728 9036 17740
rect 8991 17700 9036 17728
rect 7653 17691 7711 17697
rect 9030 17688 9036 17700
rect 9088 17688 9094 17740
rect 11692 17731 11750 17737
rect 11692 17697 11704 17731
rect 11738 17728 11750 17731
rect 12158 17728 12164 17740
rect 11738 17700 12164 17728
rect 11738 17697 11750 17700
rect 11692 17691 11750 17697
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 15105 17731 15163 17737
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 15746 17728 15752 17740
rect 15151 17700 15752 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 1486 17660 1492 17672
rect 1447 17632 1492 17660
rect 1486 17620 1492 17632
rect 1544 17620 1550 17672
rect 3988 17660 4016 17688
rect 16040 17672 16068 17768
rect 17212 17765 17224 17768
rect 17258 17796 17270 17799
rect 17862 17796 17868 17808
rect 17258 17768 17868 17796
rect 17258 17765 17270 17768
rect 17212 17759 17270 17765
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 23658 17756 23664 17808
rect 23716 17796 23722 17808
rect 23753 17799 23811 17805
rect 23753 17796 23765 17799
rect 23716 17768 23765 17796
rect 23716 17756 23722 17768
rect 23753 17765 23765 17768
rect 23799 17796 23811 17799
rect 24765 17799 24823 17805
rect 24765 17796 24777 17799
rect 23799 17768 24777 17796
rect 23799 17765 23811 17768
rect 23753 17759 23811 17765
rect 24765 17765 24777 17768
rect 24811 17765 24823 17799
rect 24765 17759 24823 17765
rect 16945 17731 17003 17737
rect 16945 17697 16957 17731
rect 16991 17728 17003 17731
rect 17034 17728 17040 17740
rect 16991 17700 17040 17728
rect 16991 17697 17003 17700
rect 16945 17691 17003 17697
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19484 17700 19717 17728
rect 19484 17688 19490 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 21168 17731 21226 17737
rect 21168 17697 21180 17731
rect 21214 17728 21226 17731
rect 21450 17728 21456 17740
rect 21214 17700 21456 17728
rect 21214 17697 21226 17700
rect 21168 17691 21226 17697
rect 21450 17688 21456 17700
rect 21508 17688 21514 17740
rect 24949 17731 25007 17737
rect 24949 17697 24961 17731
rect 24995 17728 25007 17731
rect 25866 17728 25872 17740
rect 24995 17700 25872 17728
rect 24995 17697 25007 17700
rect 24949 17691 25007 17697
rect 25866 17688 25872 17700
rect 25924 17688 25930 17740
rect 4801 17663 4859 17669
rect 4801 17660 4813 17663
rect 3988 17632 4813 17660
rect 4801 17629 4813 17632
rect 4847 17629 4859 17663
rect 7926 17660 7932 17672
rect 7887 17632 7932 17660
rect 4801 17623 4859 17629
rect 7926 17620 7932 17632
rect 7984 17620 7990 17672
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 9456 17632 10149 17660
rect 9456 17620 9462 17632
rect 10137 17629 10149 17632
rect 10183 17660 10195 17663
rect 10226 17660 10232 17672
rect 10183 17632 10232 17660
rect 10183 17629 10195 17632
rect 10137 17623 10195 17629
rect 10226 17620 10232 17632
rect 10284 17620 10290 17672
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 11330 17660 11336 17672
rect 10367 17632 11336 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 11425 17663 11483 17669
rect 11425 17629 11437 17663
rect 11471 17629 11483 17663
rect 11425 17623 11483 17629
rect 14185 17663 14243 17669
rect 14185 17629 14197 17663
rect 14231 17660 14243 17663
rect 14826 17660 14832 17672
rect 14231 17632 14832 17660
rect 14231 17629 14243 17632
rect 14185 17623 14243 17629
rect 6914 17552 6920 17604
rect 6972 17592 6978 17604
rect 7285 17595 7343 17601
rect 7285 17592 7297 17595
rect 6972 17564 7297 17592
rect 6972 17552 6978 17564
rect 7285 17561 7297 17564
rect 7331 17561 7343 17595
rect 9674 17592 9680 17604
rect 9635 17564 9680 17592
rect 7285 17555 7343 17561
rect 9674 17552 9680 17564
rect 9732 17552 9738 17604
rect 2130 17484 2136 17536
rect 2188 17524 2194 17536
rect 2590 17524 2596 17536
rect 2188 17496 2596 17524
rect 2188 17484 2194 17496
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 4430 17524 4436 17536
rect 4387 17496 4436 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 6178 17524 6184 17536
rect 6139 17496 6184 17524
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 7800 17496 8309 17524
rect 7800 17484 7806 17496
rect 8297 17493 8309 17496
rect 8343 17493 8355 17527
rect 8297 17487 8355 17493
rect 8478 17484 8484 17536
rect 8536 17524 8542 17536
rect 8665 17527 8723 17533
rect 8665 17524 8677 17527
rect 8536 17496 8677 17524
rect 8536 17484 8542 17496
rect 8665 17493 8677 17496
rect 8711 17524 8723 17527
rect 9582 17524 9588 17536
rect 8711 17496 9588 17524
rect 8711 17493 8723 17496
rect 8665 17487 8723 17493
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 11440 17524 11468 17623
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 15838 17660 15844 17672
rect 15799 17632 15844 17660
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16022 17660 16028 17672
rect 15935 17632 16028 17660
rect 16022 17620 16028 17632
rect 16080 17620 16086 17672
rect 20806 17660 20812 17672
rect 19536 17632 20812 17660
rect 15378 17592 15384 17604
rect 15339 17564 15384 17592
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 11790 17524 11796 17536
rect 11440 17496 11796 17524
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 16485 17527 16543 17533
rect 16485 17493 16497 17527
rect 16531 17524 16543 17527
rect 16574 17524 16580 17536
rect 16531 17496 16580 17524
rect 16531 17493 16543 17496
rect 16485 17487 16543 17493
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 16853 17527 16911 17533
rect 16853 17493 16865 17527
rect 16899 17524 16911 17527
rect 16942 17524 16948 17536
rect 16899 17496 16948 17524
rect 16899 17493 16911 17496
rect 16853 17487 16911 17493
rect 16942 17484 16948 17496
rect 17000 17524 17006 17536
rect 18325 17527 18383 17533
rect 18325 17524 18337 17527
rect 17000 17496 18337 17524
rect 17000 17484 17006 17496
rect 18325 17493 18337 17496
rect 18371 17493 18383 17527
rect 18325 17487 18383 17493
rect 18690 17484 18696 17536
rect 18748 17524 18754 17536
rect 19242 17524 19248 17536
rect 18748 17496 19248 17524
rect 18748 17484 18754 17496
rect 19242 17484 19248 17496
rect 19300 17524 19306 17536
rect 19536 17533 19564 17632
rect 20806 17620 20812 17632
rect 20864 17660 20870 17672
rect 20901 17663 20959 17669
rect 20901 17660 20913 17663
rect 20864 17632 20913 17660
rect 20864 17620 20870 17632
rect 20901 17629 20913 17632
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 22922 17620 22928 17672
rect 22980 17660 22986 17672
rect 23845 17663 23903 17669
rect 23845 17660 23857 17663
rect 22980 17632 23857 17660
rect 22980 17620 22986 17632
rect 23845 17629 23857 17632
rect 23891 17629 23903 17663
rect 24026 17660 24032 17672
rect 23987 17632 24032 17660
rect 23845 17623 23903 17629
rect 24026 17620 24032 17632
rect 24084 17620 24090 17672
rect 23293 17595 23351 17601
rect 23293 17561 23305 17595
rect 23339 17592 23351 17595
rect 24044 17592 24072 17620
rect 23339 17564 24072 17592
rect 23339 17561 23351 17564
rect 23293 17555 23351 17561
rect 19521 17527 19579 17533
rect 19521 17524 19533 17527
rect 19300 17496 19533 17524
rect 19300 17484 19306 17496
rect 19521 17493 19533 17496
rect 19567 17493 19579 17527
rect 19521 17487 19579 17493
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 23106 17524 23112 17536
rect 22244 17496 23112 17524
rect 22244 17484 22250 17496
rect 23106 17484 23112 17496
rect 23164 17484 23170 17536
rect 23382 17524 23388 17536
rect 23343 17496 23388 17524
rect 23382 17484 23388 17496
rect 23440 17484 23446 17536
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24397 17527 24455 17533
rect 24397 17524 24409 17527
rect 24268 17496 24409 17524
rect 24268 17484 24274 17496
rect 24397 17493 24409 17496
rect 24443 17493 24455 17527
rect 25130 17524 25136 17536
rect 25091 17496 25136 17524
rect 24397 17487 24455 17493
rect 25130 17484 25136 17496
rect 25188 17484 25194 17536
rect 25590 17524 25596 17536
rect 25551 17496 25596 17524
rect 25590 17484 25596 17496
rect 25648 17484 25654 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17280 1584 17332
rect 1636 17320 1642 17332
rect 2774 17320 2780 17332
rect 1636 17292 2780 17320
rect 1636 17280 1642 17292
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3421 17323 3479 17329
rect 3421 17289 3433 17323
rect 3467 17320 3479 17323
rect 3786 17320 3792 17332
rect 3467 17292 3792 17320
rect 3467 17289 3479 17292
rect 3421 17283 3479 17289
rect 3786 17280 3792 17292
rect 3844 17280 3850 17332
rect 4062 17320 4068 17332
rect 4023 17292 4068 17320
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 4709 17323 4767 17329
rect 4709 17320 4721 17323
rect 4212 17292 4721 17320
rect 4212 17280 4218 17292
rect 4709 17289 4721 17292
rect 4755 17320 4767 17323
rect 4755 17292 5396 17320
rect 4755 17289 4767 17292
rect 4709 17283 4767 17289
rect 1486 17212 1492 17264
rect 1544 17252 1550 17264
rect 1857 17255 1915 17261
rect 1857 17252 1869 17255
rect 1544 17224 1869 17252
rect 1544 17212 1550 17224
rect 1857 17221 1869 17224
rect 1903 17252 1915 17255
rect 1946 17252 1952 17264
rect 1903 17224 1952 17252
rect 1903 17221 1915 17224
rect 1857 17215 1915 17221
rect 1946 17212 1952 17224
rect 2004 17252 2010 17264
rect 2004 17224 2084 17252
rect 2004 17212 2010 17224
rect 2056 17193 2084 17224
rect 3970 17212 3976 17264
rect 4028 17252 4034 17264
rect 4338 17252 4344 17264
rect 4028 17224 4344 17252
rect 4028 17212 4034 17224
rect 4338 17212 4344 17224
rect 4396 17212 4402 17264
rect 5368 17196 5396 17292
rect 5442 17280 5448 17332
rect 5500 17320 5506 17332
rect 7009 17323 7067 17329
rect 7009 17320 7021 17323
rect 5500 17292 7021 17320
rect 5500 17280 5506 17292
rect 7009 17289 7021 17292
rect 7055 17289 7067 17323
rect 7834 17320 7840 17332
rect 7795 17292 7840 17320
rect 7009 17283 7067 17289
rect 7834 17280 7840 17292
rect 7892 17280 7898 17332
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 9950 17320 9956 17332
rect 9732 17292 9956 17320
rect 9732 17280 9738 17292
rect 9950 17280 9956 17292
rect 10008 17280 10014 17332
rect 10045 17323 10103 17329
rect 10045 17289 10057 17323
rect 10091 17320 10103 17323
rect 10226 17320 10232 17332
rect 10091 17292 10232 17320
rect 10091 17289 10103 17292
rect 10045 17283 10103 17289
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 11790 17320 11796 17332
rect 11751 17292 11796 17320
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 12158 17320 12164 17332
rect 12119 17292 12164 17320
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12621 17323 12679 17329
rect 12621 17289 12633 17323
rect 12667 17320 12679 17323
rect 13262 17320 13268 17332
rect 12667 17292 13268 17320
rect 12667 17289 12679 17292
rect 12621 17283 12679 17289
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 13630 17320 13636 17332
rect 13591 17292 13636 17320
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 15749 17323 15807 17329
rect 15749 17289 15761 17323
rect 15795 17320 15807 17323
rect 16022 17320 16028 17332
rect 15795 17292 16028 17320
rect 15795 17289 15807 17292
rect 15749 17283 15807 17289
rect 16022 17280 16028 17292
rect 16080 17280 16086 17332
rect 16393 17323 16451 17329
rect 16393 17289 16405 17323
rect 16439 17320 16451 17323
rect 16482 17320 16488 17332
rect 16439 17292 16488 17320
rect 16439 17289 16451 17292
rect 16393 17283 16451 17289
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 17034 17280 17040 17332
rect 17092 17320 17098 17332
rect 17405 17323 17463 17329
rect 17405 17320 17417 17323
rect 17092 17292 17417 17320
rect 17092 17280 17098 17292
rect 17405 17289 17417 17292
rect 17451 17320 17463 17323
rect 18509 17323 18567 17329
rect 18509 17320 18521 17323
rect 17451 17292 18521 17320
rect 17451 17289 17463 17292
rect 17405 17283 17463 17289
rect 18509 17289 18521 17292
rect 18555 17289 18567 17323
rect 18509 17283 18567 17289
rect 6270 17212 6276 17264
rect 6328 17252 6334 17264
rect 6641 17255 6699 17261
rect 6641 17252 6653 17255
rect 6328 17224 6653 17252
rect 6328 17212 6334 17224
rect 6641 17221 6653 17224
rect 6687 17252 6699 17255
rect 7926 17252 7932 17264
rect 6687 17224 7932 17252
rect 6687 17221 6699 17224
rect 6641 17215 6699 17221
rect 7926 17212 7932 17224
rect 7984 17212 7990 17264
rect 9398 17252 9404 17264
rect 9359 17224 9404 17252
rect 9398 17212 9404 17224
rect 9456 17212 9462 17264
rect 12710 17212 12716 17264
rect 12768 17252 12774 17264
rect 12897 17255 12955 17261
rect 12897 17252 12909 17255
rect 12768 17224 12909 17252
rect 12768 17212 12774 17224
rect 12897 17221 12909 17224
rect 12943 17221 12955 17255
rect 12897 17215 12955 17221
rect 2041 17187 2099 17193
rect 2041 17153 2053 17187
rect 2087 17153 2099 17187
rect 5350 17184 5356 17196
rect 5263 17156 5356 17184
rect 2041 17147 2099 17153
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5534 17184 5540 17196
rect 5495 17156 5540 17184
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 11422 17184 11428 17196
rect 11383 17156 11428 17184
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 13648 17184 13676 17280
rect 13725 17187 13783 17193
rect 13725 17184 13737 17187
rect 13648 17156 13737 17184
rect 13725 17153 13737 17156
rect 13771 17153 13783 17187
rect 16942 17184 16948 17196
rect 16903 17156 16948 17184
rect 13725 17147 13783 17153
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 18524 17184 18552 17283
rect 22370 17280 22376 17332
rect 22428 17320 22434 17332
rect 23198 17320 23204 17332
rect 22428 17292 23204 17320
rect 22428 17280 22434 17292
rect 23198 17280 23204 17292
rect 23256 17280 23262 17332
rect 20806 17212 20812 17264
rect 20864 17252 20870 17264
rect 20901 17255 20959 17261
rect 20901 17252 20913 17255
rect 20864 17224 20913 17252
rect 20864 17212 20870 17224
rect 20901 17221 20913 17224
rect 20947 17252 20959 17255
rect 23106 17252 23112 17264
rect 20947 17224 23112 17252
rect 20947 17221 20959 17224
rect 20901 17215 20959 17221
rect 23106 17212 23112 17224
rect 23164 17252 23170 17264
rect 23385 17255 23443 17261
rect 23385 17252 23397 17255
rect 23164 17224 23397 17252
rect 23164 17212 23170 17224
rect 23385 17221 23397 17224
rect 23431 17252 23443 17255
rect 23431 17224 23704 17252
rect 23431 17221 23443 17224
rect 23385 17215 23443 17221
rect 18690 17184 18696 17196
rect 18524 17156 18696 17184
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 21821 17187 21879 17193
rect 21821 17153 21833 17187
rect 21867 17184 21879 17187
rect 22462 17184 22468 17196
rect 21867 17156 22468 17184
rect 21867 17153 21879 17156
rect 21821 17147 21879 17153
rect 22462 17144 22468 17156
rect 22520 17144 22526 17196
rect 23676 17193 23704 17224
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17153 23719 17187
rect 23661 17147 23719 17153
rect 2314 17125 2320 17128
rect 2308 17116 2320 17125
rect 2275 17088 2320 17116
rect 2308 17079 2320 17088
rect 2314 17076 2320 17079
rect 2372 17076 2378 17128
rect 4982 17076 4988 17128
rect 5040 17116 5046 17128
rect 5261 17119 5319 17125
rect 5261 17116 5273 17119
rect 5040 17088 5273 17116
rect 5040 17076 5046 17088
rect 5261 17085 5273 17088
rect 5307 17085 5319 17119
rect 5261 17079 5319 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 6871 17088 7512 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 2590 16980 2596 16992
rect 1820 16952 2596 16980
rect 1820 16940 1826 16952
rect 2590 16940 2596 16952
rect 2648 16940 2654 16992
rect 4890 16980 4896 16992
rect 4851 16952 4896 16980
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 5994 16980 6000 16992
rect 5955 16952 6000 16980
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 7484 16989 7512 17088
rect 7742 17076 7748 17128
rect 7800 17116 7806 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7800 17088 8033 17116
rect 7800 17076 7806 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 11149 17119 11207 17125
rect 11149 17116 11161 17119
rect 10836 17088 11161 17116
rect 10836 17076 10842 17088
rect 11149 17085 11161 17088
rect 11195 17085 11207 17119
rect 11149 17079 11207 17085
rect 11241 17119 11299 17125
rect 11241 17085 11253 17119
rect 11287 17116 11299 17119
rect 11330 17116 11336 17128
rect 11287 17088 11336 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 8288 17051 8346 17057
rect 8288 17017 8300 17051
rect 8334 17048 8346 17051
rect 8478 17048 8484 17060
rect 8334 17020 8484 17048
rect 8334 17017 8346 17020
rect 8288 17011 8346 17017
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 10042 17008 10048 17060
rect 10100 17048 10106 17060
rect 10689 17051 10747 17057
rect 10689 17048 10701 17051
rect 10100 17020 10701 17048
rect 10100 17008 10106 17020
rect 10689 17017 10701 17020
rect 10735 17048 10747 17051
rect 11256 17048 11284 17079
rect 11330 17076 11336 17088
rect 11388 17076 11394 17128
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12492 17088 12537 17116
rect 12492 17076 12498 17088
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 13992 17119 14050 17125
rect 13992 17116 14004 17119
rect 13872 17088 14004 17116
rect 13872 17076 13878 17088
rect 13992 17085 14004 17088
rect 14038 17116 14050 17119
rect 15102 17116 15108 17128
rect 14038 17088 15108 17116
rect 14038 17085 14050 17088
rect 13992 17079 14050 17085
rect 15102 17076 15108 17088
rect 15160 17076 15166 17128
rect 16301 17119 16359 17125
rect 16301 17085 16313 17119
rect 16347 17116 16359 17119
rect 16758 17116 16764 17128
rect 16347 17088 16764 17116
rect 16347 17085 16359 17088
rect 16301 17079 16359 17085
rect 16758 17076 16764 17088
rect 16816 17076 16822 17128
rect 22094 17076 22100 17128
rect 22152 17116 22158 17128
rect 22281 17119 22339 17125
rect 22281 17116 22293 17119
rect 22152 17088 22293 17116
rect 22152 17076 22158 17088
rect 22281 17085 22293 17088
rect 22327 17085 22339 17119
rect 22281 17079 22339 17085
rect 10735 17020 11284 17048
rect 10735 17017 10747 17020
rect 10689 17011 10747 17017
rect 16574 17008 16580 17060
rect 16632 17048 16638 17060
rect 16853 17051 16911 17057
rect 16853 17048 16865 17051
rect 16632 17020 16865 17048
rect 16632 17008 16638 17020
rect 16853 17017 16865 17020
rect 16899 17017 16911 17051
rect 18938 17051 18996 17057
rect 18938 17048 18950 17051
rect 16853 17011 16911 17017
rect 18708 17020 18950 17048
rect 18708 16992 18736 17020
rect 18938 17017 18950 17020
rect 18984 17017 18996 17051
rect 18938 17011 18996 17017
rect 21634 17008 21640 17060
rect 21692 17048 21698 17060
rect 22373 17051 22431 17057
rect 22373 17048 22385 17051
rect 21692 17020 22385 17048
rect 21692 17008 21698 17020
rect 22373 17017 22385 17020
rect 22419 17017 22431 17051
rect 22373 17011 22431 17017
rect 23109 17051 23167 17057
rect 23109 17017 23121 17051
rect 23155 17048 23167 17051
rect 23928 17051 23986 17057
rect 23928 17048 23940 17051
rect 23155 17020 23940 17048
rect 23155 17017 23167 17020
rect 23109 17011 23167 17017
rect 23928 17017 23940 17020
rect 23974 17048 23986 17051
rect 24026 17048 24032 17060
rect 23974 17020 24032 17048
rect 23974 17017 23986 17020
rect 23928 17011 23986 17017
rect 24026 17008 24032 17020
rect 24084 17008 24090 17060
rect 7469 16983 7527 16989
rect 7469 16949 7481 16983
rect 7515 16980 7527 16983
rect 7834 16980 7840 16992
rect 7515 16952 7840 16980
rect 7515 16949 7527 16952
rect 7469 16943 7527 16949
rect 7834 16940 7840 16952
rect 7892 16940 7898 16992
rect 10778 16980 10784 16992
rect 10739 16952 10784 16980
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 14550 16940 14556 16992
rect 14608 16980 14614 16992
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 14608 16952 15117 16980
rect 14608 16940 14614 16952
rect 15105 16949 15117 16952
rect 15151 16949 15163 16983
rect 17862 16980 17868 16992
rect 17823 16952 17868 16980
rect 15105 16943 15163 16949
rect 17862 16940 17868 16952
rect 17920 16940 17926 16992
rect 18690 16940 18696 16992
rect 18748 16940 18754 16992
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 20073 16983 20131 16989
rect 20073 16980 20085 16983
rect 19576 16952 20085 16980
rect 19576 16940 19582 16952
rect 20073 16949 20085 16952
rect 20119 16949 20131 16983
rect 20073 16943 20131 16949
rect 21361 16983 21419 16989
rect 21361 16949 21373 16983
rect 21407 16980 21419 16983
rect 21450 16980 21456 16992
rect 21407 16952 21456 16980
rect 21407 16949 21419 16952
rect 21361 16943 21419 16949
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 21913 16983 21971 16989
rect 21913 16949 21925 16983
rect 21959 16980 21971 16983
rect 22922 16980 22928 16992
rect 21959 16952 22928 16980
rect 21959 16949 21971 16952
rect 21913 16943 21971 16949
rect 22922 16940 22928 16952
rect 22980 16940 22986 16992
rect 25038 16980 25044 16992
rect 24999 16952 25044 16980
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 25685 16983 25743 16989
rect 25685 16949 25697 16983
rect 25731 16980 25743 16983
rect 25866 16980 25872 16992
rect 25731 16952 25872 16980
rect 25731 16949 25743 16952
rect 25685 16943 25743 16949
rect 25866 16940 25872 16952
rect 25924 16940 25930 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1946 16776 1952 16788
rect 1728 16748 1952 16776
rect 1728 16736 1734 16748
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 2222 16776 2228 16788
rect 2183 16748 2228 16776
rect 2222 16736 2228 16748
rect 2280 16736 2286 16788
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 2866 16776 2872 16788
rect 2455 16748 2872 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 2866 16736 2872 16748
rect 2924 16736 2930 16788
rect 3142 16736 3148 16788
rect 3200 16776 3206 16788
rect 4246 16776 4252 16788
rect 3200 16748 4108 16776
rect 4207 16748 4252 16776
rect 3200 16736 3206 16748
rect 2498 16708 2504 16720
rect 1412 16680 2504 16708
rect 1412 16649 1440 16680
rect 1964 16652 1992 16680
rect 2498 16668 2504 16680
rect 2556 16668 2562 16720
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16708 2835 16711
rect 2823 16680 3924 16708
rect 2823 16677 2835 16680
rect 2777 16671 2835 16677
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16609 1455 16643
rect 1397 16603 1455 16609
rect 1946 16600 1952 16652
rect 2004 16600 2010 16652
rect 2314 16600 2320 16652
rect 2372 16640 2378 16652
rect 3896 16649 3924 16680
rect 4080 16652 4108 16748
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 4982 16776 4988 16788
rect 4943 16748 4988 16776
rect 4982 16736 4988 16748
rect 5040 16736 5046 16788
rect 5166 16736 5172 16788
rect 5224 16776 5230 16788
rect 6822 16776 6828 16788
rect 5224 16748 5856 16776
rect 6783 16748 6828 16776
rect 5224 16736 5230 16748
rect 5353 16711 5411 16717
rect 5353 16677 5365 16711
rect 5399 16708 5411 16711
rect 5534 16708 5540 16720
rect 5399 16680 5540 16708
rect 5399 16677 5411 16680
rect 5353 16671 5411 16677
rect 5534 16668 5540 16680
rect 5592 16708 5598 16720
rect 5690 16711 5748 16717
rect 5690 16708 5702 16711
rect 5592 16680 5702 16708
rect 5592 16668 5598 16680
rect 5690 16677 5702 16680
rect 5736 16677 5748 16711
rect 5828 16708 5856 16748
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 7469 16779 7527 16785
rect 7469 16745 7481 16779
rect 7515 16776 7527 16779
rect 7558 16776 7564 16788
rect 7515 16748 7564 16776
rect 7515 16745 7527 16748
rect 7469 16739 7527 16745
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 8202 16736 8208 16788
rect 8260 16736 8266 16788
rect 8386 16776 8392 16788
rect 8347 16748 8392 16776
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 9125 16779 9183 16785
rect 9125 16745 9137 16779
rect 9171 16776 9183 16779
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 9171 16748 10977 16776
rect 9171 16745 9183 16748
rect 9125 16739 9183 16745
rect 10965 16745 10977 16748
rect 11011 16776 11023 16779
rect 11422 16776 11428 16788
rect 11011 16748 11428 16776
rect 11011 16745 11023 16748
rect 10965 16739 11023 16745
rect 11422 16736 11428 16748
rect 11480 16736 11486 16788
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13357 16779 13415 16785
rect 13357 16776 13369 16779
rect 12952 16748 13369 16776
rect 12952 16736 12958 16748
rect 13357 16745 13369 16748
rect 13403 16745 13415 16779
rect 13814 16776 13820 16788
rect 13775 16748 13820 16776
rect 13357 16739 13415 16745
rect 13814 16736 13820 16748
rect 13872 16736 13878 16788
rect 15286 16776 15292 16788
rect 15247 16748 15292 16776
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15933 16779 15991 16785
rect 15933 16745 15945 16779
rect 15979 16776 15991 16779
rect 16942 16776 16948 16788
rect 15979 16748 16948 16776
rect 15979 16745 15991 16748
rect 15933 16739 15991 16745
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 17773 16779 17831 16785
rect 17773 16745 17785 16779
rect 17819 16776 17831 16779
rect 17862 16776 17868 16788
rect 17819 16748 17868 16776
rect 17819 16745 17831 16748
rect 17773 16739 17831 16745
rect 17862 16736 17868 16748
rect 17920 16736 17926 16788
rect 18690 16776 18696 16788
rect 18651 16748 18696 16776
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 18874 16776 18880 16788
rect 18835 16748 18880 16776
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 19242 16776 19248 16788
rect 19203 16748 19248 16776
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 20714 16776 20720 16788
rect 19392 16748 19437 16776
rect 20675 16748 20720 16776
rect 19392 16736 19398 16748
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 20806 16736 20812 16788
rect 20864 16776 20870 16788
rect 20901 16779 20959 16785
rect 20901 16776 20913 16779
rect 20864 16748 20913 16776
rect 20864 16736 20870 16748
rect 20901 16745 20913 16748
rect 20947 16745 20959 16779
rect 20901 16739 20959 16745
rect 21634 16736 21640 16788
rect 21692 16776 21698 16788
rect 21913 16779 21971 16785
rect 21913 16776 21925 16779
rect 21692 16748 21925 16776
rect 21692 16736 21698 16748
rect 21913 16745 21925 16748
rect 21959 16745 21971 16779
rect 21913 16739 21971 16745
rect 22094 16736 22100 16788
rect 22152 16776 22158 16788
rect 22281 16779 22339 16785
rect 22281 16776 22293 16779
rect 22152 16748 22293 16776
rect 22152 16736 22158 16748
rect 22281 16745 22293 16748
rect 22327 16745 22339 16779
rect 22922 16776 22928 16788
rect 22883 16748 22928 16776
rect 22281 16739 22339 16745
rect 22922 16736 22928 16748
rect 22980 16736 22986 16788
rect 24394 16776 24400 16788
rect 24355 16748 24400 16776
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 7745 16711 7803 16717
rect 7745 16708 7757 16711
rect 5828 16680 7757 16708
rect 5690 16671 5748 16677
rect 7745 16677 7757 16680
rect 7791 16677 7803 16711
rect 7745 16671 7803 16677
rect 3421 16643 3479 16649
rect 3421 16640 3433 16643
rect 2372 16612 3433 16640
rect 2372 16600 2378 16612
rect 3421 16609 3433 16612
rect 3467 16609 3479 16643
rect 3421 16603 3479 16609
rect 3881 16643 3939 16649
rect 3881 16609 3893 16643
rect 3927 16640 3939 16643
rect 3927 16612 4016 16640
rect 3927 16609 3939 16612
rect 3881 16603 3939 16609
rect 2869 16575 2927 16581
rect 2869 16541 2881 16575
rect 2915 16541 2927 16575
rect 3050 16572 3056 16584
rect 2963 16544 3056 16572
rect 2869 16535 2927 16541
rect 1762 16464 1768 16516
rect 1820 16504 1826 16516
rect 2590 16504 2596 16516
rect 1820 16476 2596 16504
rect 1820 16464 1826 16476
rect 2590 16464 2596 16476
rect 2648 16464 2654 16516
rect 2884 16504 2912 16535
rect 3050 16532 3056 16544
rect 3108 16572 3114 16584
rect 3988 16572 4016 16612
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4120 16612 4213 16640
rect 4120 16600 4126 16612
rect 4338 16600 4344 16652
rect 4396 16640 4402 16652
rect 5442 16640 5448 16652
rect 4396 16612 5448 16640
rect 4396 16600 4402 16612
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 7558 16600 7564 16652
rect 7616 16640 7622 16652
rect 8220 16640 8248 16736
rect 9306 16668 9312 16720
rect 9364 16708 9370 16720
rect 23290 16717 23296 16720
rect 9401 16711 9459 16717
rect 9401 16708 9413 16711
rect 9364 16680 9413 16708
rect 9364 16668 9370 16680
rect 9401 16677 9413 16680
rect 9447 16677 9459 16711
rect 23284 16708 23296 16717
rect 9401 16671 9459 16677
rect 9600 16680 10272 16708
rect 23251 16680 23296 16708
rect 7616 16612 8248 16640
rect 8481 16643 8539 16649
rect 7616 16600 7622 16612
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 9030 16640 9036 16652
rect 8527 16612 9036 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 5166 16572 5172 16584
rect 3108 16544 3924 16572
rect 3988 16544 5172 16572
rect 3108 16532 3114 16544
rect 3694 16504 3700 16516
rect 2884 16476 3700 16504
rect 3694 16464 3700 16476
rect 3752 16464 3758 16516
rect 3896 16504 3924 16544
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 8665 16575 8723 16581
rect 8665 16541 8677 16575
rect 8711 16572 8723 16575
rect 8846 16572 8852 16584
rect 8711 16544 8852 16572
rect 8711 16541 8723 16544
rect 8665 16535 8723 16541
rect 8846 16532 8852 16544
rect 8904 16532 8910 16584
rect 9490 16532 9496 16584
rect 9548 16572 9554 16584
rect 9600 16572 9628 16680
rect 10244 16649 10272 16680
rect 23284 16671 23296 16680
rect 23290 16668 23296 16671
rect 23348 16668 23354 16720
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16640 10287 16643
rect 10962 16640 10968 16652
rect 10275 16612 10968 16640
rect 10275 16609 10287 16612
rect 10229 16603 10287 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11330 16600 11336 16652
rect 11388 16640 11394 16652
rect 11681 16643 11739 16649
rect 11681 16640 11693 16643
rect 11388 16612 11693 16640
rect 11388 16600 11394 16612
rect 11681 16609 11693 16612
rect 11727 16609 11739 16643
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 11681 16603 11739 16609
rect 13832 16612 13921 16640
rect 9548 16544 9628 16572
rect 9548 16532 9554 16544
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10321 16575 10379 16581
rect 10321 16572 10333 16575
rect 10192 16544 10333 16572
rect 10192 16532 10198 16544
rect 10321 16541 10333 16544
rect 10367 16541 10379 16575
rect 10321 16535 10379 16541
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16572 10563 16575
rect 10870 16572 10876 16584
rect 10551 16544 10876 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 11425 16575 11483 16581
rect 11425 16541 11437 16575
rect 11471 16541 11483 16575
rect 11425 16535 11483 16541
rect 3970 16504 3976 16516
rect 3896 16476 3976 16504
rect 3970 16464 3976 16476
rect 4028 16504 4034 16516
rect 4246 16504 4252 16516
rect 4028 16476 4252 16504
rect 4028 16464 4034 16476
rect 4246 16464 4252 16476
rect 4304 16464 4310 16516
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 9861 16507 9919 16513
rect 9861 16504 9873 16507
rect 9640 16476 9873 16504
rect 9640 16464 9646 16476
rect 9861 16473 9873 16476
rect 9907 16473 9919 16507
rect 9861 16467 9919 16473
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 11440 16504 11468 16535
rect 12986 16532 12992 16584
rect 13044 16572 13050 16584
rect 13832 16572 13860 16612
rect 13909 16609 13921 16612
rect 13955 16609 13967 16643
rect 14366 16640 14372 16652
rect 14327 16612 14372 16640
rect 13909 16603 13967 16609
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 15102 16640 15108 16652
rect 15063 16612 15108 16640
rect 15102 16600 15108 16612
rect 15160 16600 15166 16652
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16640 16359 16643
rect 16660 16643 16718 16649
rect 16660 16640 16672 16643
rect 16347 16612 16672 16640
rect 16347 16609 16359 16612
rect 16301 16603 16359 16609
rect 16660 16609 16672 16612
rect 16706 16640 16718 16643
rect 17034 16640 17040 16652
rect 16706 16612 17040 16640
rect 16706 16609 16718 16612
rect 16660 16603 16718 16609
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19889 16643 19947 16649
rect 19889 16640 19901 16643
rect 19484 16612 19901 16640
rect 19484 16600 19490 16612
rect 19889 16609 19901 16612
rect 19935 16609 19947 16643
rect 19889 16603 19947 16609
rect 20162 16600 20168 16652
rect 20220 16640 20226 16652
rect 20438 16640 20444 16652
rect 20220 16612 20444 16640
rect 20220 16600 20226 16612
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 20714 16640 20720 16652
rect 20627 16612 20720 16640
rect 13044 16544 13860 16572
rect 13044 16532 13050 16544
rect 16206 16532 16212 16584
rect 16264 16572 16270 16584
rect 16393 16575 16451 16581
rect 16393 16572 16405 16575
rect 16264 16544 16405 16572
rect 16264 16532 16270 16544
rect 16393 16541 16405 16544
rect 16439 16541 16451 16575
rect 19518 16572 19524 16584
rect 19479 16544 19524 16572
rect 16393 16535 16451 16541
rect 19518 16532 19524 16544
rect 19576 16532 19582 16584
rect 19978 16532 19984 16584
rect 20036 16572 20042 16584
rect 20640 16572 20668 16612
rect 20714 16600 20720 16612
rect 20772 16640 20778 16652
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 20772 16612 21281 16640
rect 20772 16600 20778 16612
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 23017 16643 23075 16649
rect 23017 16609 23029 16643
rect 23063 16640 23075 16643
rect 23106 16640 23112 16652
rect 23063 16612 23112 16640
rect 23063 16609 23075 16612
rect 23017 16603 23075 16609
rect 23106 16600 23112 16612
rect 23164 16600 23170 16652
rect 21358 16572 21364 16584
rect 20036 16544 20668 16572
rect 21319 16544 21364 16572
rect 20036 16532 20042 16544
rect 21358 16532 21364 16544
rect 21416 16532 21422 16584
rect 21545 16575 21603 16581
rect 21545 16541 21557 16575
rect 21591 16572 21603 16575
rect 21910 16572 21916 16584
rect 21591 16544 21916 16572
rect 21591 16541 21603 16544
rect 21545 16535 21603 16541
rect 21910 16532 21916 16544
rect 21968 16532 21974 16584
rect 11020 16476 11468 16504
rect 11020 16464 11026 16476
rect 2222 16396 2228 16448
rect 2280 16436 2286 16448
rect 2498 16436 2504 16448
rect 2280 16408 2504 16436
rect 2280 16396 2286 16408
rect 2498 16396 2504 16408
rect 2556 16396 2562 16448
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 11241 16439 11299 16445
rect 11241 16436 11253 16439
rect 11112 16408 11253 16436
rect 11112 16396 11118 16408
rect 11241 16405 11253 16408
rect 11287 16405 11299 16439
rect 11241 16399 11299 16405
rect 11698 16396 11704 16448
rect 11756 16436 11762 16448
rect 12805 16439 12863 16445
rect 12805 16436 12817 16439
rect 11756 16408 12817 16436
rect 11756 16396 11762 16408
rect 12805 16405 12817 16408
rect 12851 16405 12863 16439
rect 18414 16436 18420 16448
rect 18375 16408 18420 16436
rect 12805 16399 12863 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 20349 16439 20407 16445
rect 20349 16405 20361 16439
rect 20395 16436 20407 16439
rect 20438 16436 20444 16448
rect 20395 16408 20444 16436
rect 20395 16405 20407 16408
rect 20349 16399 20407 16405
rect 20438 16396 20444 16408
rect 20496 16396 20502 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1670 16192 1676 16244
rect 1728 16232 1734 16244
rect 2409 16235 2467 16241
rect 2409 16232 2421 16235
rect 1728 16204 2421 16232
rect 1728 16192 1734 16204
rect 2409 16201 2421 16204
rect 2455 16201 2467 16235
rect 5166 16232 5172 16244
rect 5127 16204 5172 16232
rect 2409 16195 2467 16201
rect 2424 16096 2452 16195
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 5442 16192 5448 16244
rect 5500 16232 5506 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5500 16204 6193 16232
rect 5500 16192 5506 16204
rect 5920 16176 5948 16204
rect 6181 16201 6193 16204
rect 6227 16232 6239 16235
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6227 16204 6561 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6549 16201 6561 16204
rect 6595 16232 6607 16235
rect 7742 16232 7748 16244
rect 6595 16204 7748 16232
rect 6595 16201 6607 16204
rect 6549 16195 6607 16201
rect 5074 16164 5080 16176
rect 5035 16136 5080 16164
rect 5074 16124 5080 16136
rect 5132 16124 5138 16176
rect 5902 16124 5908 16176
rect 5960 16124 5966 16176
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 2424 16068 2605 16096
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 4706 16096 4712 16108
rect 4619 16068 4712 16096
rect 2593 16059 2651 16065
rect 4706 16056 4712 16068
rect 4764 16096 4770 16108
rect 5534 16096 5540 16108
rect 4764 16068 5540 16096
rect 4764 16056 4770 16068
rect 5534 16056 5540 16068
rect 5592 16096 5598 16108
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5592 16068 5733 16096
rect 5592 16056 5598 16068
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 6564 16096 6592 16195
rect 7742 16192 7748 16204
rect 7800 16232 7806 16244
rect 9306 16232 9312 16244
rect 7800 16204 9312 16232
rect 7800 16192 7806 16204
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16232 9827 16235
rect 10134 16232 10140 16244
rect 9815 16204 10140 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 10962 16192 10968 16244
rect 11020 16232 11026 16244
rect 11790 16232 11796 16244
rect 11020 16204 11796 16232
rect 11020 16192 11026 16204
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 13998 16232 14004 16244
rect 13959 16204 14004 16232
rect 13998 16192 14004 16204
rect 14056 16192 14062 16244
rect 14826 16192 14832 16244
rect 14884 16232 14890 16244
rect 15473 16235 15531 16241
rect 15473 16232 15485 16235
rect 14884 16204 15485 16232
rect 14884 16192 14890 16204
rect 15473 16201 15485 16204
rect 15519 16201 15531 16235
rect 15473 16195 15531 16201
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 12802 16164 12808 16176
rect 11112 16136 12808 16164
rect 11112 16124 11118 16136
rect 12802 16124 12808 16136
rect 12860 16164 12866 16176
rect 12860 16136 13032 16164
rect 12860 16124 12866 16136
rect 13004 16105 13032 16136
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6564 16068 6837 16096
rect 5721 16059 5779 16065
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16096 13047 16099
rect 13449 16099 13507 16105
rect 13449 16096 13461 16099
rect 13035 16068 13461 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 13449 16065 13461 16068
rect 13495 16065 13507 16099
rect 14550 16096 14556 16108
rect 13449 16059 13507 16065
rect 13832 16068 14556 16096
rect 13832 16040 13860 16068
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1443 16000 2084 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1578 15892 1584 15904
rect 1539 15864 1584 15892
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 2056 15901 2084 16000
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 5629 16031 5687 16037
rect 5629 16028 5641 16031
rect 4396 16000 5641 16028
rect 4396 15988 4402 16000
rect 5629 15997 5641 16000
rect 5675 16028 5687 16031
rect 5994 16028 6000 16040
rect 5675 16000 6000 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 5994 15988 6000 16000
rect 6052 15988 6058 16040
rect 9306 15988 9312 16040
rect 9364 16028 9370 16040
rect 9861 16031 9919 16037
rect 9861 16028 9873 16031
rect 9364 16000 9873 16028
rect 9364 15988 9370 16000
rect 9861 15997 9873 16000
rect 9907 15997 9919 16031
rect 13814 16028 13820 16040
rect 13775 16000 13820 16028
rect 9861 15991 9919 15997
rect 13814 15988 13820 16000
rect 13872 15988 13878 16040
rect 14366 16028 14372 16040
rect 14327 16000 14372 16028
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 15488 16028 15516 16195
rect 15746 16192 15752 16244
rect 15804 16232 15810 16244
rect 16393 16235 16451 16241
rect 16393 16232 16405 16235
rect 15804 16204 16405 16232
rect 15804 16192 15810 16204
rect 16393 16201 16405 16204
rect 16439 16201 16451 16235
rect 18046 16232 18052 16244
rect 18007 16204 18052 16232
rect 16393 16195 16451 16201
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 19334 16192 19340 16244
rect 19392 16232 19398 16244
rect 19429 16235 19487 16241
rect 19429 16232 19441 16235
rect 19392 16204 19441 16232
rect 19392 16192 19398 16204
rect 19429 16201 19441 16204
rect 19475 16201 19487 16235
rect 19978 16232 19984 16244
rect 19939 16204 19984 16232
rect 19429 16195 19487 16201
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 21358 16192 21364 16244
rect 21416 16232 21422 16244
rect 21545 16235 21603 16241
rect 21545 16232 21557 16235
rect 21416 16204 21557 16232
rect 21416 16192 21422 16204
rect 21545 16201 21557 16204
rect 21591 16232 21603 16235
rect 22002 16232 22008 16244
rect 21591 16204 22008 16232
rect 21591 16201 21603 16204
rect 21545 16195 21603 16201
rect 22002 16192 22008 16204
rect 22060 16192 22066 16244
rect 23106 16232 23112 16244
rect 23067 16204 23112 16232
rect 23106 16192 23112 16204
rect 23164 16232 23170 16244
rect 23385 16235 23443 16241
rect 23385 16232 23397 16235
rect 23164 16204 23397 16232
rect 23164 16192 23170 16204
rect 23385 16201 23397 16204
rect 23431 16201 23443 16235
rect 23385 16195 23443 16201
rect 21085 16167 21143 16173
rect 21085 16133 21097 16167
rect 21131 16164 21143 16167
rect 21910 16164 21916 16176
rect 21131 16136 21916 16164
rect 21131 16133 21143 16136
rect 21085 16127 21143 16133
rect 21910 16124 21916 16136
rect 21968 16124 21974 16176
rect 22741 16167 22799 16173
rect 22741 16133 22753 16167
rect 22787 16164 22799 16167
rect 23290 16164 23296 16176
rect 22787 16136 23296 16164
rect 22787 16133 22799 16136
rect 22741 16127 22799 16133
rect 23290 16124 23296 16136
rect 23348 16124 23354 16176
rect 17034 16096 17040 16108
rect 16947 16068 17040 16096
rect 17034 16056 17040 16068
rect 17092 16096 17098 16108
rect 18414 16096 18420 16108
rect 17092 16068 18420 16096
rect 17092 16056 17098 16068
rect 18414 16056 18420 16068
rect 18472 16096 18478 16108
rect 18601 16099 18659 16105
rect 18601 16096 18613 16099
rect 18472 16068 18613 16096
rect 18472 16056 18478 16068
rect 18601 16065 18613 16068
rect 18647 16065 18659 16099
rect 18601 16059 18659 16065
rect 19889 16099 19947 16105
rect 19889 16065 19901 16099
rect 19935 16096 19947 16099
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 19935 16068 20545 16096
rect 19935 16065 19947 16068
rect 19889 16059 19947 16065
rect 20533 16065 20545 16068
rect 20579 16096 20591 16099
rect 21361 16099 21419 16105
rect 21361 16096 21373 16099
rect 20579 16068 21373 16096
rect 20579 16065 20591 16068
rect 20533 16059 20591 16065
rect 21361 16065 21373 16068
rect 21407 16096 21419 16099
rect 21450 16096 21456 16108
rect 21407 16068 21456 16096
rect 21407 16065 21419 16068
rect 21361 16059 21419 16065
rect 21450 16056 21456 16068
rect 21508 16096 21514 16108
rect 22097 16099 22155 16105
rect 22097 16096 22109 16099
rect 21508 16068 22109 16096
rect 21508 16056 21514 16068
rect 22097 16065 22109 16068
rect 22143 16065 22155 16099
rect 23400 16096 23428 16195
rect 23661 16099 23719 16105
rect 23661 16096 23673 16099
rect 23400 16068 23673 16096
rect 22097 16059 22155 16065
rect 23661 16065 23673 16068
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 16761 16031 16819 16037
rect 16761 16028 16773 16031
rect 15488 16000 16773 16028
rect 16761 15997 16773 16000
rect 16807 15997 16819 16031
rect 16761 15991 16819 15997
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 16028 17555 16031
rect 18690 16028 18696 16040
rect 17543 16000 18696 16028
rect 17543 15997 17555 16000
rect 17497 15991 17555 15997
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 20349 16031 20407 16037
rect 20349 15997 20361 16031
rect 20395 16028 20407 16031
rect 20622 16028 20628 16040
rect 20395 16000 20628 16028
rect 20395 15997 20407 16000
rect 20349 15991 20407 15997
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 21726 15988 21732 16040
rect 21784 16028 21790 16040
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21784 16000 21925 16028
rect 21784 15988 21790 16000
rect 21913 15997 21925 16000
rect 21959 15997 21971 16031
rect 21913 15991 21971 15997
rect 2860 15963 2918 15969
rect 2860 15929 2872 15963
rect 2906 15960 2918 15963
rect 3326 15960 3332 15972
rect 2906 15932 3332 15960
rect 2906 15929 2918 15932
rect 2860 15923 2918 15929
rect 3326 15920 3332 15932
rect 3384 15920 3390 15972
rect 3804 15932 5028 15960
rect 2041 15895 2099 15901
rect 2041 15861 2053 15895
rect 2087 15892 2099 15895
rect 3804 15892 3832 15932
rect 3970 15892 3976 15904
rect 2087 15864 3832 15892
rect 3931 15864 3976 15892
rect 2087 15861 2099 15864
rect 2041 15855 2099 15861
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 5000 15892 5028 15932
rect 5074 15920 5080 15972
rect 5132 15960 5138 15972
rect 5537 15963 5595 15969
rect 5537 15960 5549 15963
rect 5132 15932 5549 15960
rect 5132 15920 5138 15932
rect 5537 15929 5549 15932
rect 5583 15929 5595 15963
rect 5537 15923 5595 15929
rect 7006 15920 7012 15972
rect 7064 15969 7070 15972
rect 7064 15963 7128 15969
rect 7064 15929 7082 15963
rect 7116 15929 7128 15963
rect 7064 15923 7128 15929
rect 10128 15963 10186 15969
rect 10128 15929 10140 15963
rect 10174 15960 10186 15963
rect 11054 15960 11060 15972
rect 10174 15932 11060 15960
rect 10174 15929 10186 15932
rect 10128 15923 10186 15929
rect 7064 15920 7070 15923
rect 11054 15920 11060 15932
rect 11112 15920 11118 15972
rect 12253 15963 12311 15969
rect 12253 15929 12265 15963
rect 12299 15960 12311 15963
rect 12805 15963 12863 15969
rect 12805 15960 12817 15963
rect 12299 15932 12817 15960
rect 12299 15929 12311 15932
rect 12253 15923 12311 15929
rect 12805 15929 12817 15932
rect 12851 15960 12863 15963
rect 12986 15960 12992 15972
rect 12851 15932 12992 15960
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 12986 15920 12992 15932
rect 13044 15920 13050 15972
rect 18874 15960 18880 15972
rect 18432 15932 18880 15960
rect 7190 15892 7196 15904
rect 5000 15864 7196 15892
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 7742 15852 7748 15904
rect 7800 15892 7806 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7800 15864 8217 15892
rect 7800 15852 7806 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 8849 15895 8907 15901
rect 8849 15861 8861 15895
rect 8895 15892 8907 15895
rect 9030 15892 9036 15904
rect 8895 15864 9036 15892
rect 8895 15861 8907 15864
rect 8849 15855 8907 15861
rect 9030 15852 9036 15864
rect 9088 15852 9094 15904
rect 11241 15895 11299 15901
rect 11241 15861 11253 15895
rect 11287 15892 11299 15895
rect 11514 15892 11520 15904
rect 11287 15864 11520 15892
rect 11287 15861 11299 15864
rect 11241 15855 11299 15861
rect 11514 15852 11520 15864
rect 11572 15852 11578 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 12897 15895 12955 15901
rect 12492 15864 12537 15892
rect 12492 15852 12498 15864
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13354 15892 13360 15904
rect 12943 15864 13360 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 14090 15852 14096 15904
rect 14148 15892 14154 15904
rect 14366 15892 14372 15904
rect 14148 15864 14372 15892
rect 14148 15852 14154 15864
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 14458 15852 14464 15904
rect 14516 15892 14522 15904
rect 15933 15895 15991 15901
rect 14516 15864 14561 15892
rect 14516 15852 14522 15864
rect 15933 15861 15945 15895
rect 15979 15892 15991 15895
rect 16206 15892 16212 15904
rect 15979 15864 16212 15892
rect 15979 15861 15991 15864
rect 15933 15855 15991 15861
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 16850 15892 16856 15904
rect 16347 15864 16856 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 17678 15852 17684 15904
rect 17736 15892 17742 15904
rect 18432 15901 18460 15932
rect 18874 15920 18880 15932
rect 18932 15920 18938 15972
rect 19153 15963 19211 15969
rect 19153 15929 19165 15963
rect 19199 15960 19211 15963
rect 19518 15960 19524 15972
rect 19199 15932 19524 15960
rect 19199 15929 19211 15932
rect 19153 15923 19211 15929
rect 19518 15920 19524 15932
rect 19576 15960 19582 15972
rect 20530 15960 20536 15972
rect 19576 15932 20536 15960
rect 19576 15920 19582 15932
rect 20530 15920 20536 15932
rect 20588 15920 20594 15972
rect 21266 15920 21272 15972
rect 21324 15960 21330 15972
rect 22005 15963 22063 15969
rect 22005 15960 22017 15963
rect 21324 15932 22017 15960
rect 21324 15920 21330 15932
rect 22005 15929 22017 15932
rect 22051 15929 22063 15963
rect 22005 15923 22063 15929
rect 23474 15920 23480 15972
rect 23532 15960 23538 15972
rect 23906 15963 23964 15969
rect 23906 15960 23918 15963
rect 23532 15932 23918 15960
rect 23532 15920 23538 15932
rect 23906 15929 23918 15932
rect 23952 15960 23964 15963
rect 24210 15960 24216 15972
rect 23952 15932 24216 15960
rect 23952 15929 23964 15932
rect 23906 15923 23964 15929
rect 24210 15920 24216 15932
rect 24268 15920 24274 15972
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 17736 15864 17785 15892
rect 17736 15852 17742 15864
rect 17773 15861 17785 15864
rect 17819 15892 17831 15895
rect 18417 15895 18475 15901
rect 18417 15892 18429 15895
rect 17819 15864 18429 15892
rect 17819 15861 17831 15864
rect 17773 15855 17831 15861
rect 18417 15861 18429 15864
rect 18463 15861 18475 15895
rect 18417 15855 18475 15861
rect 18509 15895 18567 15901
rect 18509 15861 18521 15895
rect 18555 15892 18567 15895
rect 18598 15892 18604 15904
rect 18555 15864 18604 15892
rect 18555 15861 18567 15864
rect 18509 15855 18567 15861
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 20438 15892 20444 15904
rect 20399 15864 20444 15892
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 24026 15852 24032 15904
rect 24084 15892 24090 15904
rect 25041 15895 25099 15901
rect 25041 15892 25053 15895
rect 24084 15864 25053 15892
rect 24084 15852 24090 15864
rect 25041 15861 25053 15864
rect 25087 15892 25099 15895
rect 25222 15892 25228 15904
rect 25087 15864 25228 15892
rect 25087 15861 25099 15864
rect 25041 15855 25099 15861
rect 25222 15852 25228 15864
rect 25280 15852 25286 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1854 15688 1860 15700
rect 1815 15660 1860 15688
rect 1854 15648 1860 15660
rect 1912 15648 1918 15700
rect 2038 15648 2044 15700
rect 2096 15648 2102 15700
rect 2961 15691 3019 15697
rect 2961 15657 2973 15691
rect 3007 15688 3019 15691
rect 3050 15688 3056 15700
rect 3007 15660 3056 15688
rect 3007 15657 3019 15660
rect 2961 15651 3019 15657
rect 3050 15648 3056 15660
rect 3108 15648 3114 15700
rect 3326 15688 3332 15700
rect 3287 15660 3332 15688
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 4338 15688 4344 15700
rect 4299 15660 4344 15688
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 4709 15691 4767 15697
rect 4709 15657 4721 15691
rect 4755 15688 4767 15691
rect 4798 15688 4804 15700
rect 4755 15660 4804 15688
rect 4755 15657 4767 15660
rect 4709 15651 4767 15657
rect 4798 15648 4804 15660
rect 4856 15648 4862 15700
rect 5534 15688 5540 15700
rect 5495 15660 5540 15688
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 8113 15691 8171 15697
rect 8113 15657 8125 15691
rect 8159 15688 8171 15691
rect 8202 15688 8208 15700
rect 8159 15660 8208 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 8757 15691 8815 15697
rect 8757 15688 8769 15691
rect 8720 15660 8769 15688
rect 8720 15648 8726 15660
rect 8757 15657 8769 15660
rect 8803 15657 8815 15691
rect 9490 15688 9496 15700
rect 9451 15660 9496 15688
rect 8757 15651 8815 15657
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9824 15660 9873 15688
rect 9824 15648 9830 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 9861 15651 9919 15657
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10229 15691 10287 15697
rect 10229 15688 10241 15691
rect 10008 15660 10241 15688
rect 10008 15648 10014 15660
rect 10229 15657 10241 15660
rect 10275 15657 10287 15691
rect 10870 15688 10876 15700
rect 10831 15660 10876 15688
rect 10229 15651 10287 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 11330 15688 11336 15700
rect 11291 15660 11336 15688
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 12802 15688 12808 15700
rect 12763 15660 12808 15688
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 16393 15691 16451 15697
rect 16393 15657 16405 15691
rect 16439 15688 16451 15691
rect 17034 15688 17040 15700
rect 16439 15660 17040 15688
rect 16439 15657 16451 15660
rect 16393 15651 16451 15657
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 17865 15691 17923 15697
rect 17865 15657 17877 15691
rect 17911 15688 17923 15691
rect 18414 15688 18420 15700
rect 17911 15660 18420 15688
rect 17911 15657 17923 15660
rect 17865 15651 17923 15657
rect 18414 15648 18420 15660
rect 18472 15648 18478 15700
rect 18506 15648 18512 15700
rect 18564 15688 18570 15700
rect 19334 15688 19340 15700
rect 18564 15660 18609 15688
rect 19295 15660 19340 15688
rect 18564 15648 18570 15660
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 21266 15648 21272 15700
rect 21324 15688 21330 15700
rect 21361 15691 21419 15697
rect 21361 15688 21373 15691
rect 21324 15660 21373 15688
rect 21324 15648 21330 15660
rect 21361 15657 21373 15660
rect 21407 15657 21419 15691
rect 21361 15651 21419 15657
rect 21726 15648 21732 15700
rect 21784 15648 21790 15700
rect 22462 15648 22468 15700
rect 22520 15688 22526 15700
rect 22922 15688 22928 15700
rect 22520 15660 22928 15688
rect 22520 15648 22526 15660
rect 22922 15648 22928 15660
rect 22980 15688 22986 15700
rect 23474 15688 23480 15700
rect 22980 15660 23480 15688
rect 22980 15648 22986 15660
rect 23474 15648 23480 15660
rect 23532 15648 23538 15700
rect 23842 15688 23848 15700
rect 23803 15660 23848 15688
rect 23842 15648 23848 15660
rect 23900 15648 23906 15700
rect 2056 15620 2084 15648
rect 4522 15620 4528 15632
rect 2056 15592 4528 15620
rect 4522 15580 4528 15592
rect 4580 15580 4586 15632
rect 6172 15623 6230 15629
rect 6172 15589 6184 15623
rect 6218 15620 6230 15623
rect 6270 15620 6276 15632
rect 6218 15592 6276 15620
rect 6218 15589 6230 15592
rect 6172 15583 6230 15589
rect 6270 15580 6276 15592
rect 6328 15580 6334 15632
rect 8481 15623 8539 15629
rect 8481 15589 8493 15623
rect 8527 15620 8539 15623
rect 8846 15620 8852 15632
rect 8527 15592 8852 15620
rect 8527 15589 8539 15592
rect 8481 15583 8539 15589
rect 8846 15580 8852 15592
rect 8904 15580 8910 15632
rect 11698 15629 11704 15632
rect 11692 15620 11704 15629
rect 11659 15592 11704 15620
rect 11692 15583 11704 15592
rect 11698 15580 11704 15583
rect 11756 15580 11762 15632
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 13725 15623 13783 15629
rect 13725 15620 13737 15623
rect 12492 15592 13737 15620
rect 12492 15580 12498 15592
rect 13725 15589 13737 15592
rect 13771 15589 13783 15623
rect 13725 15583 13783 15589
rect 20717 15623 20775 15629
rect 20717 15589 20729 15623
rect 20763 15620 20775 15623
rect 21744 15620 21772 15648
rect 20763 15592 21772 15620
rect 20763 15589 20775 15592
rect 20717 15583 20775 15589
rect 2038 15512 2044 15564
rect 2096 15552 2102 15564
rect 2225 15555 2283 15561
rect 2225 15552 2237 15555
rect 2096 15524 2237 15552
rect 2096 15512 2102 15524
rect 2225 15521 2237 15524
rect 2271 15521 2283 15555
rect 2225 15515 2283 15521
rect 2314 15512 2320 15564
rect 2372 15552 2378 15564
rect 3694 15552 3700 15564
rect 2372 15524 2417 15552
rect 3655 15524 3700 15552
rect 2372 15512 2378 15524
rect 3694 15512 3700 15524
rect 3752 15512 3758 15564
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 4982 15552 4988 15564
rect 4847 15524 4988 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 5902 15552 5908 15564
rect 5863 15524 5908 15552
rect 5902 15512 5908 15524
rect 5960 15512 5966 15564
rect 8570 15552 8576 15564
rect 8531 15524 8576 15552
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 10962 15552 10968 15564
rect 9364 15524 10968 15552
rect 9364 15512 9370 15524
rect 10962 15512 10968 15524
rect 11020 15552 11026 15564
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 11020 15524 11437 15552
rect 11020 15512 11026 15524
rect 11425 15521 11437 15524
rect 11471 15521 11483 15555
rect 13262 15552 13268 15564
rect 11425 15515 11483 15521
rect 11532 15524 13268 15552
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 2406 15484 2412 15496
rect 1811 15456 2412 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 3602 15444 3608 15496
rect 3660 15484 3666 15496
rect 4338 15484 4344 15496
rect 3660 15456 4344 15484
rect 3660 15444 3666 15456
rect 4338 15444 4344 15456
rect 4396 15484 4402 15496
rect 4893 15487 4951 15493
rect 4893 15484 4905 15487
rect 4396 15456 4905 15484
rect 4396 15444 4402 15456
rect 4893 15453 4905 15456
rect 4939 15484 4951 15487
rect 5442 15484 5448 15496
rect 4939 15456 5448 15484
rect 4939 15453 4951 15456
rect 4893 15447 4951 15453
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15484 10563 15487
rect 10778 15484 10784 15496
rect 10551 15456 10784 15484
rect 10551 15453 10563 15456
rect 10505 15447 10563 15453
rect 9125 15419 9183 15425
rect 9125 15385 9137 15419
rect 9171 15416 9183 15419
rect 9490 15416 9496 15428
rect 9171 15388 9496 15416
rect 9171 15385 9183 15388
rect 9125 15379 9183 15385
rect 9490 15376 9496 15388
rect 9548 15416 9554 15428
rect 10520 15416 10548 15447
rect 10778 15444 10784 15456
rect 10836 15484 10842 15496
rect 11532 15484 11560 15524
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 13909 15555 13967 15561
rect 13909 15521 13921 15555
rect 13955 15552 13967 15555
rect 13998 15552 14004 15564
rect 13955 15524 14004 15552
rect 13955 15521 13967 15524
rect 13909 15515 13967 15521
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 16758 15561 16764 15564
rect 16752 15515 16764 15561
rect 16816 15552 16822 15564
rect 16816 15524 16852 15552
rect 16758 15512 16764 15515
rect 16816 15512 16822 15524
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21801 15555 21859 15561
rect 21801 15552 21813 15555
rect 21140 15524 21813 15552
rect 21140 15512 21146 15524
rect 21801 15521 21813 15524
rect 21847 15521 21859 15555
rect 21801 15515 21859 15521
rect 23842 15512 23848 15564
rect 23900 15552 23906 15564
rect 24397 15555 24455 15561
rect 24397 15552 24409 15555
rect 23900 15524 24409 15552
rect 23900 15512 23906 15524
rect 24397 15521 24409 15524
rect 24443 15521 24455 15555
rect 24397 15515 24455 15521
rect 24489 15555 24547 15561
rect 24489 15521 24501 15555
rect 24535 15552 24547 15555
rect 24762 15552 24768 15564
rect 24535 15524 24768 15552
rect 24535 15521 24547 15524
rect 24489 15515 24547 15521
rect 24762 15512 24768 15524
rect 24820 15512 24826 15564
rect 15286 15484 15292 15496
rect 10836 15456 11560 15484
rect 15247 15456 15292 15484
rect 10836 15444 10842 15456
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 16206 15444 16212 15496
rect 16264 15484 16270 15496
rect 16485 15487 16543 15493
rect 16485 15484 16497 15487
rect 16264 15456 16497 15484
rect 16264 15444 16270 15456
rect 16485 15453 16497 15456
rect 16531 15453 16543 15487
rect 19426 15484 19432 15496
rect 19387 15456 19432 15484
rect 16485 15447 16543 15453
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 14090 15416 14096 15428
rect 9548 15388 10548 15416
rect 14051 15388 14096 15416
rect 9548 15376 9554 15388
rect 14090 15376 14096 15388
rect 14148 15376 14154 15428
rect 18877 15419 18935 15425
rect 18877 15385 18889 15419
rect 18923 15416 18935 15419
rect 19242 15416 19248 15428
rect 18923 15388 19248 15416
rect 18923 15385 18935 15388
rect 18877 15379 18935 15385
rect 19242 15376 19248 15388
rect 19300 15416 19306 15428
rect 19536 15416 19564 15447
rect 21358 15444 21364 15496
rect 21416 15484 21422 15496
rect 21545 15487 21603 15493
rect 21545 15484 21557 15487
rect 21416 15456 21557 15484
rect 21416 15444 21422 15456
rect 21545 15453 21557 15456
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 24673 15487 24731 15493
rect 24673 15453 24685 15487
rect 24719 15484 24731 15487
rect 25222 15484 25228 15496
rect 24719 15456 25228 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 19300 15388 19564 15416
rect 19300 15376 19306 15388
rect 7282 15348 7288 15360
rect 7243 15320 7288 15348
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 13354 15348 13360 15360
rect 13315 15320 13360 15348
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14369 15351 14427 15357
rect 14369 15348 14381 15351
rect 13872 15320 14381 15348
rect 13872 15308 13878 15320
rect 14369 15317 14381 15320
rect 14415 15348 14427 15351
rect 14458 15348 14464 15360
rect 14415 15320 14464 15348
rect 14415 15317 14427 15320
rect 14369 15311 14427 15317
rect 14458 15308 14464 15320
rect 14516 15308 14522 15360
rect 18966 15348 18972 15360
rect 18927 15320 18972 15348
rect 18966 15308 18972 15320
rect 19024 15308 19030 15360
rect 19978 15348 19984 15360
rect 19939 15320 19984 15348
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 24026 15348 24032 15360
rect 23987 15320 24032 15348
rect 24026 15308 24032 15320
rect 24084 15308 24090 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 4798 15104 4804 15156
rect 4856 15144 4862 15156
rect 4985 15147 5043 15153
rect 4985 15144 4997 15147
rect 4856 15116 4997 15144
rect 4856 15104 4862 15116
rect 4985 15113 4997 15116
rect 5031 15113 5043 15147
rect 4985 15107 5043 15113
rect 5994 15104 6000 15156
rect 6052 15144 6058 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 6052 15116 6193 15144
rect 6052 15104 6058 15116
rect 6181 15113 6193 15116
rect 6227 15113 6239 15147
rect 6181 15107 6239 15113
rect 2314 15036 2320 15088
rect 2372 15076 2378 15088
rect 3605 15079 3663 15085
rect 3605 15076 3617 15079
rect 2372 15048 3617 15076
rect 2372 15036 2378 15048
rect 3605 15045 3617 15048
rect 3651 15045 3663 15079
rect 6196 15076 6224 15107
rect 6270 15104 6276 15156
rect 6328 15144 6334 15156
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 6328 15116 6561 15144
rect 6328 15104 6334 15116
rect 6549 15113 6561 15116
rect 6595 15113 6607 15147
rect 7006 15144 7012 15156
rect 6967 15116 7012 15144
rect 6549 15107 6607 15113
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 9950 15144 9956 15156
rect 9911 15116 9956 15144
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 10318 15144 10324 15156
rect 10279 15116 10324 15144
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 10778 15144 10784 15156
rect 10739 15116 10784 15144
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11790 15104 11796 15116
rect 11848 15144 11854 15156
rect 12526 15144 12532 15156
rect 11848 15116 12532 15144
rect 11848 15104 11854 15116
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 12710 15144 12716 15156
rect 12671 15116 12716 15144
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 16945 15147 17003 15153
rect 16945 15144 16957 15147
rect 16816 15116 16957 15144
rect 16816 15104 16822 15116
rect 16945 15113 16957 15116
rect 16991 15144 17003 15147
rect 17586 15144 17592 15156
rect 16991 15116 17592 15144
rect 16991 15113 17003 15116
rect 16945 15107 17003 15113
rect 17586 15104 17592 15116
rect 17644 15144 17650 15156
rect 17773 15147 17831 15153
rect 17773 15144 17785 15147
rect 17644 15116 17785 15144
rect 17644 15104 17650 15116
rect 17773 15113 17785 15116
rect 17819 15113 17831 15147
rect 17773 15107 17831 15113
rect 7561 15079 7619 15085
rect 7561 15076 7573 15079
rect 6196 15048 7573 15076
rect 3605 15039 3663 15045
rect 7561 15045 7573 15048
rect 7607 15076 7619 15079
rect 7607 15048 7788 15076
rect 7607 15045 7619 15048
rect 7561 15039 7619 15045
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2498 15008 2504 15020
rect 1995 14980 2504 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2498 14968 2504 14980
rect 2556 14968 2562 15020
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 15008 2651 15011
rect 3145 15011 3203 15017
rect 3145 15008 3157 15011
rect 2639 14980 3157 15008
rect 2639 14977 2651 14980
rect 2593 14971 2651 14977
rect 3145 14977 3157 14980
rect 3191 15008 3203 15011
rect 3970 15008 3976 15020
rect 3191 14980 3976 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 2406 14900 2412 14952
rect 2464 14940 2470 14952
rect 2608 14940 2636 14971
rect 3970 14968 3976 14980
rect 4028 15008 4034 15020
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 4028 14980 4169 15008
rect 4028 14968 4034 14980
rect 4157 14977 4169 14980
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 4982 15008 4988 15020
rect 4755 14980 4988 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 4982 14968 4988 14980
rect 5040 14968 5046 15020
rect 5810 15008 5816 15020
rect 5771 14980 5816 15008
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 7760 15017 7788 15048
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 2464 14912 2636 14940
rect 2464 14900 2470 14912
rect 5166 14900 5172 14952
rect 5224 14940 5230 14952
rect 5537 14943 5595 14949
rect 5537 14940 5549 14943
rect 5224 14912 5549 14940
rect 5224 14900 5230 14912
rect 5537 14909 5549 14912
rect 5583 14909 5595 14943
rect 5537 14903 5595 14909
rect 5629 14943 5687 14949
rect 5629 14909 5641 14943
rect 5675 14940 5687 14943
rect 6822 14940 6828 14952
rect 5675 14912 6828 14940
rect 5675 14909 5687 14912
rect 5629 14903 5687 14909
rect 3973 14875 4031 14881
rect 3973 14872 3985 14875
rect 3528 14844 3985 14872
rect 3528 14816 3556 14844
rect 3973 14841 3985 14844
rect 4019 14841 4031 14875
rect 3973 14835 4031 14841
rect 4614 14832 4620 14884
rect 4672 14872 4678 14884
rect 4982 14872 4988 14884
rect 4672 14844 4988 14872
rect 4672 14832 4678 14844
rect 4982 14832 4988 14844
rect 5040 14832 5046 14884
rect 5258 14832 5264 14884
rect 5316 14872 5322 14884
rect 5644 14872 5672 14903
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7760 14940 7788 14971
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11241 15011 11299 15017
rect 11241 15008 11253 15011
rect 11112 14980 11253 15008
rect 11112 14968 11118 14980
rect 11241 14977 11253 14980
rect 11287 14977 11299 15011
rect 11241 14971 11299 14977
rect 11425 15011 11483 15017
rect 11425 14977 11437 15011
rect 11471 15008 11483 15011
rect 11698 15008 11704 15020
rect 11471 14980 11704 15008
rect 11471 14977 11483 14980
rect 11425 14971 11483 14977
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 13262 15008 13268 15020
rect 13223 14980 13268 15008
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 17788 15008 17816 15107
rect 19058 15104 19064 15156
rect 19116 15144 19122 15156
rect 19334 15144 19340 15156
rect 19116 15116 19340 15144
rect 19116 15104 19122 15116
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21082 15144 21088 15156
rect 21039 15116 21088 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 21082 15104 21088 15116
rect 21140 15144 21146 15156
rect 21913 15147 21971 15153
rect 21913 15144 21925 15147
rect 21140 15116 21925 15144
rect 21140 15104 21146 15116
rect 21913 15113 21925 15116
rect 21959 15113 21971 15147
rect 21913 15107 21971 15113
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22281 15147 22339 15153
rect 22281 15144 22293 15147
rect 22152 15116 22293 15144
rect 22152 15104 22158 15116
rect 22281 15113 22293 15116
rect 22327 15113 22339 15147
rect 22646 15144 22652 15156
rect 22607 15116 22652 15144
rect 22281 15107 22339 15113
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 23474 15144 23480 15156
rect 23435 15116 23480 15144
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 23842 15144 23848 15156
rect 23803 15116 23848 15144
rect 23842 15104 23848 15116
rect 23900 15104 23906 15156
rect 24670 15104 24676 15156
rect 24728 15144 24734 15156
rect 25593 15147 25651 15153
rect 25593 15144 25605 15147
rect 24728 15116 25605 15144
rect 24728 15104 24734 15116
rect 25593 15113 25605 15116
rect 25639 15113 25651 15147
rect 25593 15107 25651 15113
rect 18601 15011 18659 15017
rect 18601 15008 18613 15011
rect 17788 14980 18613 15008
rect 18601 14977 18613 14980
rect 18647 14977 18659 15011
rect 23492 15008 23520 15104
rect 24210 15036 24216 15088
rect 24268 15076 24274 15088
rect 24857 15079 24915 15085
rect 24857 15076 24869 15079
rect 24268 15048 24869 15076
rect 24268 15036 24274 15048
rect 24412 15020 24440 15048
rect 24857 15045 24869 15048
rect 24903 15045 24915 15079
rect 25222 15076 25228 15088
rect 25183 15048 25228 15076
rect 24857 15039 24915 15045
rect 25222 15036 25228 15048
rect 25280 15036 25286 15088
rect 24305 15011 24363 15017
rect 24305 15008 24317 15011
rect 23492 14980 24317 15008
rect 18601 14971 18659 14977
rect 24305 14977 24317 14980
rect 24351 14977 24363 15011
rect 24305 14971 24363 14977
rect 8846 14940 8852 14952
rect 7760 14912 8852 14940
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 14476 14912 14657 14940
rect 5316 14844 5672 14872
rect 5316 14832 5322 14844
rect 7834 14832 7840 14884
rect 7892 14872 7898 14884
rect 7990 14875 8048 14881
rect 7990 14872 8002 14875
rect 7892 14844 8002 14872
rect 7892 14832 7898 14844
rect 7990 14841 8002 14844
rect 8036 14841 8048 14875
rect 7990 14835 8048 14841
rect 12253 14875 12311 14881
rect 12253 14841 12265 14875
rect 12299 14872 12311 14875
rect 13170 14872 13176 14884
rect 12299 14844 13176 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 13446 14832 13452 14884
rect 13504 14872 13510 14884
rect 14476 14881 14504 14912
rect 14645 14909 14657 14912
rect 14691 14940 14703 14943
rect 16206 14940 16212 14952
rect 14691 14912 16212 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 16206 14900 16212 14912
rect 16264 14940 16270 14952
rect 16577 14943 16635 14949
rect 16577 14940 16589 14943
rect 16264 14912 16589 14940
rect 16264 14900 16270 14912
rect 16577 14909 16589 14912
rect 16623 14909 16635 14943
rect 16577 14903 16635 14909
rect 18230 14900 18236 14952
rect 18288 14940 18294 14952
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18288 14912 18521 14940
rect 18288 14900 18294 14912
rect 18509 14909 18521 14912
rect 18555 14940 18567 14943
rect 18966 14940 18972 14952
rect 18555 14912 18972 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 18966 14900 18972 14912
rect 19024 14900 19030 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 19444 14912 19625 14940
rect 14461 14875 14519 14881
rect 14461 14872 14473 14875
rect 13504 14844 14473 14872
rect 13504 14832 13510 14844
rect 14461 14841 14473 14844
rect 14507 14841 14519 14875
rect 14461 14835 14519 14841
rect 14550 14832 14556 14884
rect 14608 14872 14614 14884
rect 14890 14875 14948 14881
rect 14890 14872 14902 14875
rect 14608 14844 14902 14872
rect 14608 14832 14614 14844
rect 14890 14841 14902 14844
rect 14936 14841 14948 14875
rect 14890 14835 14948 14841
rect 17497 14875 17555 14881
rect 17497 14841 17509 14875
rect 17543 14872 17555 14875
rect 18417 14875 18475 14881
rect 18417 14872 18429 14875
rect 17543 14844 18429 14872
rect 17543 14841 17555 14844
rect 17497 14835 17555 14841
rect 18417 14841 18429 14844
rect 18463 14872 18475 14875
rect 18690 14872 18696 14884
rect 18463 14844 18696 14872
rect 18463 14841 18475 14844
rect 18417 14835 18475 14841
rect 18690 14832 18696 14844
rect 18748 14832 18754 14884
rect 19058 14872 19064 14884
rect 19019 14844 19064 14872
rect 19058 14832 19064 14844
rect 19116 14832 19122 14884
rect 2038 14804 2044 14816
rect 1999 14776 2044 14804
rect 2038 14764 2044 14776
rect 2096 14764 2102 14816
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 2498 14804 2504 14816
rect 2455 14776 2504 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 3510 14804 3516 14816
rect 3471 14776 3516 14804
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 4062 14804 4068 14816
rect 4023 14776 4068 14804
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 5074 14764 5080 14816
rect 5132 14804 5138 14816
rect 5169 14807 5227 14813
rect 5169 14804 5181 14807
rect 5132 14776 5181 14804
rect 5132 14764 5138 14776
rect 5169 14773 5181 14776
rect 5215 14773 5227 14807
rect 5169 14767 5227 14773
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 6546 14804 6552 14816
rect 6420 14776 6552 14804
rect 6420 14764 6426 14776
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 9125 14807 9183 14813
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9214 14804 9220 14816
rect 9171 14776 9220 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 10597 14807 10655 14813
rect 10597 14804 10609 14807
rect 10192 14776 10609 14804
rect 10192 14764 10198 14776
rect 10597 14773 10609 14776
rect 10643 14804 10655 14807
rect 11149 14807 11207 14813
rect 11149 14804 11161 14807
rect 10643 14776 11161 14804
rect 10643 14773 10655 14776
rect 10597 14767 10655 14773
rect 11149 14773 11161 14776
rect 11195 14773 11207 14807
rect 11149 14767 11207 14773
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 12768 14776 13093 14804
rect 12768 14764 12774 14776
rect 13081 14773 13093 14776
rect 13127 14773 13139 14807
rect 13998 14804 14004 14816
rect 13959 14776 14004 14804
rect 13081 14767 13139 14773
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 16025 14807 16083 14813
rect 16025 14773 16037 14807
rect 16071 14804 16083 14807
rect 16390 14804 16396 14816
rect 16071 14776 16396 14804
rect 16071 14773 16083 14776
rect 16025 14767 16083 14773
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 18046 14804 18052 14816
rect 18007 14776 18052 14804
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18322 14764 18328 14816
rect 18380 14804 18386 14816
rect 19444 14813 19472 14912
rect 19613 14909 19625 14912
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 21266 14900 21272 14952
rect 21324 14940 21330 14952
rect 22465 14943 22523 14949
rect 22465 14940 22477 14943
rect 21324 14912 22477 14940
rect 21324 14900 21330 14912
rect 22465 14909 22477 14912
rect 22511 14940 22523 14943
rect 23017 14943 23075 14949
rect 23017 14940 23029 14943
rect 22511 14912 23029 14940
rect 22511 14909 22523 14912
rect 22465 14903 22523 14909
rect 23017 14909 23029 14912
rect 23063 14909 23075 14943
rect 23017 14903 23075 14909
rect 23934 14900 23940 14952
rect 23992 14940 23998 14952
rect 24213 14943 24271 14949
rect 24213 14940 24225 14943
rect 23992 14912 24225 14940
rect 23992 14900 23998 14912
rect 24213 14909 24225 14912
rect 24259 14909 24271 14943
rect 24320 14940 24348 14971
rect 24394 14968 24400 15020
rect 24452 15008 24458 15020
rect 24452 14980 24545 15008
rect 24452 14968 24458 14980
rect 25409 14943 25467 14949
rect 25409 14940 25421 14943
rect 24320 14912 25421 14940
rect 24213 14903 24271 14909
rect 25409 14909 25421 14912
rect 25455 14940 25467 14943
rect 25961 14943 26019 14949
rect 25961 14940 25973 14943
rect 25455 14912 25973 14940
rect 25455 14909 25467 14912
rect 25409 14903 25467 14909
rect 25961 14909 25973 14912
rect 26007 14909 26019 14943
rect 25961 14903 26019 14909
rect 19880 14875 19938 14881
rect 19880 14841 19892 14875
rect 19926 14872 19938 14875
rect 19978 14872 19984 14884
rect 19926 14844 19984 14872
rect 19926 14841 19938 14844
rect 19880 14835 19938 14841
rect 19978 14832 19984 14844
rect 20036 14832 20042 14884
rect 19429 14807 19487 14813
rect 19429 14804 19441 14807
rect 18380 14776 19441 14804
rect 18380 14764 18386 14776
rect 19429 14773 19441 14776
rect 19475 14773 19487 14807
rect 19429 14767 19487 14773
rect 20898 14764 20904 14816
rect 20956 14804 20962 14816
rect 21358 14804 21364 14816
rect 20956 14776 21364 14804
rect 20956 14764 20962 14776
rect 21358 14764 21364 14776
rect 21416 14804 21422 14816
rect 21545 14807 21603 14813
rect 21545 14804 21557 14807
rect 21416 14776 21557 14804
rect 21416 14764 21422 14776
rect 21545 14773 21557 14776
rect 21591 14773 21603 14807
rect 21545 14767 21603 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2130 14560 2136 14612
rect 2188 14600 2194 14612
rect 2409 14603 2467 14609
rect 2409 14600 2421 14603
rect 2188 14572 2421 14600
rect 2188 14560 2194 14572
rect 2409 14569 2421 14572
rect 2455 14569 2467 14603
rect 2409 14563 2467 14569
rect 2590 14560 2596 14612
rect 2648 14600 2654 14612
rect 2869 14603 2927 14609
rect 2869 14600 2881 14603
rect 2648 14572 2881 14600
rect 2648 14560 2654 14572
rect 2869 14569 2881 14572
rect 2915 14569 2927 14603
rect 2869 14563 2927 14569
rect 3697 14603 3755 14609
rect 3697 14569 3709 14603
rect 3743 14600 3755 14603
rect 3970 14600 3976 14612
rect 3743 14572 3976 14600
rect 3743 14569 3755 14572
rect 3697 14563 3755 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4709 14603 4767 14609
rect 4709 14600 4721 14603
rect 4212 14572 4721 14600
rect 4212 14560 4218 14572
rect 4709 14569 4721 14572
rect 4755 14569 4767 14603
rect 6270 14600 6276 14612
rect 6231 14572 6276 14600
rect 4709 14563 4767 14569
rect 6270 14560 6276 14572
rect 6328 14600 6334 14612
rect 7006 14600 7012 14612
rect 6328 14572 7012 14600
rect 6328 14560 6334 14572
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 9490 14600 9496 14612
rect 9451 14572 9496 14600
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 11698 14600 11704 14612
rect 11659 14572 11704 14600
rect 11698 14560 11704 14572
rect 11756 14600 11762 14612
rect 11977 14603 12035 14609
rect 11977 14600 11989 14603
rect 11756 14572 11989 14600
rect 11756 14560 11762 14572
rect 11977 14569 11989 14572
rect 12023 14569 12035 14603
rect 12342 14600 12348 14612
rect 12303 14572 12348 14600
rect 11977 14563 12035 14569
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 13262 14600 13268 14612
rect 13219 14572 13268 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 13814 14600 13820 14612
rect 13679 14572 13820 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 17586 14600 17592 14612
rect 17547 14572 17592 14600
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 18230 14600 18236 14612
rect 18191 14572 18236 14600
rect 18230 14560 18236 14572
rect 18288 14560 18294 14612
rect 18690 14600 18696 14612
rect 18651 14572 18696 14600
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 20714 14600 20720 14612
rect 20675 14572 20720 14600
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 23845 14603 23903 14609
rect 23845 14569 23857 14603
rect 23891 14600 23903 14603
rect 24762 14600 24768 14612
rect 23891 14572 24768 14600
rect 23891 14569 23903 14572
rect 23845 14563 23903 14569
rect 24762 14560 24768 14572
rect 24820 14600 24826 14612
rect 24857 14603 24915 14609
rect 24857 14600 24869 14603
rect 24820 14572 24869 14600
rect 24820 14560 24826 14572
rect 24857 14569 24869 14572
rect 24903 14569 24915 14603
rect 24857 14563 24915 14569
rect 25593 14603 25651 14609
rect 25593 14569 25605 14603
rect 25639 14600 25651 14603
rect 25682 14600 25688 14612
rect 25639 14572 25688 14600
rect 25639 14569 25651 14572
rect 25593 14563 25651 14569
rect 25682 14560 25688 14572
rect 25740 14560 25746 14612
rect 4338 14532 4344 14544
rect 4299 14504 4344 14532
rect 4338 14492 4344 14504
rect 4396 14492 4402 14544
rect 19518 14532 19524 14544
rect 19168 14504 19524 14532
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14433 1455 14467
rect 1397 14427 1455 14433
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14464 2835 14467
rect 3142 14464 3148 14476
rect 2823 14436 3148 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 1412 14328 1440 14427
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 5074 14464 5080 14476
rect 4672 14436 5080 14464
rect 4672 14424 4678 14436
rect 5074 14424 5080 14436
rect 5132 14464 5138 14476
rect 5261 14467 5319 14473
rect 5261 14464 5273 14467
rect 5132 14436 5273 14464
rect 5132 14424 5138 14436
rect 5261 14433 5273 14436
rect 5307 14433 5319 14467
rect 5261 14427 5319 14433
rect 6270 14424 6276 14476
rect 6328 14464 6334 14476
rect 6713 14467 6771 14473
rect 6713 14464 6725 14467
rect 6328 14436 6725 14464
rect 6328 14424 6334 14436
rect 6713 14433 6725 14436
rect 6759 14464 6771 14467
rect 7282 14464 7288 14476
rect 6759 14436 7288 14464
rect 6759 14433 6771 14436
rect 6713 14427 6771 14433
rect 7282 14424 7288 14436
rect 7340 14424 7346 14476
rect 8754 14424 8760 14476
rect 8812 14464 8818 14476
rect 9944 14467 10002 14473
rect 9944 14464 9956 14467
rect 8812 14436 9956 14464
rect 8812 14424 8818 14436
rect 9944 14433 9956 14436
rect 9990 14464 10002 14467
rect 11514 14464 11520 14476
rect 9990 14436 11520 14464
rect 9990 14433 10002 14436
rect 9944 14427 10002 14433
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 12066 14424 12072 14476
rect 12124 14464 12130 14476
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 12124 14436 12173 14464
rect 12124 14424 12130 14436
rect 12161 14433 12173 14436
rect 12207 14433 12219 14467
rect 12161 14427 12219 14433
rect 13354 14424 13360 14476
rect 13412 14464 13418 14476
rect 14001 14467 14059 14473
rect 14001 14464 14013 14467
rect 13412 14436 14013 14464
rect 13412 14424 13418 14436
rect 14001 14433 14013 14436
rect 14047 14464 14059 14467
rect 14458 14464 14464 14476
rect 14047 14436 14464 14464
rect 14047 14433 14059 14436
rect 14001 14427 14059 14433
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 16206 14464 16212 14476
rect 16167 14436 16212 14464
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 16482 14473 16488 14476
rect 16476 14464 16488 14473
rect 16443 14436 16488 14464
rect 16476 14427 16488 14436
rect 16482 14424 16488 14427
rect 16540 14424 16546 14476
rect 19058 14464 19064 14476
rect 19019 14436 19064 14464
rect 19058 14424 19064 14436
rect 19116 14424 19122 14476
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2961 14399 3019 14405
rect 2961 14396 2973 14399
rect 2464 14368 2973 14396
rect 2464 14356 2470 14368
rect 2961 14365 2973 14368
rect 3007 14396 3019 14399
rect 3602 14396 3608 14408
rect 3007 14368 3608 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 3602 14356 3608 14368
rect 3660 14356 3666 14408
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14365 5411 14399
rect 5353 14359 5411 14365
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14396 5503 14399
rect 5534 14396 5540 14408
rect 5491 14368 5540 14396
rect 5491 14365 5503 14368
rect 5445 14359 5503 14365
rect 1762 14328 1768 14340
rect 1412 14300 1768 14328
rect 1762 14288 1768 14300
rect 1820 14328 1826 14340
rect 4893 14331 4951 14337
rect 4893 14328 4905 14331
rect 1820 14300 4905 14328
rect 1820 14288 1826 14300
rect 4893 14297 4905 14300
rect 4939 14297 4951 14331
rect 4893 14291 4951 14297
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 5368 14328 5396 14359
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5994 14356 6000 14408
rect 6052 14396 6058 14408
rect 6362 14396 6368 14408
rect 6052 14368 6368 14396
rect 6052 14356 6058 14368
rect 6362 14356 6368 14368
rect 6420 14396 6426 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6420 14368 6469 14396
rect 6420 14356 6426 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 8904 14368 9689 14396
rect 8904 14356 8910 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 12986 14356 12992 14408
rect 13044 14396 13050 14408
rect 13722 14396 13728 14408
rect 13044 14368 13728 14396
rect 13044 14356 13050 14368
rect 13722 14356 13728 14368
rect 13780 14396 13786 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13780 14368 14105 14396
rect 13780 14356 13786 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 14182 14356 14188 14408
rect 14240 14396 14246 14408
rect 14240 14368 14285 14396
rect 14240 14356 14246 14368
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 19168 14405 19196 14504
rect 19518 14492 19524 14504
rect 19576 14492 19582 14544
rect 21082 14492 21088 14544
rect 21140 14541 21146 14544
rect 21140 14535 21204 14541
rect 21140 14501 21158 14535
rect 21192 14501 21204 14535
rect 21140 14495 21204 14501
rect 21140 14492 21146 14495
rect 23658 14492 23664 14544
rect 23716 14532 23722 14544
rect 24213 14535 24271 14541
rect 24213 14532 24225 14535
rect 23716 14504 24225 14532
rect 23716 14492 23722 14504
rect 24213 14501 24225 14504
rect 24259 14501 24271 14535
rect 24213 14495 24271 14501
rect 22278 14424 22284 14476
rect 22336 14424 22342 14476
rect 23385 14467 23443 14473
rect 23385 14433 23397 14467
rect 23431 14464 23443 14467
rect 23842 14464 23848 14476
rect 23431 14436 23848 14464
rect 23431 14433 23443 14436
rect 23385 14427 23443 14433
rect 23842 14424 23848 14436
rect 23900 14424 23906 14476
rect 25130 14424 25136 14476
rect 25188 14464 25194 14476
rect 25409 14467 25467 14473
rect 25409 14464 25421 14467
rect 25188 14436 25421 14464
rect 25188 14424 25194 14436
rect 25409 14433 25421 14436
rect 25455 14433 25467 14467
rect 25409 14427 25467 14433
rect 19153 14399 19211 14405
rect 19153 14396 19165 14399
rect 18472 14368 19165 14396
rect 18472 14356 18478 14368
rect 19153 14365 19165 14368
rect 19199 14365 19211 14399
rect 19153 14359 19211 14365
rect 19242 14356 19248 14408
rect 19300 14396 19306 14408
rect 20898 14396 20904 14408
rect 19300 14368 19345 14396
rect 20859 14368 20904 14396
rect 19300 14356 19306 14368
rect 20898 14356 20904 14368
rect 20956 14356 20962 14408
rect 22296 14396 22324 14424
rect 23474 14396 23480 14408
rect 22296 14368 23480 14396
rect 23474 14356 23480 14368
rect 23532 14396 23538 14408
rect 24302 14396 24308 14408
rect 23532 14368 24308 14396
rect 23532 14356 23538 14368
rect 24302 14356 24308 14368
rect 24360 14356 24366 14408
rect 24394 14356 24400 14408
rect 24452 14396 24458 14408
rect 24452 14368 24497 14396
rect 24452 14356 24458 14368
rect 5132 14300 5396 14328
rect 5132 14288 5138 14300
rect 5810 14288 5816 14340
rect 5868 14328 5874 14340
rect 5905 14331 5963 14337
rect 5905 14328 5917 14331
rect 5868 14300 5917 14328
rect 5868 14288 5874 14300
rect 5905 14297 5917 14300
rect 5951 14328 5963 14331
rect 6270 14328 6276 14340
rect 5951 14300 6276 14328
rect 5951 14297 5963 14300
rect 5905 14291 5963 14297
rect 6270 14288 6276 14300
rect 6328 14288 6334 14340
rect 7834 14328 7840 14340
rect 7795 14300 7840 14328
rect 7834 14288 7840 14300
rect 7892 14328 7898 14340
rect 8389 14331 8447 14337
rect 8389 14328 8401 14331
rect 7892 14300 8401 14328
rect 7892 14288 7898 14300
rect 8389 14297 8401 14300
rect 8435 14297 8447 14331
rect 22278 14328 22284 14340
rect 22239 14300 22284 14328
rect 8389 14291 8447 14297
rect 22278 14288 22284 14300
rect 22336 14288 22342 14340
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 1670 14260 1676 14272
rect 1627 14232 1676 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 2133 14263 2191 14269
rect 2133 14229 2145 14263
rect 2179 14260 2191 14263
rect 2498 14260 2504 14272
rect 2179 14232 2504 14260
rect 2179 14229 2191 14232
rect 2133 14223 2191 14229
rect 2498 14220 2504 14232
rect 2556 14260 2562 14272
rect 6086 14260 6092 14272
rect 2556 14232 6092 14260
rect 2556 14220 2562 14232
rect 6086 14220 6092 14232
rect 6144 14260 6150 14272
rect 7098 14260 7104 14272
rect 6144 14232 7104 14260
rect 6144 14220 6150 14232
rect 7098 14220 7104 14232
rect 7156 14220 7162 14272
rect 9122 14260 9128 14272
rect 9083 14232 9128 14260
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 11054 14260 11060 14272
rect 11015 14232 11060 14260
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 12710 14260 12716 14272
rect 12671 14232 12716 14260
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 13446 14260 13452 14272
rect 13407 14232 13452 14260
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 14550 14220 14556 14272
rect 14608 14260 14614 14272
rect 14645 14263 14703 14269
rect 14645 14260 14657 14263
rect 14608 14232 14657 14260
rect 14608 14220 14614 14232
rect 14645 14229 14657 14232
rect 14691 14229 14703 14263
rect 16022 14260 16028 14272
rect 15983 14232 16028 14260
rect 14645 14223 14703 14229
rect 16022 14220 16028 14232
rect 16080 14220 16086 14272
rect 18601 14263 18659 14269
rect 18601 14229 18613 14263
rect 18647 14260 18659 14263
rect 18690 14260 18696 14272
rect 18647 14232 18696 14260
rect 18647 14229 18659 14232
rect 18601 14223 18659 14229
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 19702 14260 19708 14272
rect 19663 14232 19708 14260
rect 19702 14220 19708 14232
rect 19760 14220 19766 14272
rect 23017 14263 23075 14269
rect 23017 14229 23029 14263
rect 23063 14260 23075 14263
rect 23106 14260 23112 14272
rect 23063 14232 23112 14260
rect 23063 14229 23075 14232
rect 23017 14223 23075 14229
rect 23106 14220 23112 14232
rect 23164 14220 23170 14272
rect 23750 14260 23756 14272
rect 23711 14232 23756 14260
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 2682 14056 2688 14068
rect 2643 14028 2688 14056
rect 2682 14016 2688 14028
rect 2740 14016 2746 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 6457 14059 6515 14065
rect 6457 14056 6469 14059
rect 6420 14028 6469 14056
rect 6420 14016 6426 14028
rect 6457 14025 6469 14028
rect 6503 14025 6515 14059
rect 6457 14019 6515 14025
rect 7374 14016 7380 14068
rect 7432 14056 7438 14068
rect 7469 14059 7527 14065
rect 7469 14056 7481 14059
rect 7432 14028 7481 14056
rect 7432 14016 7438 14028
rect 7469 14025 7481 14028
rect 7515 14056 7527 14059
rect 8478 14056 8484 14068
rect 7515 14028 8484 14056
rect 7515 14025 7527 14028
rect 7469 14019 7527 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 8846 14016 8852 14068
rect 8904 14056 8910 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 8904 14028 9045 14056
rect 8904 14016 8910 14028
rect 9033 14025 9045 14028
rect 9079 14056 9091 14059
rect 9309 14059 9367 14065
rect 9309 14056 9321 14059
rect 9079 14028 9321 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 9309 14025 9321 14028
rect 9355 14056 9367 14059
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 9355 14028 9413 14056
rect 9355 14025 9367 14028
rect 9309 14019 9367 14025
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 11514 14056 11520 14068
rect 11475 14028 11520 14056
rect 9401 14019 9459 14025
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 12986 14056 12992 14068
rect 12947 14028 12992 14056
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 13354 14056 13360 14068
rect 13315 14028 13360 14056
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 15841 14059 15899 14065
rect 15841 14025 15853 14059
rect 15887 14056 15899 14059
rect 16482 14056 16488 14068
rect 15887 14028 16488 14056
rect 15887 14025 15899 14028
rect 15841 14019 15899 14025
rect 16482 14016 16488 14028
rect 16540 14056 16546 14068
rect 17865 14059 17923 14065
rect 17865 14056 17877 14059
rect 16540 14028 17877 14056
rect 16540 14016 16546 14028
rect 17865 14025 17877 14028
rect 17911 14056 17923 14059
rect 19242 14056 19248 14068
rect 17911 14028 19248 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 21266 14056 21272 14068
rect 21227 14028 21272 14056
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 21453 14059 21511 14065
rect 21453 14025 21465 14059
rect 21499 14056 21511 14059
rect 23106 14056 23112 14068
rect 21499 14028 23112 14056
rect 21499 14025 21511 14028
rect 21453 14019 21511 14025
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 23474 14056 23480 14068
rect 23435 14028 23480 14056
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 2041 13991 2099 13997
rect 2041 13957 2053 13991
rect 2087 13988 2099 13991
rect 2590 13988 2596 14000
rect 2087 13960 2596 13988
rect 2087 13957 2099 13960
rect 2041 13951 2099 13957
rect 2590 13948 2596 13960
rect 2648 13948 2654 14000
rect 5166 13988 5172 14000
rect 5127 13960 5172 13988
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 8021 13991 8079 13997
rect 8021 13957 8033 13991
rect 8067 13988 8079 13991
rect 8202 13988 8208 14000
rect 8067 13960 8208 13988
rect 8067 13957 8079 13960
rect 8021 13951 8079 13957
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 14550 13948 14556 14000
rect 14608 13988 14614 14000
rect 14829 13991 14887 13997
rect 14829 13988 14841 13991
rect 14608 13960 14841 13988
rect 14608 13948 14614 13960
rect 14829 13957 14841 13960
rect 14875 13957 14887 13991
rect 14829 13951 14887 13957
rect 16206 13948 16212 14000
rect 16264 13988 16270 14000
rect 16850 13988 16856 14000
rect 16264 13960 16856 13988
rect 16264 13948 16270 13960
rect 16850 13948 16856 13960
rect 16908 13988 16914 14000
rect 16945 13991 17003 13997
rect 16945 13988 16957 13991
rect 16908 13960 16957 13988
rect 16908 13948 16914 13960
rect 16945 13957 16957 13960
rect 16991 13957 17003 13991
rect 19978 13988 19984 14000
rect 19939 13960 19984 13988
rect 16945 13951 17003 13957
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 1670 13920 1676 13932
rect 1412 13892 1676 13920
rect 1412 13861 1440 13892
rect 1670 13880 1676 13892
rect 1728 13920 1734 13932
rect 2682 13920 2688 13932
rect 1728 13892 2688 13920
rect 1728 13880 1734 13892
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13920 3479 13923
rect 3878 13920 3884 13932
rect 3467 13892 3884 13920
rect 3467 13889 3479 13892
rect 3421 13883 3479 13889
rect 3878 13880 3884 13892
rect 3936 13920 3942 13932
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 3936 13892 4169 13920
rect 3936 13880 3942 13892
rect 4157 13889 4169 13892
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 6178 13920 6184 13932
rect 5859 13892 6184 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 8665 13923 8723 13929
rect 8665 13920 8677 13923
rect 8168 13892 8677 13920
rect 8168 13880 8174 13892
rect 8665 13889 8677 13892
rect 8711 13920 8723 13923
rect 8754 13920 8760 13932
rect 8711 13892 8760 13920
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9122 13880 9128 13932
rect 9180 13920 9186 13932
rect 9180 13892 9720 13920
rect 9180 13880 9186 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13821 1455 13855
rect 1397 13815 1455 13821
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 4709 13855 4767 13861
rect 2547 13824 3188 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 3160 13793 3188 13824
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 7834 13852 7840 13864
rect 4755 13824 5488 13852
rect 7795 13824 7840 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 3145 13787 3203 13793
rect 3145 13753 3157 13787
rect 3191 13784 3203 13787
rect 3510 13784 3516 13796
rect 3191 13756 3516 13784
rect 3191 13753 3203 13756
rect 3145 13747 3203 13753
rect 3510 13744 3516 13756
rect 3568 13744 3574 13796
rect 3878 13744 3884 13796
rect 3936 13784 3942 13796
rect 4065 13787 4123 13793
rect 4065 13784 4077 13787
rect 3936 13756 4077 13784
rect 3936 13744 3942 13756
rect 4065 13753 4077 13756
rect 4111 13753 4123 13787
rect 5460 13784 5488 13824
rect 7834 13812 7840 13824
rect 7892 13852 7898 13864
rect 8478 13852 8484 13864
rect 7892 13824 8248 13852
rect 8439 13824 8484 13852
rect 7892 13812 7898 13824
rect 5537 13787 5595 13793
rect 5537 13784 5549 13787
rect 5460 13756 5549 13784
rect 4065 13747 4123 13753
rect 5537 13753 5549 13756
rect 5583 13784 5595 13787
rect 6825 13787 6883 13793
rect 6825 13784 6837 13787
rect 5583 13756 6837 13784
rect 5583 13753 5595 13756
rect 5537 13747 5595 13753
rect 6825 13753 6837 13756
rect 6871 13753 6883 13787
rect 8220 13784 8248 13824
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 9309 13855 9367 13861
rect 9309 13821 9321 13855
rect 9355 13852 9367 13855
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9355 13824 9597 13852
rect 9355 13821 9367 13824
rect 9309 13815 9367 13821
rect 9585 13821 9597 13824
rect 9631 13821 9643 13855
rect 9692 13852 9720 13892
rect 16022 13880 16028 13932
rect 16080 13920 16086 13932
rect 16485 13923 16543 13929
rect 16485 13920 16497 13923
rect 16080 13892 16497 13920
rect 16080 13880 16086 13892
rect 16485 13889 16497 13892
rect 16531 13889 16543 13923
rect 20898 13920 20904 13932
rect 16485 13883 16543 13889
rect 19628 13892 20904 13920
rect 9852 13855 9910 13861
rect 9852 13852 9864 13855
rect 9692 13824 9864 13852
rect 9585 13815 9643 13821
rect 9852 13821 9864 13824
rect 9898 13852 9910 13855
rect 10134 13852 10140 13864
rect 9898 13824 10140 13852
rect 9898 13821 9910 13824
rect 9852 13815 9910 13821
rect 8389 13787 8447 13793
rect 8389 13784 8401 13787
rect 8220 13756 8401 13784
rect 6825 13747 6883 13753
rect 8389 13753 8401 13756
rect 8435 13753 8447 13787
rect 9600 13784 9628 13815
rect 10134 13812 10140 13824
rect 10192 13852 10198 13864
rect 11054 13852 11060 13864
rect 10192 13824 11060 13852
rect 10192 13812 10198 13824
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 13446 13852 13452 13864
rect 12584 13824 13452 13852
rect 12584 13812 12590 13824
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 15378 13852 15384 13864
rect 15339 13824 15384 13852
rect 15378 13812 15384 13824
rect 15436 13852 15442 13864
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 15436 13824 16405 13852
rect 15436 13812 15442 13824
rect 16393 13821 16405 13824
rect 16439 13821 16451 13855
rect 16393 13815 16451 13821
rect 18322 13812 18328 13864
rect 18380 13852 18386 13864
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18380 13824 18613 13852
rect 18380 13812 18386 13824
rect 18601 13821 18613 13824
rect 18647 13852 18659 13855
rect 19628 13852 19656 13892
rect 20898 13880 20904 13892
rect 20956 13880 20962 13932
rect 21284 13920 21312 14016
rect 22922 13948 22928 14000
rect 22980 13988 22986 14000
rect 23017 13991 23075 13997
rect 23017 13988 23029 13991
rect 22980 13960 23029 13988
rect 22980 13948 22986 13960
rect 23017 13957 23029 13960
rect 23063 13957 23075 13991
rect 23661 13991 23719 13997
rect 23661 13988 23673 13991
rect 23017 13951 23075 13957
rect 23124 13960 23673 13988
rect 21913 13923 21971 13929
rect 21913 13920 21925 13923
rect 21284 13892 21925 13920
rect 21913 13889 21925 13892
rect 21959 13889 21971 13923
rect 21913 13883 21971 13889
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 18647 13824 19656 13852
rect 22020 13852 22048 13883
rect 22830 13880 22836 13932
rect 22888 13920 22894 13932
rect 23124 13920 23152 13960
rect 23661 13957 23673 13960
rect 23707 13957 23719 13991
rect 23661 13951 23719 13957
rect 22888 13892 23152 13920
rect 22888 13880 22894 13892
rect 23382 13880 23388 13932
rect 23440 13920 23446 13932
rect 23750 13920 23756 13932
rect 23440 13892 23756 13920
rect 23440 13880 23446 13892
rect 23750 13880 23756 13892
rect 23808 13920 23814 13932
rect 24213 13923 24271 13929
rect 24213 13920 24225 13923
rect 23808 13892 24225 13920
rect 23808 13880 23814 13892
rect 24213 13889 24225 13892
rect 24259 13889 24271 13923
rect 24213 13883 24271 13889
rect 25130 13880 25136 13932
rect 25188 13920 25194 13932
rect 26145 13923 26203 13929
rect 26145 13920 26157 13923
rect 25188 13892 26157 13920
rect 25188 13880 25194 13892
rect 26145 13889 26157 13892
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 22020 13824 22508 13852
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 9950 13784 9956 13796
rect 9600 13756 9956 13784
rect 8389 13747 8447 13753
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 12158 13784 12164 13796
rect 12119 13756 12164 13784
rect 12158 13744 12164 13756
rect 12216 13784 12222 13796
rect 13694 13787 13752 13793
rect 13694 13784 13706 13787
rect 12216 13756 13706 13784
rect 12216 13744 12222 13756
rect 13694 13753 13706 13756
rect 13740 13784 13752 13787
rect 13814 13784 13820 13796
rect 13740 13756 13820 13784
rect 13740 13753 13752 13756
rect 13694 13747 13752 13753
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 18414 13784 18420 13796
rect 15764 13756 18420 13784
rect 3602 13716 3608 13728
rect 3563 13688 3608 13716
rect 3602 13676 3608 13688
rect 3660 13676 3666 13728
rect 3970 13716 3976 13728
rect 3931 13688 3976 13716
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4982 13716 4988 13728
rect 4943 13688 4988 13716
rect 4982 13676 4988 13688
rect 5040 13716 5046 13728
rect 5629 13719 5687 13725
rect 5629 13716 5641 13719
rect 5040 13688 5641 13716
rect 5040 13676 5046 13688
rect 5629 13685 5641 13688
rect 5675 13685 5687 13719
rect 10962 13716 10968 13728
rect 10923 13688 10968 13716
rect 5629 13679 5687 13685
rect 10962 13676 10968 13688
rect 11020 13676 11026 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12492 13688 12537 13716
rect 12492 13676 12498 13688
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 15764 13716 15792 13756
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 18690 13744 18696 13796
rect 18748 13784 18754 13796
rect 18846 13787 18904 13793
rect 18846 13784 18858 13787
rect 18748 13756 18858 13784
rect 18748 13744 18754 13756
rect 18846 13753 18858 13756
rect 18892 13753 18904 13787
rect 18846 13747 18904 13753
rect 22480 13728 22508 13824
rect 23106 13812 23112 13864
rect 23164 13852 23170 13864
rect 24121 13855 24179 13861
rect 23164 13824 23428 13852
rect 23164 13812 23170 13824
rect 23400 13784 23428 13824
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 24302 13852 24308 13864
rect 24167 13824 24308 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 24302 13812 24308 13824
rect 24360 13852 24366 13864
rect 25041 13855 25099 13861
rect 25041 13852 25053 13855
rect 24360 13824 25053 13852
rect 24360 13812 24366 13824
rect 25041 13821 25053 13824
rect 25087 13821 25099 13855
rect 25222 13852 25228 13864
rect 25183 13824 25228 13852
rect 25041 13815 25099 13821
rect 25222 13812 25228 13824
rect 25280 13852 25286 13864
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25280 13824 25789 13852
rect 25280 13812 25286 13824
rect 25777 13821 25789 13824
rect 25823 13821 25835 13855
rect 25777 13815 25835 13821
rect 24029 13787 24087 13793
rect 24029 13784 24041 13787
rect 23400 13756 24041 13784
rect 24029 13753 24041 13756
rect 24075 13753 24087 13787
rect 24029 13747 24087 13753
rect 15930 13716 15936 13728
rect 12768 13688 15792 13716
rect 15891 13688 15936 13716
rect 12768 13676 12774 13688
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16298 13716 16304 13728
rect 16259 13688 16304 13716
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 20625 13719 20683 13725
rect 20625 13685 20637 13719
rect 20671 13716 20683 13719
rect 21821 13719 21879 13725
rect 21821 13716 21833 13719
rect 20671 13688 21833 13716
rect 20671 13685 20683 13688
rect 20625 13679 20683 13685
rect 21821 13685 21833 13688
rect 21867 13716 21879 13719
rect 22094 13716 22100 13728
rect 21867 13688 22100 13716
rect 21867 13685 21879 13688
rect 21821 13679 21879 13685
rect 22094 13676 22100 13688
rect 22152 13676 22158 13728
rect 22462 13716 22468 13728
rect 22423 13688 22468 13716
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 23658 13676 23664 13728
rect 23716 13716 23722 13728
rect 24673 13719 24731 13725
rect 24673 13716 24685 13719
rect 23716 13688 24685 13716
rect 23716 13676 23722 13688
rect 24673 13685 24685 13688
rect 24719 13685 24731 13719
rect 25406 13716 25412 13728
rect 25367 13688 25412 13716
rect 24673 13679 24731 13685
rect 25406 13676 25412 13688
rect 25464 13676 25470 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 1946 13512 1952 13524
rect 1907 13484 1952 13512
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 2314 13512 2320 13524
rect 2275 13484 2320 13512
rect 2314 13472 2320 13484
rect 2372 13472 2378 13524
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 3605 13515 3663 13521
rect 3605 13512 3617 13515
rect 2924 13484 3617 13512
rect 2924 13472 2930 13484
rect 3605 13481 3617 13484
rect 3651 13512 3663 13515
rect 3878 13512 3884 13524
rect 3651 13484 3884 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 3970 13472 3976 13524
rect 4028 13512 4034 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 4028 13484 4261 13512
rect 4028 13472 4034 13484
rect 4249 13481 4261 13484
rect 4295 13512 4307 13515
rect 4433 13515 4491 13521
rect 4433 13512 4445 13515
rect 4295 13484 4445 13512
rect 4295 13481 4307 13484
rect 4249 13475 4307 13481
rect 4433 13481 4445 13484
rect 4479 13481 4491 13515
rect 4890 13512 4896 13524
rect 4851 13484 4896 13512
rect 4433 13475 4491 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 6454 13512 6460 13524
rect 6415 13484 6460 13512
rect 6454 13472 6460 13484
rect 6512 13472 6518 13524
rect 7929 13515 7987 13521
rect 7929 13481 7941 13515
rect 7975 13512 7987 13515
rect 8110 13512 8116 13524
rect 7975 13484 8116 13512
rect 7975 13481 7987 13484
rect 7929 13475 7987 13481
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 8478 13512 8484 13524
rect 8439 13484 8484 13512
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 13814 13512 13820 13524
rect 13775 13484 13820 13512
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14369 13515 14427 13521
rect 14369 13512 14381 13515
rect 14240 13484 14381 13512
rect 14240 13472 14246 13484
rect 14369 13481 14381 13484
rect 14415 13481 14427 13515
rect 14369 13475 14427 13481
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 18693 13515 18751 13521
rect 18693 13512 18705 13515
rect 18380 13484 18705 13512
rect 18380 13472 18386 13484
rect 18693 13481 18705 13484
rect 18739 13481 18751 13515
rect 21082 13512 21088 13524
rect 21043 13484 21088 13512
rect 18693 13475 18751 13481
rect 21082 13472 21088 13484
rect 21140 13512 21146 13524
rect 22741 13515 22799 13521
rect 22741 13512 22753 13515
rect 21140 13484 22753 13512
rect 21140 13472 21146 13484
rect 22741 13481 22753 13484
rect 22787 13512 22799 13515
rect 23382 13512 23388 13524
rect 22787 13484 23388 13512
rect 22787 13481 22799 13484
rect 22741 13475 22799 13481
rect 23382 13472 23388 13484
rect 23440 13472 23446 13524
rect 23750 13512 23756 13524
rect 23711 13484 23756 13512
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 24026 13472 24032 13524
rect 24084 13512 24090 13524
rect 24213 13515 24271 13521
rect 24213 13512 24225 13515
rect 24084 13484 24225 13512
rect 24084 13472 24090 13484
rect 24213 13481 24225 13484
rect 24259 13481 24271 13515
rect 24213 13475 24271 13481
rect 25593 13515 25651 13521
rect 25593 13481 25605 13515
rect 25639 13512 25651 13515
rect 25774 13512 25780 13524
rect 25639 13484 25780 13512
rect 25639 13481 25651 13484
rect 25593 13475 25651 13481
rect 25774 13472 25780 13484
rect 25832 13472 25838 13524
rect 5905 13447 5963 13453
rect 5905 13413 5917 13447
rect 5951 13444 5963 13447
rect 6178 13444 6184 13456
rect 5951 13416 6184 13444
rect 5951 13413 5963 13416
rect 5905 13407 5963 13413
rect 6178 13404 6184 13416
rect 6236 13404 6242 13456
rect 6472 13444 6500 13472
rect 7377 13447 7435 13453
rect 7377 13444 7389 13447
rect 6472 13416 7389 13444
rect 7377 13413 7389 13416
rect 7423 13413 7435 13447
rect 7377 13407 7435 13413
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 9309 13447 9367 13453
rect 9309 13444 9321 13447
rect 8352 13416 9321 13444
rect 8352 13404 8358 13416
rect 9309 13413 9321 13416
rect 9355 13444 9367 13447
rect 9582 13444 9588 13456
rect 9355 13416 9588 13444
rect 9355 13413 9367 13416
rect 9309 13407 9367 13413
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 12704 13447 12762 13453
rect 12704 13413 12716 13447
rect 12750 13444 12762 13447
rect 12894 13444 12900 13456
rect 12750 13416 12900 13444
rect 12750 13413 12762 13416
rect 12704 13407 12762 13413
rect 12894 13404 12900 13416
rect 12952 13404 12958 13456
rect 16390 13404 16396 13456
rect 16448 13444 16454 13456
rect 17006 13447 17064 13453
rect 17006 13444 17018 13447
rect 16448 13416 17018 13444
rect 16448 13404 16454 13416
rect 17006 13413 17018 13416
rect 17052 13413 17064 13447
rect 17006 13407 17064 13413
rect 23290 13404 23296 13456
rect 23348 13444 23354 13456
rect 24305 13447 24363 13453
rect 24305 13444 24317 13447
rect 23348 13416 24317 13444
rect 23348 13404 23354 13416
rect 24305 13413 24317 13416
rect 24351 13444 24363 13447
rect 25038 13444 25044 13456
rect 24351 13416 25044 13444
rect 24351 13413 24363 13416
rect 24305 13407 24363 13413
rect 25038 13404 25044 13416
rect 25096 13404 25102 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2314 13376 2320 13388
rect 1443 13348 2320 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 3050 13376 3056 13388
rect 2547 13348 3056 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 4798 13376 4804 13388
rect 4759 13348 4804 13376
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 5537 13379 5595 13385
rect 5537 13345 5549 13379
rect 5583 13376 5595 13379
rect 5626 13376 5632 13388
rect 5583 13348 5632 13376
rect 5583 13345 5595 13348
rect 5537 13339 5595 13345
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 6362 13376 6368 13388
rect 6323 13348 6368 13376
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 8754 13376 8760 13388
rect 8435 13348 8760 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 9950 13376 9956 13388
rect 9911 13348 9956 13376
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10220 13379 10278 13385
rect 10220 13345 10232 13379
rect 10266 13376 10278 13379
rect 10962 13376 10968 13388
rect 10266 13348 10968 13376
rect 10266 13345 10278 13348
rect 10220 13339 10278 13345
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 12437 13379 12495 13385
rect 12437 13345 12449 13379
rect 12483 13376 12495 13379
rect 12526 13376 12532 13388
rect 12483 13348 12532 13376
rect 12483 13345 12495 13348
rect 12437 13339 12495 13345
rect 12526 13336 12532 13348
rect 12584 13336 12590 13388
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 16850 13376 16856 13388
rect 16807 13348 16856 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13376 19671 13379
rect 20622 13376 20628 13388
rect 19659 13348 20628 13376
rect 19659 13345 19671 13348
rect 19613 13339 19671 13345
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 20898 13336 20904 13388
rect 20956 13376 20962 13388
rect 21361 13379 21419 13385
rect 21361 13376 21373 13379
rect 20956 13348 21373 13376
rect 20956 13336 20962 13348
rect 21361 13345 21373 13348
rect 21407 13345 21419 13379
rect 21361 13339 21419 13345
rect 21628 13379 21686 13385
rect 21628 13345 21640 13379
rect 21674 13376 21686 13379
rect 22462 13376 22468 13388
rect 21674 13348 22468 13376
rect 21674 13345 21686 13348
rect 21628 13339 21686 13345
rect 22462 13336 22468 13348
rect 22520 13336 22526 13388
rect 25314 13336 25320 13388
rect 25372 13376 25378 13388
rect 25409 13379 25467 13385
rect 25409 13376 25421 13379
rect 25372 13348 25421 13376
rect 25372 13336 25378 13348
rect 25409 13345 25421 13348
rect 25455 13345 25467 13379
rect 25409 13339 25467 13345
rect 4246 13268 4252 13320
rect 4304 13308 4310 13320
rect 4985 13311 5043 13317
rect 4985 13308 4997 13311
rect 4304 13280 4997 13308
rect 4304 13268 4310 13280
rect 4985 13277 4997 13280
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 6086 13268 6092 13320
rect 6144 13308 6150 13320
rect 6270 13308 6276 13320
rect 6144 13280 6276 13308
rect 6144 13268 6150 13280
rect 6270 13268 6276 13280
rect 6328 13308 6334 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6328 13280 6561 13308
rect 6328 13268 6334 13280
rect 6549 13277 6561 13280
rect 6595 13308 6607 13311
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6595 13280 7021 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 7009 13277 7021 13280
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 9398 13308 9404 13320
rect 8711 13280 9404 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 2222 13200 2228 13252
rect 2280 13240 2286 13252
rect 2685 13243 2743 13249
rect 2685 13240 2697 13243
rect 2280 13212 2697 13240
rect 2280 13200 2286 13212
rect 2685 13209 2697 13212
rect 2731 13209 2743 13243
rect 8018 13240 8024 13252
rect 7979 13212 8024 13240
rect 2685 13203 2743 13209
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 8110 13200 8116 13252
rect 8168 13240 8174 13252
rect 8680 13240 8708 13271
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 15746 13308 15752 13320
rect 15707 13280 15752 13308
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 19058 13308 19064 13320
rect 19019 13280 19064 13308
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 8168 13212 8708 13240
rect 19720 13240 19748 13271
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 19852 13280 19897 13308
rect 19852 13268 19858 13280
rect 23842 13268 23848 13320
rect 23900 13308 23906 13320
rect 24118 13308 24124 13320
rect 23900 13280 24124 13308
rect 23900 13268 23906 13280
rect 24118 13268 24124 13280
rect 24176 13308 24182 13320
rect 24397 13311 24455 13317
rect 24397 13308 24409 13311
rect 24176 13280 24409 13308
rect 24176 13268 24182 13280
rect 24397 13277 24409 13280
rect 24443 13277 24455 13311
rect 24397 13271 24455 13277
rect 19720 13212 20392 13240
rect 8168 13200 8174 13212
rect 20364 13184 20392 13212
rect 3142 13172 3148 13184
rect 3103 13144 3148 13172
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 5074 13132 5080 13184
rect 5132 13172 5138 13184
rect 5997 13175 6055 13181
rect 5997 13172 6009 13175
rect 5132 13144 6009 13172
rect 5132 13132 5138 13144
rect 5997 13141 6009 13144
rect 6043 13141 6055 13175
rect 5997 13135 6055 13141
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 11422 13172 11428 13184
rect 11379 13144 11428 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 12161 13175 12219 13181
rect 12161 13172 12173 13175
rect 12124 13144 12173 13172
rect 12124 13132 12130 13144
rect 12161 13141 12173 13144
rect 12207 13141 12219 13175
rect 15470 13172 15476 13184
rect 15431 13144 15476 13172
rect 12161 13135 12219 13141
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 16298 13172 16304 13184
rect 16259 13144 16304 13172
rect 16298 13132 16304 13144
rect 16356 13132 16362 13184
rect 18141 13175 18199 13181
rect 18141 13141 18153 13175
rect 18187 13172 18199 13175
rect 18598 13172 18604 13184
rect 18187 13144 18604 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 19242 13172 19248 13184
rect 19203 13144 19248 13172
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 20346 13172 20352 13184
rect 20307 13144 20352 13172
rect 20346 13132 20352 13144
rect 20404 13132 20410 13184
rect 23382 13172 23388 13184
rect 23343 13144 23388 13172
rect 23382 13132 23388 13144
rect 23440 13132 23446 13184
rect 23842 13172 23848 13184
rect 23803 13144 23848 13172
rect 23842 13132 23848 13144
rect 23900 13132 23906 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1486 12928 1492 12980
rect 1544 12968 1550 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 1544 12940 1593 12968
rect 1544 12928 1550 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 1581 12931 1639 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3513 12971 3571 12977
rect 3513 12937 3525 12971
rect 3559 12968 3571 12971
rect 3602 12968 3608 12980
rect 3559 12940 3608 12968
rect 3559 12937 3571 12940
rect 3513 12931 3571 12937
rect 3602 12928 3608 12940
rect 3660 12928 3666 12980
rect 4246 12968 4252 12980
rect 4207 12940 4252 12968
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 4706 12968 4712 12980
rect 4667 12940 4712 12968
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 4798 12928 4804 12980
rect 4856 12968 4862 12980
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 4856 12940 5181 12968
rect 4856 12928 4862 12940
rect 5169 12937 5181 12940
rect 5215 12937 5227 12971
rect 6178 12968 6184 12980
rect 6139 12940 6184 12968
rect 5169 12931 5227 12937
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 6822 12968 6828 12980
rect 6420 12940 6828 12968
rect 6420 12928 6426 12940
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 8110 12968 8116 12980
rect 8071 12940 8116 12968
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8478 12968 8484 12980
rect 8439 12940 8484 12968
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 8754 12968 8760 12980
rect 8715 12940 8760 12968
rect 8754 12928 8760 12940
rect 8812 12968 8818 12980
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 8812 12940 9321 12968
rect 8812 12928 8818 12940
rect 9309 12937 9321 12940
rect 9355 12937 9367 12971
rect 9309 12931 9367 12937
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 10008 12940 10333 12968
rect 10008 12928 10014 12940
rect 10321 12937 10333 12940
rect 10367 12937 10379 12971
rect 10321 12931 10379 12937
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 10962 12968 10968 12980
rect 10827 12940 10968 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 13538 12968 13544 12980
rect 13499 12940 13544 12968
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 15013 12971 15071 12977
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 16301 12971 16359 12977
rect 15059 12940 15792 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 2409 12903 2467 12909
rect 2409 12869 2421 12903
rect 2455 12900 2467 12903
rect 3789 12903 3847 12909
rect 3789 12900 3801 12903
rect 2455 12872 3801 12900
rect 2455 12869 2467 12872
rect 2409 12863 2467 12869
rect 2516 12773 2544 12872
rect 3789 12869 3801 12872
rect 3835 12869 3847 12903
rect 6196 12900 6224 12928
rect 6196 12872 7420 12900
rect 3789 12863 3847 12869
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 7392 12841 7420 12872
rect 14826 12860 14832 12912
rect 14884 12900 14890 12912
rect 15105 12903 15163 12909
rect 15105 12900 15117 12903
rect 14884 12872 15117 12900
rect 14884 12860 14890 12872
rect 15105 12869 15117 12872
rect 15151 12869 15163 12903
rect 15105 12863 15163 12869
rect 6549 12835 6607 12841
rect 5776 12804 5821 12832
rect 5776 12792 5782 12804
rect 6549 12801 6561 12835
rect 6595 12832 6607 12835
rect 7377 12835 7435 12841
rect 6595 12804 7236 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 2501 12767 2559 12773
rect 1443 12736 2084 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2056 12637 2084 12736
rect 2501 12733 2513 12767
rect 2547 12733 2559 12767
rect 3602 12764 3608 12776
rect 3563 12736 3608 12764
rect 2501 12727 2559 12733
rect 3602 12724 3608 12736
rect 3660 12724 3666 12776
rect 5534 12764 5540 12776
rect 5447 12736 5540 12764
rect 5534 12724 5540 12736
rect 5592 12764 5598 12776
rect 6638 12764 6644 12776
rect 5592 12736 6644 12764
rect 5592 12724 5598 12736
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 7208 12773 7236 12804
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 9582 12792 9588 12844
rect 9640 12832 9646 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9640 12804 9873 12832
rect 9640 12792 9646 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 13722 12832 13728 12844
rect 12575 12804 13728 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 14458 12832 14464 12844
rect 14231 12804 14464 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 15764 12841 15792 12940
rect 16301 12937 16313 12971
rect 16347 12968 16359 12971
rect 16390 12968 16396 12980
rect 16347 12940 16396 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17126 12968 17132 12980
rect 17087 12940 17132 12968
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 18046 12968 18052 12980
rect 18007 12940 18052 12968
rect 18046 12928 18052 12940
rect 18104 12928 18110 12980
rect 19337 12971 19395 12977
rect 19337 12937 19349 12971
rect 19383 12968 19395 12971
rect 19426 12968 19432 12980
rect 19383 12940 19432 12968
rect 19383 12937 19395 12940
rect 19337 12931 19395 12937
rect 19426 12928 19432 12940
rect 19484 12968 19490 12980
rect 19794 12968 19800 12980
rect 19484 12940 19800 12968
rect 19484 12928 19490 12940
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 20165 12971 20223 12977
rect 20165 12937 20177 12971
rect 20211 12968 20223 12971
rect 20438 12968 20444 12980
rect 20211 12940 20444 12968
rect 20211 12937 20223 12940
rect 20165 12931 20223 12937
rect 20438 12928 20444 12940
rect 20496 12928 20502 12980
rect 20898 12928 20904 12980
rect 20956 12968 20962 12980
rect 21361 12971 21419 12977
rect 21361 12968 21373 12971
rect 20956 12940 21373 12968
rect 20956 12928 20962 12940
rect 21361 12937 21373 12940
rect 21407 12937 21419 12971
rect 21910 12968 21916 12980
rect 21871 12940 21916 12968
rect 21361 12931 21419 12937
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 23382 12968 23388 12980
rect 22388 12940 23388 12968
rect 16868 12900 16896 12928
rect 18322 12900 18328 12912
rect 16868 12872 18328 12900
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 20530 12860 20536 12912
rect 20588 12900 20594 12912
rect 20588 12872 20760 12900
rect 20588 12860 20594 12872
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12832 14703 12835
rect 15749 12835 15807 12841
rect 14691 12804 15608 12832
rect 14691 12801 14703 12804
rect 14645 12795 14703 12801
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12764 7251 12767
rect 7650 12764 7656 12776
rect 7239 12736 7656 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 9030 12764 9036 12776
rect 8956 12736 9036 12764
rect 4706 12656 4712 12708
rect 4764 12696 4770 12708
rect 5718 12696 5724 12708
rect 4764 12668 5724 12696
rect 4764 12656 4770 12668
rect 5718 12656 5724 12668
rect 5776 12656 5782 12708
rect 7282 12696 7288 12708
rect 7243 12668 7288 12696
rect 7282 12656 7288 12668
rect 7340 12696 7346 12708
rect 7926 12696 7932 12708
rect 7340 12668 7932 12696
rect 7340 12656 7346 12668
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 2041 12631 2099 12637
rect 2041 12597 2053 12631
rect 2087 12628 2099 12631
rect 2130 12628 2136 12640
rect 2087 12600 2136 12628
rect 2087 12597 2099 12600
rect 2041 12591 2099 12597
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 2682 12628 2688 12640
rect 2643 12600 2688 12628
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 3418 12588 3424 12640
rect 3476 12628 3482 12640
rect 4982 12628 4988 12640
rect 3476 12600 4988 12628
rect 3476 12588 3482 12600
rect 4982 12588 4988 12600
rect 5040 12628 5046 12640
rect 5629 12631 5687 12637
rect 5629 12628 5641 12631
rect 5040 12600 5641 12628
rect 5040 12588 5046 12600
rect 5629 12597 5641 12600
rect 5675 12597 5687 12631
rect 5629 12591 5687 12597
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 8956 12628 8984 12736
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 9769 12767 9827 12773
rect 9769 12764 9781 12767
rect 9732 12736 9781 12764
rect 9732 12724 9738 12736
rect 9769 12733 9781 12736
rect 9815 12764 9827 12767
rect 10042 12764 10048 12776
rect 9815 12736 10048 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 13446 12764 13452 12776
rect 13359 12736 13452 12764
rect 13446 12724 13452 12736
rect 13504 12764 13510 12776
rect 13998 12764 14004 12776
rect 13504 12736 14004 12764
rect 13504 12724 13510 12736
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 15470 12764 15476 12776
rect 15431 12736 15476 12764
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 15580 12773 15608 12804
rect 15749 12801 15761 12835
rect 15795 12832 15807 12835
rect 16482 12832 16488 12844
rect 15795 12804 16488 12832
rect 15795 12801 15807 12804
rect 15749 12795 15807 12801
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 18414 12832 18420 12844
rect 17543 12804 18420 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 18414 12792 18420 12804
rect 18472 12832 18478 12844
rect 20732 12841 20760 12872
rect 22388 12841 22416 12940
rect 23382 12928 23388 12940
rect 23440 12968 23446 12980
rect 23661 12971 23719 12977
rect 23661 12968 23673 12971
rect 23440 12940 23673 12968
rect 23440 12928 23446 12940
rect 23661 12937 23673 12940
rect 23707 12937 23719 12971
rect 23661 12931 23719 12937
rect 24118 12928 24124 12980
rect 24176 12968 24182 12980
rect 24673 12971 24731 12977
rect 24673 12968 24685 12971
rect 24176 12940 24685 12968
rect 24176 12928 24182 12940
rect 24673 12937 24685 12940
rect 24719 12937 24731 12971
rect 25038 12968 25044 12980
rect 24999 12940 25044 12968
rect 24673 12931 24731 12937
rect 25038 12928 25044 12940
rect 25096 12928 25102 12980
rect 23474 12900 23480 12912
rect 23435 12872 23480 12900
rect 23474 12860 23480 12872
rect 23532 12860 23538 12912
rect 24026 12860 24032 12912
rect 24084 12900 24090 12912
rect 24394 12900 24400 12912
rect 24084 12872 24400 12900
rect 24084 12860 24090 12872
rect 24394 12860 24400 12872
rect 24452 12860 24458 12912
rect 25314 12860 25320 12912
rect 25372 12900 25378 12912
rect 26145 12903 26203 12909
rect 26145 12900 26157 12903
rect 25372 12872 26157 12900
rect 25372 12860 25378 12872
rect 26145 12869 26157 12872
rect 26191 12869 26203 12903
rect 26145 12863 26203 12869
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 18472 12804 18613 12832
rect 18472 12792 18478 12804
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12801 20775 12835
rect 20717 12795 20775 12801
rect 22373 12835 22431 12841
rect 22373 12801 22385 12835
rect 22419 12801 22431 12835
rect 22554 12832 22560 12844
rect 22515 12804 22560 12832
rect 22373 12795 22431 12801
rect 22554 12792 22560 12804
rect 22612 12792 22618 12844
rect 23106 12832 23112 12844
rect 23019 12804 23112 12832
rect 23106 12792 23112 12804
rect 23164 12832 23170 12844
rect 24213 12835 24271 12841
rect 24213 12832 24225 12835
rect 23164 12804 24225 12832
rect 23164 12792 23170 12804
rect 24213 12801 24225 12804
rect 24259 12801 24271 12835
rect 24213 12795 24271 12801
rect 24302 12792 24308 12844
rect 24360 12832 24366 12844
rect 24670 12832 24676 12844
rect 24360 12804 24676 12832
rect 24360 12792 24366 12804
rect 24670 12792 24676 12804
rect 24728 12792 24734 12844
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12764 15623 12767
rect 15930 12764 15936 12776
rect 15611 12736 15936 12764
rect 15611 12733 15623 12736
rect 15565 12727 15623 12733
rect 15930 12724 15936 12736
rect 15988 12724 15994 12776
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 16301 12767 16359 12773
rect 16301 12764 16313 12767
rect 16264 12736 16313 12764
rect 16264 12724 16270 12736
rect 16301 12733 16313 12736
rect 16347 12733 16359 12767
rect 16942 12764 16948 12776
rect 16903 12736 16948 12764
rect 16301 12727 16359 12733
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 17865 12767 17923 12773
rect 17865 12733 17877 12767
rect 17911 12764 17923 12767
rect 18230 12764 18236 12776
rect 17911 12736 18236 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18230 12724 18236 12736
rect 18288 12764 18294 12776
rect 18509 12767 18567 12773
rect 18509 12764 18521 12767
rect 18288 12736 18521 12764
rect 18288 12724 18294 12736
rect 18509 12733 18521 12736
rect 18555 12764 18567 12767
rect 19150 12764 19156 12776
rect 18555 12736 19156 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 19392 12736 19717 12764
rect 19392 12724 19398 12736
rect 19705 12733 19717 12736
rect 19751 12764 19763 12767
rect 20625 12767 20683 12773
rect 20625 12764 20637 12767
rect 19751 12736 20637 12764
rect 19751 12733 19763 12736
rect 19705 12727 19763 12733
rect 20625 12733 20637 12736
rect 20671 12764 20683 12767
rect 22186 12764 22192 12776
rect 20671 12736 22192 12764
rect 20671 12733 20683 12736
rect 20625 12727 20683 12733
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 23474 12724 23480 12776
rect 23532 12764 23538 12776
rect 24029 12767 24087 12773
rect 24029 12764 24041 12767
rect 23532 12736 24041 12764
rect 23532 12724 23538 12736
rect 24029 12733 24041 12736
rect 24075 12733 24087 12767
rect 24029 12727 24087 12733
rect 25038 12724 25044 12776
rect 25096 12764 25102 12776
rect 25225 12767 25283 12773
rect 25225 12764 25237 12767
rect 25096 12736 25237 12764
rect 25096 12724 25102 12736
rect 25225 12733 25237 12736
rect 25271 12764 25283 12767
rect 25777 12767 25835 12773
rect 25777 12764 25789 12767
rect 25271 12736 25789 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 25777 12733 25789 12736
rect 25823 12733 25835 12767
rect 25777 12727 25835 12733
rect 9490 12656 9496 12708
rect 9548 12696 9554 12708
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 9548 12668 10977 12696
rect 9548 12656 9554 12668
rect 10965 12665 10977 12668
rect 11011 12665 11023 12699
rect 10965 12659 11023 12665
rect 11606 12656 11612 12708
rect 11664 12696 11670 12708
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 11664 12668 12173 12696
rect 11664 12656 11670 12668
rect 12161 12665 12173 12668
rect 12207 12665 12219 12699
rect 12161 12659 12219 12665
rect 13538 12656 13544 12708
rect 13596 12696 13602 12708
rect 13909 12699 13967 12705
rect 13909 12696 13921 12699
rect 13596 12668 13921 12696
rect 13596 12656 13602 12668
rect 13909 12665 13921 12668
rect 13955 12696 13967 12699
rect 14182 12696 14188 12708
rect 13955 12668 14188 12696
rect 13955 12665 13967 12668
rect 13909 12659 13967 12665
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 15654 12656 15660 12708
rect 15712 12696 15718 12708
rect 16114 12696 16120 12708
rect 15712 12668 16120 12696
rect 15712 12656 15718 12668
rect 16114 12656 16120 12668
rect 16172 12656 16178 12708
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 20073 12699 20131 12705
rect 20073 12696 20085 12699
rect 19576 12668 20085 12696
rect 19576 12656 19582 12668
rect 20073 12665 20085 12668
rect 20119 12696 20131 12699
rect 20438 12696 20444 12708
rect 20119 12668 20444 12696
rect 20119 12665 20131 12668
rect 20073 12659 20131 12665
rect 20438 12656 20444 12668
rect 20496 12696 20502 12708
rect 20533 12699 20591 12705
rect 20533 12696 20545 12699
rect 20496 12668 20545 12696
rect 20496 12656 20502 12668
rect 20533 12665 20545 12668
rect 20579 12665 20591 12699
rect 20533 12659 20591 12665
rect 21542 12656 21548 12708
rect 21600 12696 21606 12708
rect 22462 12696 22468 12708
rect 21600 12668 22468 12696
rect 21600 12656 21606 12668
rect 22462 12656 22468 12668
rect 22520 12656 22526 12708
rect 23934 12656 23940 12708
rect 23992 12696 23998 12708
rect 24302 12696 24308 12708
rect 23992 12668 24308 12696
rect 23992 12656 23998 12668
rect 24302 12656 24308 12668
rect 24360 12656 24366 12708
rect 8904 12600 8984 12628
rect 8904 12588 8910 12600
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 9125 12631 9183 12637
rect 9125 12628 9137 12631
rect 9088 12600 9137 12628
rect 9088 12588 9094 12600
rect 9125 12597 9137 12600
rect 9171 12628 9183 12631
rect 9677 12631 9735 12637
rect 9677 12628 9689 12631
rect 9171 12600 9689 12628
rect 9171 12597 9183 12600
rect 9125 12591 9183 12597
rect 9677 12597 9689 12600
rect 9723 12628 9735 12631
rect 9766 12628 9772 12640
rect 9723 12600 9772 12628
rect 9723 12597 9735 12600
rect 9677 12591 9735 12597
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 12618 12588 12624 12640
rect 12676 12628 12682 12640
rect 12989 12631 13047 12637
rect 12989 12628 13001 12631
rect 12676 12600 13001 12628
rect 12676 12588 12682 12600
rect 12989 12597 13001 12600
rect 13035 12597 13047 12631
rect 12989 12591 13047 12597
rect 15562 12588 15568 12640
rect 15620 12628 15626 12640
rect 15930 12628 15936 12640
rect 15620 12600 15936 12628
rect 15620 12588 15626 12600
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 18138 12588 18144 12640
rect 18196 12628 18202 12640
rect 18417 12631 18475 12637
rect 18417 12628 18429 12631
rect 18196 12600 18429 12628
rect 18196 12588 18202 12600
rect 18417 12597 18429 12600
rect 18463 12597 18475 12631
rect 18417 12591 18475 12597
rect 21821 12631 21879 12637
rect 21821 12597 21833 12631
rect 21867 12628 21879 12631
rect 22281 12631 22339 12637
rect 22281 12628 22293 12631
rect 21867 12600 22293 12628
rect 21867 12597 21879 12600
rect 21821 12591 21879 12597
rect 22281 12597 22293 12600
rect 22327 12628 22339 12631
rect 22922 12628 22928 12640
rect 22327 12600 22928 12628
rect 22327 12597 22339 12600
rect 22281 12591 22339 12597
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 23750 12588 23756 12640
rect 23808 12628 23814 12640
rect 24121 12631 24179 12637
rect 24121 12628 24133 12631
rect 23808 12600 24133 12628
rect 23808 12588 23814 12600
rect 24121 12597 24133 12600
rect 24167 12628 24179 12631
rect 24578 12628 24584 12640
rect 24167 12600 24584 12628
rect 24167 12597 24179 12600
rect 24121 12591 24179 12597
rect 24578 12588 24584 12600
rect 24636 12588 24642 12640
rect 25406 12628 25412 12640
rect 25367 12600 25412 12628
rect 25406 12588 25412 12600
rect 25464 12588 25470 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 2038 12424 2044 12436
rect 1999 12396 2044 12424
rect 2038 12384 2044 12396
rect 2096 12384 2102 12436
rect 2314 12424 2320 12436
rect 2275 12396 2320 12424
rect 2314 12384 2320 12396
rect 2372 12424 2378 12436
rect 2685 12427 2743 12433
rect 2685 12424 2697 12427
rect 2372 12396 2697 12424
rect 2372 12384 2378 12396
rect 2685 12393 2697 12396
rect 2731 12393 2743 12427
rect 2685 12387 2743 12393
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 2961 12427 3019 12433
rect 2961 12424 2973 12427
rect 2832 12396 2973 12424
rect 2832 12384 2838 12396
rect 2961 12393 2973 12396
rect 3007 12393 3019 12427
rect 2961 12387 3019 12393
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 4614 12424 4620 12436
rect 3927 12396 4620 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 4798 12424 4804 12436
rect 4759 12396 4804 12424
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 5626 12424 5632 12436
rect 5587 12396 5632 12424
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 6917 12427 6975 12433
rect 6917 12393 6929 12427
rect 6963 12424 6975 12427
rect 7006 12424 7012 12436
rect 6963 12396 7012 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8352 12396 8953 12424
rect 8352 12384 8358 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 8941 12387 8999 12393
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 9582 12424 9588 12436
rect 9447 12396 9588 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 4525 12359 4583 12365
rect 4525 12325 4537 12359
rect 4571 12356 4583 12359
rect 4890 12356 4896 12368
rect 4571 12328 4896 12356
rect 4571 12325 4583 12328
rect 4525 12319 4583 12325
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 7374 12316 7380 12368
rect 7432 12356 7438 12368
rect 7653 12359 7711 12365
rect 7653 12356 7665 12359
rect 7432 12328 7665 12356
rect 7432 12316 7438 12328
rect 7653 12325 7665 12328
rect 7699 12325 7711 12359
rect 8956 12356 8984 12387
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 12894 12424 12900 12436
rect 11664 12396 12900 12424
rect 11664 12384 11670 12396
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13538 12424 13544 12436
rect 13499 12396 13544 12424
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 20349 12427 20407 12433
rect 20349 12393 20361 12427
rect 20395 12424 20407 12427
rect 20530 12424 20536 12436
rect 20395 12396 20536 12424
rect 20395 12393 20407 12396
rect 20349 12387 20407 12393
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 21177 12427 21235 12433
rect 21177 12393 21189 12427
rect 21223 12424 21235 12427
rect 21223 12396 21956 12424
rect 21223 12393 21235 12396
rect 21177 12387 21235 12393
rect 10137 12359 10195 12365
rect 10137 12356 10149 12359
rect 8956 12328 10149 12356
rect 7653 12319 7711 12325
rect 10137 12325 10149 12328
rect 10183 12325 10195 12359
rect 21634 12356 21640 12368
rect 10137 12319 10195 12325
rect 21284 12328 21640 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1578 12288 1584 12300
rect 1443 12260 1584 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12288 2559 12291
rect 2590 12288 2596 12300
rect 2547 12260 2596 12288
rect 2547 12257 2559 12260
rect 2501 12251 2559 12257
rect 2590 12248 2596 12260
rect 2648 12288 2654 12300
rect 2958 12288 2964 12300
rect 2648 12260 2964 12288
rect 2648 12248 2654 12260
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 5442 12288 5448 12300
rect 5307 12260 5448 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 5994 12288 6000 12300
rect 5955 12260 6000 12288
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12288 6147 12291
rect 6270 12288 6276 12300
rect 6135 12260 6276 12288
rect 6135 12257 6147 12260
rect 6089 12251 6147 12257
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7561 12291 7619 12297
rect 7561 12288 7573 12291
rect 7248 12260 7573 12288
rect 7248 12248 7254 12260
rect 7561 12257 7573 12260
rect 7607 12288 7619 12291
rect 7834 12288 7840 12300
rect 7607 12260 7840 12288
rect 7607 12257 7619 12260
rect 7561 12251 7619 12257
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 11422 12248 11428 12300
rect 11480 12288 11486 12300
rect 11784 12291 11842 12297
rect 11784 12288 11796 12291
rect 11480 12260 11796 12288
rect 11480 12248 11486 12260
rect 11784 12257 11796 12260
rect 11830 12288 11842 12291
rect 12158 12288 12164 12300
rect 11830 12260 12164 12288
rect 11830 12257 11842 12260
rect 11784 12251 11842 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12288 15347 12291
rect 15378 12288 15384 12300
rect 15335 12260 15384 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 15562 12297 15568 12300
rect 15556 12288 15568 12297
rect 15475 12260 15568 12288
rect 15556 12251 15568 12260
rect 15620 12288 15626 12300
rect 16850 12288 16856 12300
rect 15620 12260 16856 12288
rect 15562 12248 15568 12251
rect 15620 12248 15626 12260
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 18598 12297 18604 12300
rect 18592 12288 18604 12297
rect 18559 12260 18604 12288
rect 18592 12251 18604 12260
rect 18598 12248 18604 12251
rect 18656 12248 18662 12300
rect 20438 12248 20444 12300
rect 20496 12288 20502 12300
rect 21284 12297 21312 12328
rect 21634 12316 21640 12328
rect 21692 12316 21698 12368
rect 21928 12365 21956 12396
rect 24394 12384 24400 12436
rect 24452 12424 24458 12436
rect 24673 12427 24731 12433
rect 24673 12424 24685 12427
rect 24452 12396 24685 12424
rect 24452 12384 24458 12396
rect 24673 12393 24685 12396
rect 24719 12393 24731 12427
rect 24673 12387 24731 12393
rect 24857 12427 24915 12433
rect 24857 12393 24869 12427
rect 24903 12424 24915 12427
rect 24946 12424 24952 12436
rect 24903 12396 24952 12424
rect 24903 12393 24915 12396
rect 24857 12387 24915 12393
rect 24946 12384 24952 12396
rect 25004 12384 25010 12436
rect 25225 12427 25283 12433
rect 25225 12393 25237 12427
rect 25271 12424 25283 12427
rect 25590 12424 25596 12436
rect 25271 12396 25596 12424
rect 25271 12393 25283 12396
rect 25225 12387 25283 12393
rect 25590 12384 25596 12396
rect 25648 12384 25654 12436
rect 21913 12359 21971 12365
rect 21913 12325 21925 12359
rect 21959 12356 21971 12359
rect 22554 12356 22560 12368
rect 21959 12328 22560 12356
rect 21959 12325 21971 12328
rect 21913 12319 21971 12325
rect 22554 12316 22560 12328
rect 22612 12356 22618 12368
rect 22612 12328 23244 12356
rect 22612 12316 22618 12328
rect 21269 12291 21327 12297
rect 21269 12288 21281 12291
rect 20496 12260 21281 12288
rect 20496 12248 20502 12260
rect 21269 12257 21281 12260
rect 21315 12257 21327 12291
rect 21269 12251 21327 12257
rect 22281 12291 22339 12297
rect 22281 12257 22293 12291
rect 22327 12288 22339 12291
rect 22640 12291 22698 12297
rect 22640 12288 22652 12291
rect 22327 12260 22652 12288
rect 22327 12257 22339 12260
rect 22281 12251 22339 12257
rect 22640 12257 22652 12260
rect 22686 12288 22698 12291
rect 23106 12288 23112 12300
rect 22686 12260 23112 12288
rect 22686 12257 22698 12260
rect 22640 12251 22698 12257
rect 23106 12248 23112 12260
rect 23164 12248 23170 12300
rect 23216 12288 23244 12328
rect 24578 12316 24584 12368
rect 24636 12356 24642 12368
rect 25317 12359 25375 12365
rect 25317 12356 25329 12359
rect 24636 12328 25329 12356
rect 24636 12316 24642 12328
rect 23216 12260 23796 12288
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6454 12220 6460 12232
rect 6227 12192 6460 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 7742 12220 7748 12232
rect 7703 12192 7748 12220
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 10192 12192 10241 12220
rect 10192 12180 10198 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 11514 12220 11520 12232
rect 11475 12192 11520 12220
rect 10229 12183 10287 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 14182 12220 14188 12232
rect 14143 12192 14188 12220
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 18322 12220 18328 12232
rect 18283 12192 18328 12220
rect 18322 12180 18328 12192
rect 18380 12180 18386 12232
rect 20714 12220 20720 12232
rect 20675 12192 20720 12220
rect 20714 12180 20720 12192
rect 20772 12180 20778 12232
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22373 12223 22431 12229
rect 22373 12220 22385 12223
rect 22244 12192 22385 12220
rect 22244 12180 22250 12192
rect 22373 12189 22385 12192
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7193 12155 7251 12161
rect 7193 12152 7205 12155
rect 6972 12124 7205 12152
rect 6972 12112 6978 12124
rect 7193 12121 7205 12124
rect 7239 12121 7251 12155
rect 7193 12115 7251 12121
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 8665 12155 8723 12161
rect 8665 12152 8677 12155
rect 8628 12124 8677 12152
rect 8628 12112 8634 12124
rect 8665 12121 8677 12124
rect 8711 12152 8723 12155
rect 9677 12155 9735 12161
rect 9677 12152 9689 12155
rect 8711 12124 9689 12152
rect 8711 12121 8723 12124
rect 8665 12115 8723 12121
rect 9677 12121 9689 12124
rect 9723 12121 9735 12155
rect 9677 12115 9735 12121
rect 10873 12155 10931 12161
rect 10873 12121 10885 12155
rect 10919 12152 10931 12155
rect 11422 12152 11428 12164
rect 10919 12124 11428 12152
rect 10919 12121 10931 12124
rect 10873 12115 10931 12121
rect 11422 12112 11428 12124
rect 11480 12112 11486 12164
rect 21453 12155 21511 12161
rect 21453 12121 21465 12155
rect 21499 12152 21511 12155
rect 22002 12152 22008 12164
rect 21499 12124 22008 12152
rect 21499 12121 21511 12124
rect 21453 12115 21511 12121
rect 22002 12112 22008 12124
rect 22060 12112 22066 12164
rect 23768 12161 23796 12260
rect 25056 12232 25084 12328
rect 25317 12325 25329 12328
rect 25363 12325 25375 12359
rect 25317 12319 25375 12325
rect 25038 12180 25044 12232
rect 25096 12180 25102 12232
rect 25409 12223 25467 12229
rect 25409 12189 25421 12223
rect 25455 12189 25467 12223
rect 25409 12183 25467 12189
rect 23753 12155 23811 12161
rect 23753 12121 23765 12155
rect 23799 12121 23811 12155
rect 24302 12152 24308 12164
rect 24263 12124 24308 12152
rect 23753 12115 23811 12121
rect 24302 12112 24308 12124
rect 24360 12152 24366 12164
rect 25424 12152 25452 12183
rect 26142 12152 26148 12164
rect 24360 12124 26148 12152
rect 24360 12112 24366 12124
rect 26142 12112 26148 12124
rect 26200 12112 26206 12164
rect 8294 12084 8300 12096
rect 8255 12056 8300 12084
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 11238 12084 11244 12096
rect 11199 12056 11244 12084
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 11514 12044 11520 12096
rect 11572 12084 11578 12096
rect 12618 12084 12624 12096
rect 11572 12056 12624 12084
rect 11572 12044 11578 12056
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 14001 12087 14059 12093
rect 14001 12053 14013 12087
rect 14047 12084 14059 12087
rect 14458 12084 14464 12096
rect 14047 12056 14464 12084
rect 14047 12053 14059 12056
rect 14001 12047 14059 12053
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 16206 12084 16212 12096
rect 15151 12056 16212 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 16666 12084 16672 12096
rect 16627 12056 16672 12084
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17313 12087 17371 12093
rect 17313 12084 17325 12087
rect 17000 12056 17325 12084
rect 17000 12044 17006 12056
rect 17313 12053 17325 12056
rect 17359 12084 17371 12087
rect 17862 12084 17868 12096
rect 17359 12056 17868 12084
rect 17359 12053 17371 12056
rect 17313 12047 17371 12053
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 18138 12084 18144 12096
rect 18099 12056 18144 12084
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 19705 12087 19763 12093
rect 19705 12084 19717 12087
rect 19484 12056 19717 12084
rect 19484 12044 19490 12056
rect 19705 12053 19717 12056
rect 19751 12053 19763 12087
rect 19705 12047 19763 12053
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 20438 12084 20444 12096
rect 20220 12056 20444 12084
rect 20220 12044 20226 12056
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 24210 12044 24216 12096
rect 24268 12084 24274 12096
rect 24320 12084 24348 12112
rect 24268 12056 24348 12084
rect 24268 12044 24274 12056
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11880 1642 11892
rect 1857 11883 1915 11889
rect 1857 11880 1869 11883
rect 1636 11852 1869 11880
rect 1636 11840 1642 11852
rect 1857 11849 1869 11852
rect 1903 11849 1915 11883
rect 2590 11880 2596 11892
rect 2551 11852 2596 11880
rect 1857 11843 1915 11849
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 4985 11883 5043 11889
rect 4985 11849 4997 11883
rect 5031 11880 5043 11883
rect 5258 11880 5264 11892
rect 5031 11852 5264 11880
rect 5031 11849 5043 11852
rect 4985 11843 5043 11849
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 6086 11880 6092 11892
rect 6047 11852 6092 11880
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 7190 11880 7196 11892
rect 7151 11852 7196 11880
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7558 11880 7564 11892
rect 7519 11852 7564 11880
rect 7558 11840 7564 11852
rect 7616 11880 7622 11892
rect 7616 11852 8156 11880
rect 7616 11840 7622 11852
rect 4617 11815 4675 11821
rect 4617 11781 4629 11815
rect 4663 11812 4675 11815
rect 5074 11812 5080 11824
rect 4663 11784 5080 11812
rect 4663 11781 4675 11784
rect 4617 11775 4675 11781
rect 5074 11772 5080 11784
rect 5132 11772 5138 11824
rect 6270 11772 6276 11824
rect 6328 11812 6334 11824
rect 7653 11815 7711 11821
rect 7653 11812 7665 11815
rect 6328 11784 7665 11812
rect 6328 11772 6334 11784
rect 7653 11781 7665 11784
rect 7699 11781 7711 11815
rect 7653 11775 7711 11781
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 6288 11744 6316 11772
rect 5307 11716 6316 11744
rect 6641 11747 6699 11753
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 7742 11744 7748 11756
rect 6687 11716 7748 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 8128 11753 8156 11852
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 9180 11852 9229 11880
rect 9180 11840 9186 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9217 11843 9275 11849
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 10100 11852 10241 11880
rect 10100 11840 10106 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 10778 11880 10784 11892
rect 10739 11852 10784 11880
rect 10229 11843 10287 11849
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11572 11852 11805 11880
rect 11572 11840 11578 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15749 11883 15807 11889
rect 15749 11880 15761 11883
rect 15528 11852 15761 11880
rect 15528 11840 15534 11852
rect 15749 11849 15761 11852
rect 15795 11849 15807 11883
rect 15749 11843 15807 11849
rect 21634 11840 21640 11892
rect 21692 11880 21698 11892
rect 21821 11883 21879 11889
rect 21821 11880 21833 11883
rect 21692 11852 21833 11880
rect 21692 11840 21698 11852
rect 21821 11849 21833 11852
rect 21867 11849 21879 11883
rect 21821 11843 21879 11849
rect 22649 11883 22707 11889
rect 22649 11849 22661 11883
rect 22695 11880 22707 11883
rect 22830 11880 22836 11892
rect 22695 11852 22836 11880
rect 22695 11849 22707 11852
rect 22649 11843 22707 11849
rect 22830 11840 22836 11852
rect 22888 11840 22894 11892
rect 23014 11880 23020 11892
rect 22975 11852 23020 11880
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 23658 11880 23664 11892
rect 23619 11852 23664 11880
rect 23658 11840 23664 11852
rect 23716 11840 23722 11892
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25409 11883 25467 11889
rect 25409 11880 25421 11883
rect 24912 11852 25421 11880
rect 24912 11840 24918 11852
rect 25409 11849 25421 11852
rect 25455 11849 25467 11883
rect 26142 11880 26148 11892
rect 26103 11852 26148 11880
rect 25409 11843 25467 11849
rect 26142 11840 26148 11852
rect 26200 11840 26206 11892
rect 9306 11772 9312 11824
rect 9364 11812 9370 11824
rect 9364 11784 9812 11812
rect 9364 11772 9370 11784
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11744 9183 11747
rect 9398 11744 9404 11756
rect 9171 11716 9404 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11676 1458 11688
rect 2225 11679 2283 11685
rect 2225 11676 2237 11679
rect 1452 11648 2237 11676
rect 1452 11636 1458 11648
rect 2225 11645 2237 11648
rect 2271 11645 2283 11679
rect 2225 11639 2283 11645
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 6454 11676 6460 11688
rect 5767 11648 6460 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 8021 11679 8079 11685
rect 8021 11676 8033 11679
rect 7156 11648 8033 11676
rect 7156 11636 7162 11648
rect 8021 11645 8033 11648
rect 8067 11645 8079 11679
rect 8312 11676 8340 11707
rect 9398 11704 9404 11716
rect 9456 11744 9462 11756
rect 9784 11753 9812 11784
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 14645 11815 14703 11821
rect 14645 11812 14657 11815
rect 14516 11784 14657 11812
rect 14516 11772 14522 11784
rect 14645 11781 14657 11784
rect 14691 11812 14703 11815
rect 15562 11812 15568 11824
rect 14691 11784 15568 11812
rect 14691 11781 14703 11784
rect 14645 11775 14703 11781
rect 15562 11772 15568 11784
rect 15620 11772 15626 11824
rect 16022 11772 16028 11824
rect 16080 11812 16086 11824
rect 24949 11815 25007 11821
rect 16080 11784 16436 11812
rect 16080 11772 16086 11784
rect 9769 11747 9827 11753
rect 9456 11716 9628 11744
rect 9456 11704 9462 11716
rect 8570 11676 8576 11688
rect 8312 11648 8576 11676
rect 8021 11639 8079 11645
rect 8570 11636 8576 11648
rect 8628 11676 8634 11688
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8628 11648 8769 11676
rect 8628 11636 8634 11648
rect 8757 11645 8769 11648
rect 8803 11676 8815 11679
rect 9214 11676 9220 11688
rect 8803 11648 9220 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 9214 11636 9220 11648
rect 9272 11636 9278 11688
rect 9600 11685 9628 11716
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 11238 11744 11244 11756
rect 11199 11716 11244 11744
rect 9769 11707 9827 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11422 11744 11428 11756
rect 11383 11716 11428 11744
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 16206 11744 16212 11756
rect 16167 11716 16212 11744
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 16408 11753 16436 11784
rect 24949 11781 24961 11815
rect 24995 11812 25007 11815
rect 25038 11812 25044 11824
rect 24995 11784 25044 11812
rect 24995 11781 25007 11784
rect 24949 11775 25007 11781
rect 25038 11772 25044 11784
rect 25096 11772 25102 11824
rect 16393 11747 16451 11753
rect 16393 11713 16405 11747
rect 16439 11744 16451 11747
rect 16666 11744 16672 11756
rect 16439 11716 16672 11744
rect 16439 11713 16451 11716
rect 16393 11707 16451 11713
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 17497 11747 17555 11753
rect 17497 11744 17509 11747
rect 16908 11716 17509 11744
rect 16908 11704 16914 11716
rect 17497 11713 17509 11716
rect 17543 11744 17555 11747
rect 18414 11744 18420 11756
rect 17543 11716 18420 11744
rect 17543 11713 17555 11716
rect 17497 11707 17555 11713
rect 18414 11704 18420 11716
rect 18472 11744 18478 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 18472 11716 18613 11744
rect 18472 11704 18478 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 24210 11744 24216 11756
rect 24171 11716 24216 11744
rect 18601 11707 18659 11713
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11676 10747 11679
rect 11146 11676 11152 11688
rect 10735 11648 11152 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 13081 11679 13139 11685
rect 13081 11676 13093 11679
rect 12676 11648 13093 11676
rect 12676 11636 12682 11648
rect 13081 11645 13093 11648
rect 13127 11676 13139 11679
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 13127 11648 13277 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 13265 11645 13277 11648
rect 13311 11676 13323 11679
rect 17681 11679 17739 11685
rect 13311 11648 15332 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 8294 11568 8300 11620
rect 8352 11608 8358 11620
rect 9674 11608 9680 11620
rect 8352 11580 9680 11608
rect 8352 11568 8358 11580
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 12158 11608 12164 11620
rect 12119 11580 12164 11608
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 12805 11611 12863 11617
rect 12805 11577 12817 11611
rect 12851 11608 12863 11611
rect 13170 11608 13176 11620
rect 12851 11580 13176 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 13170 11568 13176 11580
rect 13228 11608 13234 11620
rect 13510 11611 13568 11617
rect 13510 11608 13522 11611
rect 13228 11580 13522 11608
rect 13228 11568 13234 11580
rect 13510 11577 13522 11580
rect 13556 11577 13568 11611
rect 13510 11571 13568 11577
rect 15304 11552 15332 11648
rect 17681 11645 17693 11679
rect 17727 11676 17739 11679
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 17727 11648 18521 11676
rect 17727 11645 17739 11648
rect 17681 11639 17739 11645
rect 18509 11645 18521 11648
rect 18555 11676 18567 11679
rect 19518 11676 19524 11688
rect 18555 11648 19524 11676
rect 18555 11645 18567 11648
rect 18509 11639 18567 11645
rect 19518 11636 19524 11648
rect 19576 11636 19582 11688
rect 19889 11679 19947 11685
rect 19889 11645 19901 11679
rect 19935 11676 19947 11679
rect 20714 11676 20720 11688
rect 19935 11648 20720 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 16117 11611 16175 11617
rect 16117 11577 16129 11611
rect 16163 11608 16175 11611
rect 16163 11580 18092 11608
rect 16163 11577 16175 11580
rect 16117 11571 16175 11577
rect 18064 11552 18092 11580
rect 18322 11568 18328 11620
rect 18380 11608 18386 11620
rect 19061 11611 19119 11617
rect 19061 11608 19073 11611
rect 18380 11580 19073 11608
rect 18380 11568 18386 11580
rect 19061 11577 19073 11580
rect 19107 11608 19119 11611
rect 19705 11611 19763 11617
rect 19705 11608 19717 11611
rect 19107 11580 19717 11608
rect 19107 11577 19119 11580
rect 19061 11571 19119 11577
rect 19705 11577 19717 11580
rect 19751 11608 19763 11611
rect 19904 11608 19932 11639
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 22278 11636 22284 11688
rect 22336 11676 22342 11688
rect 22465 11679 22523 11685
rect 22465 11676 22477 11679
rect 22336 11648 22477 11676
rect 22336 11636 22342 11648
rect 22465 11645 22477 11648
rect 22511 11676 22523 11679
rect 23014 11676 23020 11688
rect 22511 11648 23020 11676
rect 22511 11645 22523 11648
rect 22465 11639 22523 11645
rect 23014 11636 23020 11648
rect 23072 11636 23078 11688
rect 24026 11676 24032 11688
rect 23987 11648 24032 11676
rect 24026 11636 24032 11648
rect 24084 11636 24090 11688
rect 25225 11679 25283 11685
rect 25225 11645 25237 11679
rect 25271 11676 25283 11679
rect 25682 11676 25688 11688
rect 25271 11648 25688 11676
rect 25271 11645 25283 11648
rect 25225 11639 25283 11645
rect 25682 11636 25688 11648
rect 25740 11676 25746 11688
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 25740 11648 25789 11676
rect 25740 11636 25746 11648
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 20162 11617 20168 11620
rect 20156 11608 20168 11617
rect 19751 11580 19932 11608
rect 20123 11580 20168 11608
rect 19751 11577 19763 11580
rect 19705 11571 19763 11577
rect 20156 11571 20168 11580
rect 20162 11568 20168 11571
rect 20220 11568 20226 11620
rect 24121 11611 24179 11617
rect 24121 11608 24133 11611
rect 23492 11580 24133 11608
rect 23492 11552 23520 11580
rect 24121 11577 24133 11580
rect 24167 11577 24179 11611
rect 24121 11571 24179 11577
rect 15286 11540 15292 11552
rect 15247 11512 15292 11540
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 17681 11543 17739 11549
rect 17681 11540 17693 11543
rect 17460 11512 17693 11540
rect 17460 11500 17466 11512
rect 17681 11509 17693 11512
rect 17727 11540 17739 11543
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 17727 11512 17785 11540
rect 17727 11509 17739 11512
rect 17681 11503 17739 11509
rect 17773 11509 17785 11512
rect 17819 11509 17831 11543
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 17773 11503 17831 11509
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18138 11500 18144 11552
rect 18196 11540 18202 11552
rect 18417 11543 18475 11549
rect 18417 11540 18429 11543
rect 18196 11512 18429 11540
rect 18196 11500 18202 11512
rect 18417 11509 18429 11512
rect 18463 11509 18475 11543
rect 18417 11503 18475 11509
rect 21269 11543 21327 11549
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 21450 11540 21456 11552
rect 21315 11512 21456 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21450 11500 21456 11512
rect 21508 11500 21514 11552
rect 22186 11500 22192 11552
rect 22244 11540 22250 11552
rect 22373 11543 22431 11549
rect 22373 11540 22385 11543
rect 22244 11512 22385 11540
rect 22244 11500 22250 11512
rect 22373 11509 22385 11512
rect 22419 11540 22431 11543
rect 22462 11540 22468 11552
rect 22419 11512 22468 11540
rect 22419 11509 22431 11512
rect 22373 11503 22431 11509
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 23474 11540 23480 11552
rect 23435 11512 23480 11540
rect 23474 11500 23480 11512
rect 23532 11500 23538 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1762 11336 1768 11348
rect 1719 11308 1768 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 5166 11336 5172 11348
rect 5127 11308 5172 11336
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 6089 11339 6147 11345
rect 6089 11305 6101 11339
rect 6135 11336 6147 11339
rect 6822 11336 6828 11348
rect 6135 11308 6828 11336
rect 6135 11305 6147 11308
rect 6089 11299 6147 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7285 11339 7343 11345
rect 7285 11305 7297 11339
rect 7331 11336 7343 11339
rect 7374 11336 7380 11348
rect 7331 11308 7380 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 8389 11339 8447 11345
rect 8389 11305 8401 11339
rect 8435 11336 8447 11339
rect 8478 11336 8484 11348
rect 8435 11308 8484 11336
rect 8435 11305 8447 11308
rect 8389 11299 8447 11305
rect 8478 11296 8484 11308
rect 8536 11336 8542 11348
rect 8938 11336 8944 11348
rect 8536 11308 8944 11336
rect 8536 11296 8542 11308
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9306 11336 9312 11348
rect 9267 11308 9312 11336
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11057 11339 11115 11345
rect 11057 11305 11069 11339
rect 11103 11336 11115 11339
rect 11238 11336 11244 11348
rect 11103 11308 11244 11336
rect 11103 11305 11115 11308
rect 11057 11299 11115 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 14274 11296 14280 11348
rect 14332 11336 14338 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 14332 11308 14381 11336
rect 14332 11296 14338 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 15654 11296 15660 11348
rect 15712 11336 15718 11348
rect 15930 11336 15936 11348
rect 15712 11308 15936 11336
rect 15712 11296 15718 11308
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 16574 11296 16580 11348
rect 16632 11336 16638 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16632 11308 16681 11336
rect 16632 11296 16638 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 17313 11339 17371 11345
rect 17313 11305 17325 11339
rect 17359 11336 17371 11339
rect 18046 11336 18052 11348
rect 17359 11308 18052 11336
rect 17359 11305 17371 11308
rect 17313 11299 17371 11305
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 18138 11296 18144 11348
rect 18196 11336 18202 11348
rect 18196 11308 18241 11336
rect 18196 11296 18202 11308
rect 18598 11296 18604 11348
rect 18656 11296 18662 11348
rect 21177 11339 21235 11345
rect 21177 11305 21189 11339
rect 21223 11336 21235 11339
rect 21266 11336 21272 11348
rect 21223 11308 21272 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 23106 11296 23112 11348
rect 23164 11336 23170 11348
rect 23477 11339 23535 11345
rect 23477 11336 23489 11339
rect 23164 11308 23489 11336
rect 23164 11296 23170 11308
rect 23477 11305 23489 11308
rect 23523 11305 23535 11339
rect 24026 11336 24032 11348
rect 23987 11308 24032 11336
rect 23477 11299 23535 11305
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 24946 11296 24952 11348
rect 25004 11336 25010 11348
rect 25406 11336 25412 11348
rect 25004 11308 25412 11336
rect 25004 11296 25010 11308
rect 25406 11296 25412 11308
rect 25464 11296 25470 11348
rect 25590 11336 25596 11348
rect 25551 11308 25596 11336
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 7653 11271 7711 11277
rect 7653 11268 7665 11271
rect 7156 11240 7665 11268
rect 7156 11228 7162 11240
rect 7653 11237 7665 11240
rect 7699 11237 7711 11271
rect 7653 11231 7711 11237
rect 9677 11271 9735 11277
rect 9677 11237 9689 11271
rect 9723 11268 9735 11271
rect 10042 11268 10048 11280
rect 9723 11240 10048 11268
rect 9723 11237 9735 11240
rect 9677 11231 9735 11237
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 11146 11228 11152 11280
rect 11204 11268 11210 11280
rect 11517 11271 11575 11277
rect 11517 11268 11529 11271
rect 11204 11240 11529 11268
rect 11204 11228 11210 11240
rect 11517 11237 11529 11240
rect 11563 11268 11575 11271
rect 12250 11268 12256 11280
rect 11563 11240 12256 11268
rect 11563 11237 11575 11240
rect 11517 11231 11575 11237
rect 12250 11228 12256 11240
rect 12308 11228 12314 11280
rect 15562 11277 15568 11280
rect 15105 11271 15163 11277
rect 15105 11237 15117 11271
rect 15151 11268 15163 11271
rect 15556 11268 15568 11277
rect 15151 11240 15568 11268
rect 15151 11237 15163 11240
rect 15105 11231 15163 11237
rect 15556 11231 15568 11240
rect 15620 11268 15626 11280
rect 16022 11268 16028 11280
rect 15620 11240 16028 11268
rect 15562 11228 15568 11231
rect 15620 11228 15626 11240
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 17773 11271 17831 11277
rect 17773 11237 17785 11271
rect 17819 11268 17831 11271
rect 18616 11268 18644 11296
rect 17819 11240 18644 11268
rect 22005 11271 22063 11277
rect 17819 11237 17831 11240
rect 17773 11231 17831 11237
rect 22005 11237 22017 11271
rect 22051 11268 22063 11271
rect 22342 11271 22400 11277
rect 22342 11268 22354 11271
rect 22051 11240 22354 11268
rect 22051 11237 22063 11240
rect 22005 11231 22063 11237
rect 22342 11237 22354 11240
rect 22388 11268 22400 11271
rect 23290 11268 23296 11280
rect 22388 11240 23296 11268
rect 22388 11237 22400 11240
rect 22342 11231 22400 11237
rect 23290 11228 23296 11240
rect 23348 11228 23354 11280
rect 8386 11160 8392 11212
rect 8444 11200 8450 11212
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 8444 11172 8493 11200
rect 8444 11160 8450 11172
rect 8481 11169 8493 11172
rect 8527 11169 8539 11203
rect 8481 11163 8539 11169
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 11790 11200 11796 11212
rect 11471 11172 11796 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12989 11203 13047 11209
rect 12989 11200 13001 11203
rect 12492 11172 13001 11200
rect 12492 11160 12498 11172
rect 12989 11169 13001 11172
rect 13035 11169 13047 11203
rect 12989 11163 13047 11169
rect 14185 11203 14243 11209
rect 14185 11169 14197 11203
rect 14231 11169 14243 11203
rect 15286 11200 15292 11212
rect 15199 11172 15292 11200
rect 14185 11163 14243 11169
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 11698 11132 11704 11144
rect 8628 11104 8673 11132
rect 11659 11104 11704 11132
rect 8628 11092 8634 11104
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12894 11132 12900 11144
rect 12207 11104 12900 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12894 11092 12900 11104
rect 12952 11132 12958 11144
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12952 11104 13093 11132
rect 12952 11092 12958 11104
rect 13081 11101 13093 11104
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 13814 11132 13820 11144
rect 13228 11104 13820 11132
rect 13228 11092 13234 11104
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 5721 11067 5779 11073
rect 5721 11033 5733 11067
rect 5767 11064 5779 11067
rect 5994 11064 6000 11076
rect 5767 11036 6000 11064
rect 5767 11033 5779 11036
rect 5721 11027 5779 11033
rect 5994 11024 6000 11036
rect 6052 11064 6058 11076
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 6052 11036 8033 11064
rect 6052 11024 6058 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 10870 11064 10876 11076
rect 10831 11036 10876 11064
rect 8021 11027 8079 11033
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 11716 11064 11744 11092
rect 14200 11076 14228 11163
rect 15286 11160 15292 11172
rect 15344 11200 15350 11212
rect 15930 11200 15936 11212
rect 15344 11172 15936 11200
rect 15344 11160 15350 11172
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 18046 11160 18052 11212
rect 18104 11200 18110 11212
rect 18592 11203 18650 11209
rect 18592 11200 18604 11203
rect 18104 11172 18604 11200
rect 18104 11160 18110 11172
rect 18592 11169 18604 11172
rect 18638 11200 18650 11203
rect 19426 11200 19432 11212
rect 18638 11172 19432 11200
rect 18638 11169 18650 11172
rect 18592 11163 18650 11169
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 20993 11203 21051 11209
rect 20993 11169 21005 11203
rect 21039 11200 21051 11203
rect 24946 11200 24952 11212
rect 21039 11172 21680 11200
rect 24907 11172 24952 11200
rect 21039 11169 21051 11172
rect 20993 11163 21051 11169
rect 18322 11132 18328 11144
rect 18283 11104 18328 11132
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 11072 11036 11744 11064
rect 12621 11067 12679 11073
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 11072 10996 11100 11036
rect 12621 11033 12633 11067
rect 12667 11064 12679 11067
rect 14182 11064 14188 11076
rect 12667 11036 14188 11064
rect 12667 11033 12679 11036
rect 12621 11027 12679 11033
rect 14182 11024 14188 11036
rect 14240 11024 14246 11076
rect 19334 11024 19340 11076
rect 19392 11064 19398 11076
rect 19705 11067 19763 11073
rect 19705 11064 19717 11067
rect 19392 11036 19717 11064
rect 19392 11024 19398 11036
rect 19705 11033 19717 11036
rect 19751 11064 19763 11067
rect 20162 11064 20168 11076
rect 19751 11036 20168 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20162 11024 20168 11036
rect 20220 11064 20226 11076
rect 21652 11073 21680 11172
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 22097 11135 22155 11141
rect 22097 11101 22109 11135
rect 22143 11101 22155 11135
rect 22097 11095 22155 11101
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 20220 11036 20269 11064
rect 20220 11024 20226 11036
rect 20257 11033 20269 11036
rect 20303 11033 20315 11067
rect 20257 11027 20315 11033
rect 21637 11067 21695 11073
rect 21637 11033 21649 11067
rect 21683 11064 21695 11067
rect 21726 11064 21732 11076
rect 21683 11036 21732 11064
rect 21683 11033 21695 11036
rect 21637 11027 21695 11033
rect 21726 11024 21732 11036
rect 21784 11024 21790 11076
rect 12526 10996 12532 11008
rect 10836 10968 11100 10996
rect 12487 10968 12532 10996
rect 10836 10956 10842 10968
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 21910 10956 21916 11008
rect 21968 10996 21974 11008
rect 22112 10996 22140 11095
rect 24854 11092 24860 11144
rect 24912 11132 24918 11144
rect 25041 11135 25099 11141
rect 25041 11132 25053 11135
rect 24912 11104 25053 11132
rect 24912 11092 24918 11104
rect 25041 11101 25053 11104
rect 25087 11101 25099 11135
rect 25041 11095 25099 11101
rect 25133 11135 25191 11141
rect 25133 11101 25145 11135
rect 25179 11101 25191 11135
rect 25133 11095 25191 11101
rect 22462 10996 22468 11008
rect 21968 10968 22468 10996
rect 21968 10956 21974 10968
rect 22462 10956 22468 10968
rect 22520 10996 22526 11008
rect 23014 10996 23020 11008
rect 22520 10968 23020 10996
rect 22520 10956 22526 10968
rect 23014 10956 23020 10968
rect 23072 10956 23078 11008
rect 24118 10956 24124 11008
rect 24176 10996 24182 11008
rect 24581 10999 24639 11005
rect 24581 10996 24593 10999
rect 24176 10968 24593 10996
rect 24176 10956 24182 10968
rect 24581 10965 24593 10968
rect 24627 10965 24639 10999
rect 24581 10959 24639 10965
rect 25038 10956 25044 11008
rect 25096 10996 25102 11008
rect 25148 10996 25176 11095
rect 25096 10968 25176 10996
rect 25096 10956 25102 10968
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 8113 10795 8171 10801
rect 8113 10761 8125 10795
rect 8159 10792 8171 10795
rect 8202 10792 8208 10804
rect 8159 10764 8208 10792
rect 8159 10761 8171 10764
rect 8113 10755 8171 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8478 10792 8484 10804
rect 8439 10764 8484 10792
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 9214 10792 9220 10804
rect 9175 10764 9220 10792
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 9732 10764 10793 10792
rect 9732 10752 9738 10764
rect 10781 10761 10793 10764
rect 10827 10761 10839 10795
rect 10781 10755 10839 10761
rect 12158 10752 12164 10804
rect 12216 10792 12222 10804
rect 12253 10795 12311 10801
rect 12253 10792 12265 10795
rect 12216 10764 12265 10792
rect 12216 10752 12222 10764
rect 12253 10761 12265 10764
rect 12299 10792 12311 10795
rect 12618 10792 12624 10804
rect 12299 10764 12624 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 7745 10727 7803 10733
rect 7745 10693 7757 10727
rect 7791 10724 7803 10727
rect 8570 10724 8576 10736
rect 7791 10696 8576 10724
rect 7791 10693 7803 10696
rect 7745 10687 7803 10693
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 10321 10727 10379 10733
rect 10321 10693 10333 10727
rect 10367 10724 10379 10727
rect 11146 10724 11152 10736
rect 10367 10696 11152 10724
rect 10367 10693 10379 10696
rect 10321 10687 10379 10693
rect 11146 10684 11152 10696
rect 11204 10684 11210 10736
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9364 10628 9781 10656
rect 9364 10616 9370 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 11238 10656 11244 10668
rect 11199 10628 11244 10656
rect 9769 10619 9827 10625
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11425 10659 11483 10665
rect 11425 10625 11437 10659
rect 11471 10656 11483 10659
rect 11606 10656 11612 10668
rect 11471 10628 11612 10656
rect 11471 10625 11483 10628
rect 11425 10619 11483 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12452 10665 12480 10764
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 13814 10792 13820 10804
rect 13775 10764 13820 10792
rect 13814 10752 13820 10764
rect 13872 10792 13878 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 13872 10764 14381 10792
rect 13872 10752 13878 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 14369 10755 14427 10761
rect 16390 10752 16396 10804
rect 16448 10792 16454 10804
rect 17037 10795 17095 10801
rect 17037 10792 17049 10795
rect 16448 10764 17049 10792
rect 16448 10752 16454 10764
rect 17037 10761 17049 10764
rect 17083 10761 17095 10795
rect 17037 10755 17095 10761
rect 17954 10752 17960 10804
rect 18012 10792 18018 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 18012 10764 18245 10792
rect 18012 10752 18018 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 19242 10792 19248 10804
rect 18233 10755 18291 10761
rect 18708 10764 19248 10792
rect 17497 10727 17555 10733
rect 17497 10693 17509 10727
rect 17543 10724 17555 10727
rect 18046 10724 18052 10736
rect 17543 10696 18052 10724
rect 17543 10693 17555 10696
rect 17497 10687 17555 10693
rect 18046 10684 18052 10696
rect 18104 10684 18110 10736
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 15010 10616 15016 10668
rect 15068 10656 15074 10668
rect 18708 10665 18736 10764
rect 19242 10752 19248 10764
rect 19300 10792 19306 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19300 10764 19625 10792
rect 19300 10752 19306 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 20772 10764 20913 10792
rect 20772 10752 20778 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 23014 10792 23020 10804
rect 22975 10764 23020 10792
rect 20901 10755 20959 10761
rect 19978 10724 19984 10736
rect 19939 10696 19984 10724
rect 19978 10684 19984 10696
rect 20036 10684 20042 10736
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15068 10628 15485 10656
rect 15068 10616 15074 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10656 18843 10659
rect 19334 10656 19340 10668
rect 18831 10628 19340 10656
rect 18831 10625 18843 10628
rect 18785 10619 18843 10625
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9490 10588 9496 10600
rect 9171 10560 9496 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9490 10548 9496 10560
rect 9548 10588 9554 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 9548 10560 9597 10588
rect 9548 10548 9554 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 12693 10591 12751 10597
rect 12693 10588 12705 10591
rect 12584 10560 12705 10588
rect 12584 10548 12590 10560
rect 12693 10557 12705 10560
rect 12739 10557 12751 10591
rect 12693 10551 12751 10557
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 14875 10560 15332 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 15304 10532 15332 10560
rect 16684 10560 16865 10588
rect 10134 10480 10140 10532
rect 10192 10520 10198 10532
rect 10597 10523 10655 10529
rect 10597 10520 10609 10523
rect 10192 10492 10609 10520
rect 10192 10480 10198 10492
rect 10597 10489 10609 10492
rect 10643 10520 10655 10523
rect 11149 10523 11207 10529
rect 11149 10520 11161 10523
rect 10643 10492 11161 10520
rect 10643 10489 10655 10492
rect 10597 10483 10655 10489
rect 11149 10489 11161 10492
rect 11195 10489 11207 10523
rect 11149 10483 11207 10489
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 15286 10520 15292 10532
rect 13872 10492 14964 10520
rect 15247 10492 15292 10520
rect 13872 10480 13878 10492
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 9732 10424 9777 10452
rect 9732 10412 9738 10424
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 10870 10452 10876 10464
rect 10744 10424 10876 10452
rect 10744 10412 10750 10424
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 11790 10452 11796 10464
rect 11751 10424 11796 10452
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 14936 10461 14964 10492
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 16301 10523 16359 10529
rect 16301 10520 16313 10523
rect 15396 10492 16313 10520
rect 15396 10464 15424 10492
rect 16301 10489 16313 10492
rect 16347 10489 16359 10523
rect 16301 10483 16359 10489
rect 14921 10455 14979 10461
rect 14921 10421 14933 10455
rect 14967 10421 14979 10455
rect 14921 10415 14979 10421
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 16022 10452 16028 10464
rect 15436 10424 15481 10452
rect 15983 10424 16028 10452
rect 15436 10412 15442 10424
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16684 10461 16712 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 16853 10551 16911 10557
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18800 10588 18828 10619
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 20916 10656 20944 10755
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 23566 10792 23572 10804
rect 23523 10764 23572 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 23566 10752 23572 10764
rect 23624 10752 23630 10804
rect 23842 10752 23848 10804
rect 23900 10792 23906 10804
rect 24026 10792 24032 10804
rect 23900 10764 24032 10792
rect 23900 10752 23906 10764
rect 24026 10752 24032 10764
rect 24084 10752 24090 10804
rect 24946 10752 24952 10804
rect 25004 10792 25010 10804
rect 25041 10795 25099 10801
rect 25041 10792 25053 10795
rect 25004 10764 25053 10792
rect 25004 10752 25010 10764
rect 25041 10761 25053 10764
rect 25087 10761 25099 10795
rect 25041 10755 25099 10761
rect 25409 10795 25467 10801
rect 25409 10761 25421 10795
rect 25455 10792 25467 10795
rect 25498 10792 25504 10804
rect 25455 10764 25504 10792
rect 25455 10761 25467 10764
rect 25409 10755 25467 10761
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 21085 10659 21143 10665
rect 21085 10656 21097 10659
rect 20916 10628 21097 10656
rect 21085 10625 21097 10628
rect 21131 10625 21143 10659
rect 23584 10656 23612 10752
rect 23661 10727 23719 10733
rect 23661 10693 23673 10727
rect 23707 10724 23719 10727
rect 25314 10724 25320 10736
rect 23707 10696 25320 10724
rect 23707 10693 23719 10696
rect 23661 10687 23719 10693
rect 25314 10684 25320 10696
rect 25372 10684 25378 10736
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23584 10628 24225 10656
rect 21085 10619 21143 10625
rect 24213 10625 24225 10628
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 17911 10560 18828 10588
rect 19797 10591 19855 10597
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 19797 10557 19809 10591
rect 19843 10588 19855 10591
rect 20254 10588 20260 10600
rect 19843 10560 20260 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 24029 10591 24087 10597
rect 24029 10557 24041 10591
rect 24075 10588 24087 10591
rect 24118 10588 24124 10600
rect 24075 10560 24124 10588
rect 24075 10557 24087 10560
rect 24029 10551 24087 10557
rect 24118 10548 24124 10560
rect 24176 10548 24182 10600
rect 25222 10588 25228 10600
rect 25183 10560 25228 10588
rect 25222 10548 25228 10560
rect 25280 10588 25286 10600
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25280 10560 25789 10588
rect 25280 10548 25286 10560
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 20625 10523 20683 10529
rect 20625 10489 20637 10523
rect 20671 10520 20683 10523
rect 21352 10523 21410 10529
rect 21352 10520 21364 10523
rect 20671 10492 21364 10520
rect 20671 10489 20683 10492
rect 20625 10483 20683 10489
rect 21352 10489 21364 10492
rect 21398 10520 21410 10523
rect 21450 10520 21456 10532
rect 21398 10492 21456 10520
rect 21398 10489 21410 10492
rect 21352 10483 21410 10489
rect 21450 10480 21456 10492
rect 21508 10480 21514 10532
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 16632 10424 16681 10452
rect 16632 10412 16638 10424
rect 16669 10421 16681 10424
rect 16715 10421 16727 10455
rect 18598 10452 18604 10464
rect 18559 10424 18604 10452
rect 16669 10415 16727 10421
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 18966 10412 18972 10464
rect 19024 10452 19030 10464
rect 19245 10455 19303 10461
rect 19245 10452 19257 10455
rect 19024 10424 19257 10452
rect 19024 10412 19030 10424
rect 19245 10421 19257 10424
rect 19291 10421 19303 10455
rect 19245 10415 19303 10421
rect 22186 10412 22192 10464
rect 22244 10452 22250 10464
rect 22465 10455 22523 10461
rect 22465 10452 22477 10455
rect 22244 10424 22477 10452
rect 22244 10412 22250 10424
rect 22465 10421 22477 10424
rect 22511 10421 22523 10455
rect 22465 10415 22523 10421
rect 23842 10412 23848 10464
rect 23900 10452 23906 10464
rect 24121 10455 24179 10461
rect 24121 10452 24133 10455
rect 23900 10424 24133 10452
rect 23900 10412 23906 10424
rect 24121 10421 24133 10424
rect 24167 10421 24179 10455
rect 24121 10415 24179 10421
rect 24210 10412 24216 10464
rect 24268 10452 24274 10464
rect 24673 10455 24731 10461
rect 24673 10452 24685 10455
rect 24268 10424 24685 10452
rect 24268 10412 24274 10424
rect 24673 10421 24685 10424
rect 24719 10452 24731 10455
rect 24854 10452 24860 10464
rect 24719 10424 24860 10452
rect 24719 10421 24731 10424
rect 24673 10415 24731 10421
rect 24854 10412 24860 10424
rect 24912 10412 24918 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 9306 10248 9312 10260
rect 9267 10220 9312 10248
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10686 10248 10692 10260
rect 10183 10220 10692 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10686 10208 10692 10220
rect 10744 10248 10750 10260
rect 10962 10248 10968 10260
rect 10744 10220 10968 10248
rect 10744 10208 10750 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11606 10248 11612 10260
rect 11567 10220 11612 10248
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 14182 10248 14188 10260
rect 14143 10220 14188 10248
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 15010 10248 15016 10260
rect 14971 10220 15016 10248
rect 15010 10208 15016 10220
rect 15068 10248 15074 10260
rect 15286 10248 15292 10260
rect 15068 10220 15292 10248
rect 15068 10208 15074 10220
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15562 10248 15568 10260
rect 15523 10220 15568 10248
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 23014 10208 23020 10260
rect 23072 10248 23078 10260
rect 23290 10248 23296 10260
rect 23072 10220 23296 10248
rect 23072 10208 23078 10220
rect 23290 10208 23296 10220
rect 23348 10208 23354 10260
rect 24118 10208 24124 10260
rect 24176 10248 24182 10260
rect 24213 10251 24271 10257
rect 24213 10248 24225 10251
rect 24176 10220 24225 10248
rect 24176 10208 24182 10220
rect 24213 10217 24225 10220
rect 24259 10217 24271 10251
rect 24213 10211 24271 10217
rect 24578 10208 24584 10260
rect 24636 10248 24642 10260
rect 25038 10248 25044 10260
rect 24636 10220 25044 10248
rect 24636 10208 24642 10220
rect 25038 10208 25044 10220
rect 25096 10248 25102 10260
rect 25409 10251 25467 10257
rect 25409 10248 25421 10251
rect 25096 10220 25421 10248
rect 25096 10208 25102 10220
rect 25409 10217 25421 10220
rect 25455 10217 25467 10251
rect 25409 10211 25467 10217
rect 10505 10183 10563 10189
rect 10505 10149 10517 10183
rect 10551 10180 10563 10183
rect 10778 10180 10784 10192
rect 10551 10152 10784 10180
rect 10551 10149 10563 10152
rect 10505 10143 10563 10149
rect 10778 10140 10784 10152
rect 10836 10140 10842 10192
rect 12428 10183 12486 10189
rect 12428 10149 12440 10183
rect 12474 10180 12486 10183
rect 15028 10180 15056 10208
rect 12474 10152 15056 10180
rect 16292 10183 16350 10189
rect 12474 10149 12486 10152
rect 12428 10143 12486 10149
rect 16292 10149 16304 10183
rect 16338 10180 16350 10183
rect 16390 10180 16396 10192
rect 16338 10152 16396 10180
rect 16338 10149 16350 10152
rect 16292 10143 16350 10149
rect 16390 10140 16396 10152
rect 16448 10140 16454 10192
rect 20901 10183 20959 10189
rect 20901 10149 20913 10183
rect 20947 10180 20959 10183
rect 24765 10183 24823 10189
rect 24765 10180 24777 10183
rect 20947 10152 24777 10180
rect 20947 10149 20959 10152
rect 20901 10143 20959 10149
rect 24765 10149 24777 10152
rect 24811 10180 24823 10183
rect 24854 10180 24860 10192
rect 24811 10152 24860 10180
rect 24811 10149 24823 10152
rect 24765 10143 24823 10149
rect 24854 10140 24860 10152
rect 24912 10140 24918 10192
rect 10962 10112 10968 10124
rect 10923 10084 10968 10112
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 11514 10112 11520 10124
rect 11103 10084 11520 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 12158 10112 12164 10124
rect 12119 10084 12164 10112
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 16022 10112 16028 10124
rect 15983 10084 16028 10112
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 18966 10072 18972 10124
rect 19024 10112 19030 10124
rect 22186 10121 22192 10124
rect 19153 10115 19211 10121
rect 19153 10112 19165 10115
rect 19024 10084 19165 10112
rect 19024 10072 19030 10084
rect 19153 10081 19165 10084
rect 19199 10081 19211 10115
rect 19153 10075 19211 10081
rect 21729 10115 21787 10121
rect 21729 10081 21741 10115
rect 21775 10112 21787 10115
rect 22180 10112 22192 10121
rect 21775 10084 22192 10112
rect 21775 10081 21787 10084
rect 21729 10075 21787 10081
rect 22180 10075 22192 10084
rect 22244 10112 22250 10124
rect 24118 10112 24124 10124
rect 22244 10084 24124 10112
rect 22186 10072 22192 10075
rect 22244 10072 22250 10084
rect 24118 10072 24124 10084
rect 24176 10112 24182 10124
rect 24176 10084 24992 10112
rect 24176 10072 24182 10084
rect 11238 10044 11244 10056
rect 11199 10016 11244 10044
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 18049 10047 18107 10053
rect 18049 10013 18061 10047
rect 18095 10044 18107 10047
rect 19242 10044 19248 10056
rect 18095 10016 19248 10044
rect 18095 10013 18107 10016
rect 18049 10007 18107 10013
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 19426 10044 19432 10056
rect 19387 10016 19432 10044
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 21910 10044 21916 10056
rect 20772 10016 21916 10044
rect 20772 10004 20778 10016
rect 21910 10004 21916 10016
rect 21968 10004 21974 10056
rect 24964 10053 24992 10084
rect 24857 10047 24915 10053
rect 24857 10013 24869 10047
rect 24903 10013 24915 10047
rect 24857 10007 24915 10013
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10013 25007 10047
rect 24949 10007 25007 10013
rect 8941 9979 8999 9985
rect 8941 9945 8953 9979
rect 8987 9976 8999 9979
rect 9582 9976 9588 9988
rect 8987 9948 9588 9976
rect 8987 9945 8999 9948
rect 8941 9939 8999 9945
rect 9582 9936 9588 9948
rect 9640 9936 9646 9988
rect 10597 9979 10655 9985
rect 10597 9945 10609 9979
rect 10643 9976 10655 9979
rect 11977 9979 12035 9985
rect 11977 9976 11989 9979
rect 10643 9948 11989 9976
rect 10643 9945 10655 9948
rect 10597 9939 10655 9945
rect 11977 9945 11989 9948
rect 12023 9945 12035 9979
rect 11977 9939 12035 9945
rect 11992 9908 12020 9939
rect 18598 9936 18604 9988
rect 18656 9976 18662 9988
rect 18785 9979 18843 9985
rect 18785 9976 18797 9979
rect 18656 9948 18797 9976
rect 18656 9936 18662 9948
rect 18785 9945 18797 9948
rect 18831 9976 18843 9979
rect 19797 9979 19855 9985
rect 19797 9976 19809 9979
rect 18831 9948 19809 9976
rect 18831 9945 18843 9948
rect 18785 9939 18843 9945
rect 19797 9945 19809 9948
rect 19843 9945 19855 9979
rect 19797 9939 19855 9945
rect 23106 9936 23112 9988
rect 23164 9976 23170 9988
rect 24397 9979 24455 9985
rect 24397 9976 24409 9979
rect 23164 9948 24409 9976
rect 23164 9936 23170 9948
rect 24397 9945 24409 9948
rect 24443 9945 24455 9979
rect 24397 9939 24455 9945
rect 12342 9908 12348 9920
rect 11992 9880 12348 9908
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 13446 9908 13452 9920
rect 12584 9880 13452 9908
rect 12584 9868 12590 9880
rect 13446 9868 13452 9880
rect 13504 9908 13510 9920
rect 13541 9911 13599 9917
rect 13541 9908 13553 9911
rect 13504 9880 13553 9908
rect 13504 9868 13510 9880
rect 13541 9877 13553 9880
rect 13587 9877 13599 9911
rect 13541 9871 13599 9877
rect 17405 9911 17463 9917
rect 17405 9877 17417 9911
rect 17451 9908 17463 9911
rect 17678 9908 17684 9920
rect 17451 9880 17684 9908
rect 17451 9877 17463 9880
rect 17405 9871 17463 9877
rect 17678 9868 17684 9880
rect 17736 9868 17742 9920
rect 18322 9908 18328 9920
rect 18283 9880 18328 9908
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 20254 9908 20260 9920
rect 20215 9880 20260 9908
rect 20254 9868 20260 9880
rect 20312 9868 20318 9920
rect 23842 9908 23848 9920
rect 23803 9880 23848 9908
rect 23842 9868 23848 9880
rect 23900 9868 23906 9920
rect 24872 9908 24900 10007
rect 24946 9908 24952 9920
rect 24872 9880 24952 9908
rect 24946 9868 24952 9880
rect 25004 9908 25010 9920
rect 25682 9908 25688 9920
rect 25004 9880 25688 9908
rect 25004 9868 25010 9880
rect 25682 9868 25688 9880
rect 25740 9868 25746 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 12158 9704 12164 9716
rect 12119 9676 12164 9704
rect 12158 9664 12164 9676
rect 12216 9704 12222 9716
rect 12802 9704 12808 9716
rect 12216 9676 12808 9704
rect 12216 9664 12222 9676
rect 12802 9664 12808 9676
rect 12860 9704 12866 9716
rect 13541 9707 13599 9713
rect 13541 9704 13553 9707
rect 12860 9676 13553 9704
rect 12860 9664 12866 9676
rect 13541 9673 13553 9676
rect 13587 9673 13599 9707
rect 13541 9667 13599 9673
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 10045 9639 10103 9645
rect 10045 9636 10057 9639
rect 9732 9608 10057 9636
rect 9732 9596 9738 9608
rect 10045 9605 10057 9608
rect 10091 9605 10103 9639
rect 10045 9599 10103 9605
rect 11149 9639 11207 9645
rect 11149 9605 11161 9639
rect 11195 9636 11207 9639
rect 11238 9636 11244 9648
rect 11195 9608 11244 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 11238 9596 11244 9608
rect 11296 9636 11302 9648
rect 12526 9636 12532 9648
rect 11296 9608 12532 9636
rect 11296 9596 11302 9608
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10134 9568 10140 9580
rect 10008 9540 10140 9568
rect 10008 9528 10014 9540
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10686 9568 10692 9580
rect 10647 9540 10692 9568
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 13556 9568 13584 9667
rect 14734 9664 14740 9716
rect 14792 9704 14798 9716
rect 15105 9707 15163 9713
rect 15105 9704 15117 9707
rect 14792 9676 15117 9704
rect 14792 9664 14798 9676
rect 15105 9673 15117 9676
rect 15151 9704 15163 9707
rect 15286 9704 15292 9716
rect 15151 9676 15292 9704
rect 15151 9673 15163 9676
rect 15105 9667 15163 9673
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 16390 9664 16396 9716
rect 16448 9704 16454 9716
rect 16448 9676 16528 9704
rect 16448 9664 16454 9676
rect 16206 9636 16212 9648
rect 16167 9608 16212 9636
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 16500 9636 16528 9676
rect 16758 9664 16764 9716
rect 16816 9704 16822 9716
rect 16942 9704 16948 9716
rect 16816 9676 16948 9704
rect 16816 9664 16822 9676
rect 16942 9664 16948 9676
rect 17000 9664 17006 9716
rect 17770 9704 17776 9716
rect 17604 9676 17776 9704
rect 17221 9639 17279 9645
rect 17221 9636 17233 9639
rect 16500 9608 17233 9636
rect 17221 9605 17233 9608
rect 17267 9605 17279 9639
rect 17604 9636 17632 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 21910 9664 21916 9716
rect 21968 9704 21974 9716
rect 22649 9707 22707 9713
rect 22649 9704 22661 9707
rect 21968 9676 22661 9704
rect 21968 9664 21974 9676
rect 22649 9673 22661 9676
rect 22695 9673 22707 9707
rect 22649 9667 22707 9673
rect 23014 9664 23020 9716
rect 23072 9704 23078 9716
rect 23290 9704 23296 9716
rect 23072 9676 23296 9704
rect 23072 9664 23078 9676
rect 23290 9664 23296 9676
rect 23348 9664 23354 9716
rect 23658 9704 23664 9716
rect 23492 9676 23664 9704
rect 18230 9636 18236 9648
rect 17604 9608 18236 9636
rect 17221 9599 17279 9605
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 20257 9639 20315 9645
rect 20257 9636 20269 9639
rect 19484 9608 20269 9636
rect 19484 9596 19490 9608
rect 20257 9605 20269 9608
rect 20303 9605 20315 9639
rect 20257 9599 20315 9605
rect 20438 9596 20444 9648
rect 20496 9636 20502 9648
rect 20496 9608 23428 9636
rect 20496 9596 20502 9608
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13556 9540 13737 9568
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 16850 9568 16856 9580
rect 16811 9540 16856 9568
rect 13725 9531 13783 9537
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 22186 9568 22192 9580
rect 22147 9540 22192 9568
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 10100 9472 10517 9500
rect 10100 9460 10106 9472
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 15749 9503 15807 9509
rect 15749 9500 15761 9503
rect 10505 9463 10563 9469
rect 10612 9472 15761 9500
rect 9950 9392 9956 9444
rect 10008 9432 10014 9444
rect 10612 9432 10640 9472
rect 15749 9469 15761 9472
rect 15795 9500 15807 9503
rect 16577 9503 16635 9509
rect 16577 9500 16589 9503
rect 15795 9472 16589 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 16577 9469 16589 9472
rect 16623 9500 16635 9503
rect 17034 9500 17040 9512
rect 16623 9472 17040 9500
rect 16623 9469 16635 9472
rect 16577 9463 16635 9469
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 18322 9500 18328 9512
rect 17788 9472 18328 9500
rect 10008 9404 10640 9432
rect 13265 9435 13323 9441
rect 10008 9392 10014 9404
rect 13265 9401 13277 9435
rect 13311 9432 13323 9435
rect 13992 9435 14050 9441
rect 13992 9432 14004 9435
rect 13311 9404 14004 9432
rect 13311 9401 13323 9404
rect 13265 9395 13323 9401
rect 13992 9401 14004 9404
rect 14038 9432 14050 9435
rect 14274 9432 14280 9444
rect 14038 9404 14280 9432
rect 14038 9401 14050 9404
rect 13992 9395 14050 9401
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 16117 9435 16175 9441
rect 16117 9401 16129 9435
rect 16163 9432 16175 9435
rect 16163 9404 16712 9432
rect 16163 9401 16175 9404
rect 16117 9395 16175 9401
rect 9858 9364 9864 9376
rect 9819 9336 9864 9364
rect 9858 9324 9864 9336
rect 9916 9364 9922 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 9916 9336 10425 9364
rect 9916 9324 9922 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 11514 9364 11520 9376
rect 11475 9336 11520 9364
rect 10413 9327 10471 9333
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 11885 9367 11943 9373
rect 11885 9333 11897 9367
rect 11931 9364 11943 9367
rect 12342 9364 12348 9376
rect 11931 9336 12348 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 12526 9364 12532 9376
rect 12487 9336 12532 9364
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 16684 9373 16712 9404
rect 16669 9367 16727 9373
rect 16669 9333 16681 9367
rect 16715 9364 16727 9367
rect 16942 9364 16948 9376
rect 16715 9336 16948 9364
rect 16715 9333 16727 9336
rect 16669 9327 16727 9333
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17126 9324 17132 9376
rect 17184 9364 17190 9376
rect 17788 9373 17816 9472
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 21545 9503 21603 9509
rect 21545 9469 21557 9503
rect 21591 9500 21603 9503
rect 22002 9500 22008 9512
rect 21591 9472 22008 9500
rect 21591 9469 21603 9472
rect 21545 9463 21603 9469
rect 22002 9460 22008 9472
rect 22060 9460 22066 9512
rect 18506 9392 18512 9444
rect 18564 9441 18570 9444
rect 18564 9435 18628 9441
rect 18564 9401 18582 9435
rect 18616 9401 18628 9435
rect 18564 9395 18628 9401
rect 18564 9392 18570 9395
rect 20898 9392 20904 9444
rect 20956 9432 20962 9444
rect 21177 9435 21235 9441
rect 21177 9432 21189 9435
rect 20956 9404 21189 9432
rect 20956 9392 20962 9404
rect 21177 9401 21189 9404
rect 21223 9432 21235 9435
rect 22097 9435 22155 9441
rect 22097 9432 22109 9435
rect 21223 9404 22109 9432
rect 21223 9401 21235 9404
rect 21177 9395 21235 9401
rect 22097 9401 22109 9404
rect 22143 9401 22155 9435
rect 23400 9432 23428 9608
rect 23492 9500 23520 9676
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 24118 9704 24124 9716
rect 24079 9676 24124 9704
rect 24118 9664 24124 9676
rect 24176 9664 24182 9716
rect 24670 9596 24676 9648
rect 24728 9636 24734 9648
rect 24765 9639 24823 9645
rect 24765 9636 24777 9639
rect 24728 9608 24777 9636
rect 24728 9596 24734 9608
rect 24765 9605 24777 9608
rect 24811 9605 24823 9639
rect 24765 9599 24823 9605
rect 24854 9596 24860 9648
rect 24912 9636 24918 9648
rect 25133 9639 25191 9645
rect 25133 9636 25145 9639
rect 24912 9608 25145 9636
rect 24912 9596 24918 9608
rect 25133 9605 25145 9608
rect 25179 9605 25191 9639
rect 25133 9599 25191 9605
rect 23658 9500 23664 9512
rect 23492 9472 23664 9500
rect 23658 9460 23664 9472
rect 23716 9460 23722 9512
rect 23934 9460 23940 9512
rect 23992 9500 23998 9512
rect 24581 9503 24639 9509
rect 24581 9500 24593 9503
rect 23992 9472 24593 9500
rect 23992 9460 23998 9472
rect 24581 9469 24593 9472
rect 24627 9500 24639 9503
rect 25501 9503 25559 9509
rect 25501 9500 25513 9503
rect 24627 9472 25513 9500
rect 24627 9469 24639 9472
rect 24581 9463 24639 9469
rect 25501 9469 25513 9472
rect 25547 9469 25559 9503
rect 25501 9463 25559 9469
rect 24397 9435 24455 9441
rect 24397 9432 24409 9435
rect 23400 9404 24409 9432
rect 22097 9395 22155 9401
rect 24397 9401 24409 9404
rect 24443 9432 24455 9435
rect 24946 9432 24952 9444
rect 24443 9404 24952 9432
rect 24443 9401 24455 9404
rect 24397 9395 24455 9401
rect 24946 9392 24952 9404
rect 25004 9392 25010 9444
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17184 9336 17785 9364
rect 17184 9324 17190 9336
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 17773 9327 17831 9333
rect 19518 9324 19524 9376
rect 19576 9364 19582 9376
rect 19705 9367 19763 9373
rect 19705 9364 19717 9367
rect 19576 9336 19717 9364
rect 19576 9324 19582 9336
rect 19705 9333 19717 9336
rect 19751 9364 19763 9367
rect 20530 9364 20536 9376
rect 19751 9336 20536 9364
rect 19751 9333 19763 9336
rect 19705 9327 19763 9333
rect 20530 9324 20536 9336
rect 20588 9364 20594 9376
rect 21082 9364 21088 9376
rect 20588 9336 21088 9364
rect 20588 9324 20594 9336
rect 21082 9324 21088 9336
rect 21140 9324 21146 9376
rect 21634 9364 21640 9376
rect 21595 9336 21640 9364
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 10042 9160 10048 9172
rect 10003 9132 10048 9160
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 10689 9163 10747 9169
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 10962 9160 10968 9172
rect 10735 9132 10968 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 10962 9120 10968 9132
rect 11020 9160 11026 9172
rect 11977 9163 12035 9169
rect 11977 9160 11989 9163
rect 11020 9132 11989 9160
rect 11020 9120 11026 9132
rect 11977 9129 11989 9132
rect 12023 9129 12035 9163
rect 11977 9123 12035 9129
rect 12066 9120 12072 9172
rect 12124 9160 12130 9172
rect 12437 9163 12495 9169
rect 12437 9160 12449 9163
rect 12124 9132 12449 9160
rect 12124 9120 12130 9132
rect 12437 9129 12449 9132
rect 12483 9129 12495 9163
rect 12437 9123 12495 9129
rect 13081 9163 13139 9169
rect 13081 9129 13093 9163
rect 13127 9160 13139 9163
rect 13722 9160 13728 9172
rect 13127 9132 13728 9160
rect 13127 9129 13139 9132
rect 13081 9123 13139 9129
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 13909 9163 13967 9169
rect 13909 9160 13921 9163
rect 13832 9132 13921 9160
rect 13832 9036 13860 9132
rect 13909 9129 13921 9132
rect 13955 9160 13967 9163
rect 14642 9160 14648 9172
rect 13955 9132 14648 9160
rect 13955 9129 13967 9132
rect 13909 9123 13967 9129
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 15565 9163 15623 9169
rect 15565 9129 15577 9163
rect 15611 9160 15623 9163
rect 16482 9160 16488 9172
rect 15611 9132 16488 9160
rect 15611 9129 15623 9132
rect 15565 9123 15623 9129
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16850 9120 16856 9172
rect 16908 9160 16914 9172
rect 16945 9163 17003 9169
rect 16945 9160 16957 9163
rect 16908 9132 16957 9160
rect 16908 9120 16914 9132
rect 16945 9129 16957 9132
rect 16991 9129 17003 9163
rect 19518 9160 19524 9172
rect 19479 9132 19524 9160
rect 16945 9123 17003 9129
rect 19518 9120 19524 9132
rect 19576 9120 19582 9172
rect 20530 9160 20536 9172
rect 20491 9132 20536 9160
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 20898 9160 20904 9172
rect 20859 9132 20904 9160
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 21634 9120 21640 9172
rect 21692 9160 21698 9172
rect 22462 9160 22468 9172
rect 21692 9132 22324 9160
rect 22423 9132 22468 9160
rect 21692 9120 21698 9132
rect 14550 9092 14556 9104
rect 14511 9064 14556 9092
rect 14550 9052 14556 9064
rect 14608 9052 14614 9104
rect 22005 9095 22063 9101
rect 22005 9061 22017 9095
rect 22051 9092 22063 9095
rect 22186 9092 22192 9104
rect 22051 9064 22192 9092
rect 22051 9061 22063 9064
rect 22005 9055 22063 9061
rect 22186 9052 22192 9064
rect 22244 9052 22250 9104
rect 22296 9092 22324 9132
rect 22462 9120 22468 9132
rect 22520 9120 22526 9172
rect 22833 9163 22891 9169
rect 22833 9129 22845 9163
rect 22879 9160 22891 9163
rect 23106 9160 23112 9172
rect 22879 9132 23112 9160
rect 22879 9129 22891 9132
rect 22833 9123 22891 9129
rect 23106 9120 23112 9132
rect 23164 9120 23170 9172
rect 24762 9160 24768 9172
rect 24723 9132 24768 9160
rect 24762 9120 24768 9132
rect 24820 9120 24826 9172
rect 22922 9092 22928 9104
rect 22296 9064 22928 9092
rect 22922 9052 22928 9064
rect 22980 9052 22986 9104
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 9732 8996 10977 9024
rect 9732 8984 9738 8996
rect 10965 8993 10977 8996
rect 11011 8993 11023 9027
rect 10965 8987 11023 8993
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 9024 12403 9027
rect 12526 9024 12532 9036
rect 12391 8996 12532 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 13814 8984 13820 9036
rect 13872 8984 13878 9036
rect 13906 8984 13912 9036
rect 13964 9024 13970 9036
rect 14001 9027 14059 9033
rect 14001 9024 14013 9027
rect 13964 8996 14013 9024
rect 13964 8984 13970 8996
rect 14001 8993 14013 8996
rect 14047 8993 14059 9027
rect 15930 9024 15936 9036
rect 15891 8996 15936 9024
rect 14001 8987 14059 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 17396 9027 17454 9033
rect 17396 8993 17408 9027
rect 17442 9024 17454 9027
rect 17770 9024 17776 9036
rect 17442 8996 17776 9024
rect 17442 8993 17454 8996
rect 17396 8987 17454 8993
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 21266 9024 21272 9036
rect 21227 8996 21272 9024
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 23842 8984 23848 9036
rect 23900 9024 23906 9036
rect 24581 9027 24639 9033
rect 24581 9024 24593 9027
rect 23900 8996 24593 9024
rect 23900 8984 23906 8996
rect 24581 8993 24593 8996
rect 24627 9024 24639 9027
rect 25038 9024 25044 9036
rect 24627 8996 25044 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 25038 8984 25044 8996
rect 25096 8984 25102 9036
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8956 12679 8959
rect 14185 8959 14243 8965
rect 12667 8928 14136 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 12636 8888 12664 8919
rect 13538 8888 13544 8900
rect 12400 8860 12664 8888
rect 13499 8860 13544 8888
rect 12400 8848 12406 8860
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 14108 8888 14136 8928
rect 14185 8925 14197 8959
rect 14231 8956 14243 8959
rect 14274 8956 14280 8968
rect 14231 8928 14280 8956
rect 14231 8925 14243 8928
rect 14185 8919 14243 8925
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8956 15163 8959
rect 16022 8956 16028 8968
rect 15151 8928 16028 8956
rect 15151 8925 15163 8928
rect 15105 8919 15163 8925
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 16114 8916 16120 8968
rect 16172 8956 16178 8968
rect 17126 8956 17132 8968
rect 16172 8928 16217 8956
rect 16592 8928 17132 8956
rect 16172 8916 16178 8928
rect 14734 8888 14740 8900
rect 14108 8860 14740 8888
rect 14734 8848 14740 8860
rect 14792 8848 14798 8900
rect 16592 8832 16620 8928
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 19610 8956 19616 8968
rect 19571 8928 19616 8956
rect 19610 8916 19616 8928
rect 19668 8916 19674 8968
rect 19886 8916 19892 8968
rect 19944 8956 19950 8968
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 19944 8928 21373 8956
rect 19944 8916 19950 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 23109 8959 23167 8965
rect 21508 8928 21553 8956
rect 21508 8916 21514 8928
rect 23109 8925 23121 8959
rect 23155 8956 23167 8959
rect 23290 8956 23296 8968
rect 23155 8928 23296 8956
rect 23155 8925 23167 8928
rect 23109 8919 23167 8925
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 18506 8888 18512 8900
rect 18467 8860 18512 8888
rect 18506 8848 18512 8860
rect 18564 8888 18570 8900
rect 19061 8891 19119 8897
rect 19061 8888 19073 8891
rect 18564 8860 19073 8888
rect 18564 8848 18570 8860
rect 19061 8857 19073 8860
rect 19107 8857 19119 8891
rect 19061 8851 19119 8857
rect 13354 8820 13360 8832
rect 13315 8792 13360 8820
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 16574 8820 16580 8832
rect 16535 8792 16580 8820
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 12621 8619 12679 8625
rect 12621 8616 12633 8619
rect 12584 8588 12633 8616
rect 12584 8576 12590 8588
rect 12621 8585 12633 8588
rect 12667 8585 12679 8619
rect 12894 8616 12900 8628
rect 12855 8588 12900 8616
rect 12621 8579 12679 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13906 8616 13912 8628
rect 13867 8588 13912 8616
rect 13906 8576 13912 8588
rect 13964 8616 13970 8628
rect 15378 8616 15384 8628
rect 13964 8588 15384 8616
rect 13964 8576 13970 8588
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15657 8619 15715 8625
rect 15657 8585 15669 8619
rect 15703 8616 15715 8619
rect 16114 8616 16120 8628
rect 15703 8588 16120 8616
rect 15703 8585 15715 8588
rect 15657 8579 15715 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 17184 8588 17417 8616
rect 17184 8576 17190 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 18966 8616 18972 8628
rect 18927 8588 18972 8616
rect 17405 8579 17463 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 19392 8588 20545 8616
rect 19392 8576 19398 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 21266 8576 21272 8628
rect 21324 8616 21330 8628
rect 21545 8619 21603 8625
rect 21545 8616 21557 8619
rect 21324 8588 21557 8616
rect 21324 8576 21330 8588
rect 21545 8585 21557 8588
rect 21591 8585 21603 8619
rect 22922 8616 22928 8628
rect 22883 8588 22928 8616
rect 21545 8579 21603 8585
rect 22922 8576 22928 8588
rect 22980 8576 22986 8628
rect 23106 8576 23112 8628
rect 23164 8616 23170 8628
rect 23385 8619 23443 8625
rect 23385 8616 23397 8619
rect 23164 8588 23397 8616
rect 23164 8576 23170 8588
rect 23385 8585 23397 8588
rect 23431 8585 23443 8619
rect 23385 8579 23443 8585
rect 24026 8576 24032 8628
rect 24084 8616 24090 8628
rect 24121 8619 24179 8625
rect 24121 8616 24133 8619
rect 24084 8588 24133 8616
rect 24084 8576 24090 8588
rect 24121 8585 24133 8588
rect 24167 8585 24179 8619
rect 24854 8616 24860 8628
rect 24815 8588 24860 8616
rect 24121 8579 24179 8585
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25038 8576 25044 8628
rect 25096 8616 25102 8628
rect 25133 8619 25191 8625
rect 25133 8616 25145 8619
rect 25096 8588 25145 8616
rect 25096 8576 25102 8588
rect 25133 8585 25145 8588
rect 25179 8585 25191 8619
rect 25133 8579 25191 8585
rect 13354 8508 13360 8560
rect 13412 8548 13418 8560
rect 14461 8551 14519 8557
rect 14461 8548 14473 8551
rect 13412 8520 14473 8548
rect 13412 8508 13418 8520
rect 14461 8517 14473 8520
rect 14507 8517 14519 8551
rect 14461 8511 14519 8517
rect 14826 8508 14832 8560
rect 14884 8548 14890 8560
rect 15930 8548 15936 8560
rect 14884 8520 15936 8548
rect 14884 8508 14890 8520
rect 15930 8508 15936 8520
rect 15988 8548 15994 8560
rect 16393 8551 16451 8557
rect 16393 8548 16405 8551
rect 15988 8520 16405 8548
rect 15988 8508 15994 8520
rect 16393 8517 16405 8520
rect 16439 8517 16451 8551
rect 16393 8511 16451 8517
rect 19886 8508 19892 8560
rect 19944 8548 19950 8560
rect 19981 8551 20039 8557
rect 19981 8548 19993 8551
rect 19944 8520 19993 8548
rect 19944 8508 19950 8520
rect 19981 8517 19993 8520
rect 20027 8517 20039 8551
rect 19981 8511 20039 8517
rect 22649 8551 22707 8557
rect 22649 8517 22661 8551
rect 22695 8548 22707 8551
rect 23290 8548 23296 8560
rect 22695 8520 23296 8548
rect 22695 8517 22707 8520
rect 22649 8511 22707 8517
rect 23290 8508 23296 8520
rect 23348 8508 23354 8560
rect 23845 8551 23903 8557
rect 23845 8517 23857 8551
rect 23891 8548 23903 8551
rect 25406 8548 25412 8560
rect 23891 8520 25412 8548
rect 23891 8517 23903 8520
rect 23845 8511 23903 8517
rect 25406 8508 25412 8520
rect 25464 8508 25470 8560
rect 11330 8480 11336 8492
rect 11291 8452 11336 8480
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 13446 8480 13452 8492
rect 13407 8452 13452 8480
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 14734 8440 14740 8492
rect 14792 8480 14798 8492
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14792 8452 15025 8480
rect 14792 8440 14798 8452
rect 15013 8449 15025 8452
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16356 8452 16957 8480
rect 16356 8440 16362 8452
rect 16945 8449 16957 8452
rect 16991 8480 17003 8483
rect 17770 8480 17776 8492
rect 16991 8452 17776 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 17770 8440 17776 8452
rect 17828 8440 17834 8492
rect 19518 8480 19524 8492
rect 19479 8452 19524 8480
rect 19518 8440 19524 8452
rect 19576 8440 19582 8492
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 20898 8480 20904 8492
rect 20680 8452 20904 8480
rect 20680 8440 20686 8452
rect 20898 8440 20904 8452
rect 20956 8480 20962 8492
rect 20993 8483 21051 8489
rect 20993 8480 21005 8483
rect 20956 8452 21005 8480
rect 20956 8440 20962 8452
rect 20993 8449 21005 8452
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 21082 8440 21088 8492
rect 21140 8480 21146 8492
rect 21140 8452 21185 8480
rect 21140 8440 21146 8452
rect 22094 8440 22100 8492
rect 22152 8480 22158 8492
rect 22152 8452 22197 8480
rect 22152 8440 22158 8452
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8412 13323 8415
rect 13354 8412 13360 8424
rect 13311 8384 13360 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14608 8384 14933 8412
rect 14608 8372 14614 8384
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 16758 8412 16764 8424
rect 16719 8384 16764 8412
rect 14921 8375 14979 8381
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 19337 8415 19395 8421
rect 19337 8412 19349 8415
rect 18555 8384 19349 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 19337 8381 19349 8384
rect 19383 8412 19395 8415
rect 19610 8412 19616 8424
rect 19383 8384 19616 8412
rect 19383 8381 19395 8384
rect 19337 8375 19395 8381
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 21358 8412 21364 8424
rect 20364 8384 21364 8412
rect 11974 8344 11980 8356
rect 11935 8316 11980 8344
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 13722 8344 13728 8356
rect 13372 8316 13728 8344
rect 11238 8276 11244 8288
rect 11199 8248 11244 8276
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 13372 8285 13400 8316
rect 13722 8304 13728 8316
rect 13780 8304 13786 8356
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8344 14427 8347
rect 14642 8344 14648 8356
rect 14415 8316 14648 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 14642 8304 14648 8316
rect 14700 8344 14706 8356
rect 14829 8347 14887 8353
rect 14829 8344 14841 8347
rect 14700 8316 14841 8344
rect 14700 8304 14706 8316
rect 14829 8313 14841 8316
rect 14875 8313 14887 8347
rect 14829 8307 14887 8313
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 16853 8347 16911 8353
rect 16853 8344 16865 8347
rect 16632 8316 16865 8344
rect 16632 8304 16638 8316
rect 16853 8313 16865 8316
rect 16899 8344 16911 8347
rect 17862 8344 17868 8356
rect 16899 8316 17868 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 17862 8304 17868 8316
rect 17920 8304 17926 8356
rect 18782 8344 18788 8356
rect 18743 8316 18788 8344
rect 18782 8304 18788 8316
rect 18840 8344 18846 8356
rect 19429 8347 19487 8353
rect 19429 8344 19441 8347
rect 18840 8316 19441 8344
rect 18840 8304 18846 8316
rect 19429 8313 19441 8316
rect 19475 8344 19487 8347
rect 20364 8344 20392 8384
rect 21358 8372 21364 8384
rect 21416 8372 21422 8424
rect 23661 8415 23719 8421
rect 23661 8381 23673 8415
rect 23707 8412 23719 8415
rect 24026 8412 24032 8424
rect 23707 8384 24032 8412
rect 23707 8381 23719 8384
rect 23661 8375 23719 8381
rect 24026 8372 24032 8384
rect 24084 8372 24090 8424
rect 24673 8415 24731 8421
rect 24673 8381 24685 8415
rect 24719 8412 24731 8415
rect 24762 8412 24768 8424
rect 24719 8384 24768 8412
rect 24719 8381 24731 8384
rect 24673 8375 24731 8381
rect 24762 8372 24768 8384
rect 24820 8412 24826 8424
rect 25501 8415 25559 8421
rect 25501 8412 25513 8415
rect 24820 8384 25513 8412
rect 24820 8372 24826 8384
rect 25501 8381 25513 8384
rect 25547 8381 25559 8415
rect 25501 8375 25559 8381
rect 19475 8316 20392 8344
rect 20441 8347 20499 8353
rect 19475 8313 19487 8316
rect 19429 8307 19487 8313
rect 20441 8313 20453 8347
rect 20487 8344 20499 8347
rect 20898 8344 20904 8356
rect 20487 8316 20904 8344
rect 20487 8313 20499 8316
rect 20441 8307 20499 8313
rect 20898 8304 20904 8316
rect 20956 8304 20962 8356
rect 13357 8279 13415 8285
rect 13357 8245 13369 8279
rect 13403 8245 13415 8279
rect 16298 8276 16304 8288
rect 16259 8248 16304 8276
rect 13357 8239 13415 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 24026 8236 24032 8288
rect 24084 8276 24090 8288
rect 25774 8276 25780 8288
rect 24084 8248 25780 8276
rect 24084 8236 24090 8248
rect 25774 8236 25780 8248
rect 25832 8236 25838 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 11572 8044 11897 8072
rect 11572 8032 11578 8044
rect 11885 8041 11897 8044
rect 11931 8041 11943 8075
rect 11885 8035 11943 8041
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 13446 8072 13452 8084
rect 13035 8044 13452 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13722 8072 13728 8084
rect 13679 8044 13728 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14090 8032 14096 8084
rect 14148 8072 14154 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 14148 8044 14197 8072
rect 14148 8032 14154 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 14734 8072 14740 8084
rect 14695 8044 14740 8072
rect 14185 8035 14243 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8072 16451 8075
rect 16758 8072 16764 8084
rect 16439 8044 16764 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 16758 8032 16764 8044
rect 16816 8072 16822 8084
rect 18969 8075 19027 8081
rect 18969 8072 18981 8075
rect 16816 8044 18981 8072
rect 16816 8032 16822 8044
rect 18969 8041 18981 8044
rect 19015 8041 19027 8075
rect 20622 8072 20628 8084
rect 20583 8044 20628 8072
rect 18969 8035 19027 8041
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 21450 8072 21456 8084
rect 21411 8044 21456 8072
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 22554 8032 22560 8084
rect 22612 8072 22618 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 22612 8044 22937 8072
rect 22612 8032 22618 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 23934 8072 23940 8084
rect 23895 8044 23940 8072
rect 22925 8035 22983 8041
rect 23934 8032 23940 8044
rect 23992 8032 23998 8084
rect 24949 8075 25007 8081
rect 24949 8041 24961 8075
rect 24995 8072 25007 8075
rect 25130 8072 25136 8084
rect 24995 8044 25136 8072
rect 24995 8041 25007 8044
rect 24949 8035 25007 8041
rect 25130 8032 25136 8044
rect 25188 8032 25194 8084
rect 11238 7964 11244 8016
rect 11296 8004 11302 8016
rect 12342 8004 12348 8016
rect 11296 7976 12348 8004
rect 11296 7964 11302 7976
rect 12342 7964 12348 7976
rect 12400 7964 12406 8016
rect 16025 8007 16083 8013
rect 16025 7973 16037 8007
rect 16071 8004 16083 8007
rect 16482 8004 16488 8016
rect 16071 7976 16488 8004
rect 16071 7973 16083 7976
rect 16025 7967 16083 7973
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 19334 8004 19340 8016
rect 19295 7976 19340 8004
rect 19334 7964 19340 7976
rect 19392 7964 19398 8016
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12253 7939 12311 7945
rect 12253 7936 12265 7939
rect 11940 7908 12265 7936
rect 11940 7896 11946 7908
rect 12253 7905 12265 7908
rect 12299 7905 12311 7939
rect 12360 7936 12388 7964
rect 16752 7939 16810 7945
rect 12360 7908 12480 7936
rect 12253 7899 12311 7905
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 12452 7877 12480 7908
rect 16752 7905 16764 7939
rect 16798 7936 16810 7939
rect 17678 7936 17684 7948
rect 16798 7908 17684 7936
rect 16798 7905 16810 7908
rect 16752 7899 16810 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 20901 7939 20959 7945
rect 20901 7905 20913 7939
rect 20947 7936 20959 7939
rect 20990 7936 20996 7948
rect 20947 7908 20996 7936
rect 20947 7905 20959 7908
rect 20901 7899 20959 7905
rect 20990 7896 20996 7908
rect 21048 7896 21054 7948
rect 22741 7939 22799 7945
rect 22741 7905 22753 7939
rect 22787 7936 22799 7939
rect 23198 7936 23204 7948
rect 22787 7908 23204 7936
rect 22787 7905 22799 7908
rect 22741 7899 22799 7905
rect 23198 7896 23204 7908
rect 23256 7896 23262 7948
rect 23658 7896 23664 7948
rect 23716 7936 23722 7948
rect 23753 7939 23811 7945
rect 23753 7936 23765 7939
rect 23716 7908 23765 7936
rect 23716 7896 23722 7908
rect 23753 7905 23765 7908
rect 23799 7905 23811 7939
rect 24762 7936 24768 7948
rect 24723 7908 24768 7936
rect 23753 7899 23811 7905
rect 24762 7896 24768 7908
rect 24820 7896 24826 7948
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 12216 7840 12357 7868
rect 12216 7828 12222 7840
rect 12345 7837 12357 7840
rect 12391 7837 12403 7871
rect 12345 7831 12403 7837
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7837 12495 7871
rect 15470 7868 15476 7880
rect 15431 7840 15476 7868
rect 12437 7831 12495 7837
rect 12360 7800 12388 7831
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 16482 7868 16488 7880
rect 16443 7840 16488 7868
rect 16482 7828 16488 7840
rect 16540 7828 16546 7880
rect 17494 7828 17500 7880
rect 17552 7868 17558 7880
rect 19058 7868 19064 7880
rect 17552 7840 19064 7868
rect 17552 7828 17558 7840
rect 19058 7828 19064 7840
rect 19116 7868 19122 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 19116 7840 19441 7868
rect 19116 7828 19122 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19610 7868 19616 7880
rect 19523 7840 19616 7868
rect 19429 7831 19487 7837
rect 19610 7828 19616 7840
rect 19668 7868 19674 7880
rect 20622 7868 20628 7880
rect 19668 7840 20628 7868
rect 19668 7828 19674 7840
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 12710 7800 12716 7812
rect 12360 7772 12716 7800
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 17865 7803 17923 7809
rect 17865 7800 17877 7803
rect 17828 7772 17877 7800
rect 17828 7760 17834 7772
rect 17865 7769 17877 7772
rect 17911 7769 17923 7803
rect 21082 7800 21088 7812
rect 21043 7772 21088 7800
rect 17865 7763 17923 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 14001 7735 14059 7741
rect 14001 7701 14013 7735
rect 14047 7732 14059 7735
rect 14274 7732 14280 7744
rect 14047 7704 14280 7732
rect 14047 7701 14059 7704
rect 14001 7695 14059 7701
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11296 7500 11529 7528
rect 11296 7488 11302 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 14826 7528 14832 7540
rect 14787 7500 14832 7528
rect 11517 7491 11575 7497
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 15286 7528 15292 7540
rect 15247 7500 15292 7528
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15565 7531 15623 7537
rect 15565 7497 15577 7531
rect 15611 7528 15623 7531
rect 15746 7528 15752 7540
rect 15611 7500 15752 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 16393 7531 16451 7537
rect 16393 7528 16405 7531
rect 16080 7500 16405 7528
rect 16080 7488 16086 7500
rect 16393 7497 16405 7500
rect 16439 7497 16451 7531
rect 16393 7491 16451 7497
rect 17862 7488 17868 7540
rect 17920 7528 17926 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 17920 7500 18061 7528
rect 17920 7488 17926 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 19058 7528 19064 7540
rect 19019 7500 19064 7528
rect 18049 7491 18107 7497
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 19613 7531 19671 7537
rect 19613 7497 19625 7531
rect 19659 7528 19671 7531
rect 19978 7528 19984 7540
rect 19659 7500 19984 7528
rect 19659 7497 19671 7500
rect 19613 7491 19671 7497
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 20622 7528 20628 7540
rect 20583 7500 20628 7528
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 20990 7528 20996 7540
rect 20951 7500 20996 7528
rect 20990 7488 20996 7500
rect 21048 7488 21054 7540
rect 22925 7531 22983 7537
rect 22925 7497 22937 7531
rect 22971 7528 22983 7531
rect 23198 7528 23204 7540
rect 22971 7500 23204 7528
rect 22971 7497 22983 7500
rect 22925 7491 22983 7497
rect 23198 7488 23204 7500
rect 23256 7488 23262 7540
rect 23658 7488 23664 7540
rect 23716 7528 23722 7540
rect 24489 7531 24547 7537
rect 24489 7528 24501 7531
rect 23716 7500 24501 7528
rect 23716 7488 23722 7500
rect 24489 7497 24501 7500
rect 24535 7497 24547 7531
rect 24489 7491 24547 7497
rect 24762 7488 24768 7540
rect 24820 7528 24826 7540
rect 25133 7531 25191 7537
rect 25133 7528 25145 7531
rect 24820 7500 25145 7528
rect 24820 7488 24826 7500
rect 25133 7497 25145 7500
rect 25179 7497 25191 7531
rect 25133 7491 25191 7497
rect 16209 7463 16267 7469
rect 16209 7429 16221 7463
rect 16255 7460 16267 7463
rect 16482 7460 16488 7472
rect 16255 7432 16488 7460
rect 16255 7429 16267 7432
rect 16209 7423 16267 7429
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 23845 7463 23903 7469
rect 23845 7429 23857 7463
rect 23891 7460 23903 7463
rect 24026 7460 24032 7472
rect 23891 7432 24032 7460
rect 23891 7429 23903 7432
rect 23845 7423 23903 7429
rect 24026 7420 24032 7432
rect 24084 7420 24090 7472
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7392 15991 7395
rect 16298 7392 16304 7404
rect 15979 7364 16304 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16298 7352 16304 7364
rect 16356 7392 16362 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16356 7364 16957 7392
rect 16356 7352 16362 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17497 7395 17555 7401
rect 17497 7361 17509 7395
rect 17543 7392 17555 7395
rect 17678 7392 17684 7404
rect 17543 7364 17684 7392
rect 17543 7361 17555 7364
rect 17497 7355 17555 7361
rect 17678 7352 17684 7364
rect 17736 7392 17742 7404
rect 18693 7395 18751 7401
rect 18693 7392 18705 7395
rect 17736 7364 18705 7392
rect 17736 7352 17742 7364
rect 18693 7361 18705 7364
rect 18739 7392 18751 7395
rect 19610 7392 19616 7404
rect 18739 7364 19616 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 19610 7352 19616 7364
rect 19668 7352 19674 7404
rect 20070 7392 20076 7404
rect 20031 7364 20076 7392
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20346 7392 20352 7404
rect 20303 7364 20352 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 21174 7392 21180 7404
rect 21135 7364 21180 7392
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 22370 7392 22376 7404
rect 22331 7364 22376 7392
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 24673 7395 24731 7401
rect 24673 7392 24685 7395
rect 23808 7364 24685 7392
rect 23808 7352 23814 7364
rect 24673 7361 24685 7364
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 12710 7324 12716 7336
rect 12671 7296 12716 7324
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 15381 7327 15439 7333
rect 15381 7324 15393 7327
rect 15344 7296 15393 7324
rect 15344 7284 15350 7296
rect 15381 7293 15393 7296
rect 15427 7293 15439 7327
rect 16758 7324 16764 7336
rect 16719 7296 16764 7324
rect 15381 7287 15439 7293
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 23658 7324 23664 7336
rect 23619 7296 23664 7324
rect 23658 7284 23664 7296
rect 23716 7324 23722 7336
rect 24121 7327 24179 7333
rect 24121 7324 24133 7327
rect 23716 7296 24133 7324
rect 23716 7284 23722 7296
rect 24121 7293 24133 7296
rect 24167 7293 24179 7327
rect 24121 7287 24179 7293
rect 14734 7216 14740 7268
rect 14792 7256 14798 7268
rect 17773 7259 17831 7265
rect 17773 7256 17785 7259
rect 14792 7228 17785 7256
rect 14792 7216 14798 7228
rect 17773 7225 17785 7228
rect 17819 7256 17831 7259
rect 18506 7256 18512 7268
rect 17819 7228 18512 7256
rect 17819 7225 17831 7228
rect 17773 7219 17831 7225
rect 18506 7216 18512 7228
rect 18564 7216 18570 7268
rect 19521 7259 19579 7265
rect 19521 7225 19533 7259
rect 19567 7256 19579 7259
rect 19981 7259 20039 7265
rect 19981 7256 19993 7259
rect 19567 7228 19993 7256
rect 19567 7225 19579 7228
rect 19521 7219 19579 7225
rect 19981 7225 19993 7228
rect 20027 7256 20039 7259
rect 20162 7256 20168 7268
rect 20027 7228 20168 7256
rect 20027 7225 20039 7228
rect 19981 7219 20039 7225
rect 20162 7216 20168 7228
rect 20220 7216 20226 7268
rect 11882 7188 11888 7200
rect 11843 7160 11888 7188
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 16850 7148 16856 7200
rect 16908 7188 16914 7200
rect 16908 7160 16953 7188
rect 16908 7148 16914 7160
rect 18230 7148 18236 7200
rect 18288 7188 18294 7200
rect 18417 7191 18475 7197
rect 18417 7188 18429 7191
rect 18288 7160 18429 7188
rect 18288 7148 18294 7160
rect 18417 7157 18429 7160
rect 18463 7157 18475 7191
rect 18417 7151 18475 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 15470 6944 15476 6996
rect 15528 6984 15534 6996
rect 17494 6984 17500 6996
rect 15528 6956 17500 6984
rect 15528 6944 15534 6956
rect 17494 6944 17500 6956
rect 17552 6944 17558 6996
rect 20073 6987 20131 6993
rect 20073 6953 20085 6987
rect 20119 6984 20131 6987
rect 20346 6984 20352 6996
rect 20119 6956 20352 6984
rect 20119 6953 20131 6956
rect 20073 6947 20131 6953
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 15930 6916 15936 6928
rect 15891 6888 15936 6916
rect 15930 6876 15936 6888
rect 15988 6876 15994 6928
rect 17586 6916 17592 6928
rect 17547 6888 17592 6916
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 16025 6851 16083 6857
rect 16025 6848 16037 6851
rect 15436 6820 16037 6848
rect 15436 6808 15442 6820
rect 16025 6817 16037 6820
rect 16071 6817 16083 6851
rect 16390 6848 16396 6860
rect 16025 6811 16083 6817
rect 16224 6820 16396 6848
rect 16224 6789 16252 6820
rect 16390 6808 16396 6820
rect 16448 6848 16454 6860
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16448 6820 16681 6848
rect 16448 6808 16454 6820
rect 16669 6817 16681 6820
rect 16715 6848 16727 6851
rect 19061 6851 19119 6857
rect 16715 6820 17724 6848
rect 16715 6817 16727 6820
rect 16669 6811 16727 6817
rect 17696 6792 17724 6820
rect 19061 6817 19073 6851
rect 19107 6848 19119 6851
rect 19242 6848 19248 6860
rect 19107 6820 19248 6848
rect 19107 6817 19119 6820
rect 19061 6811 19119 6817
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 19705 6851 19763 6857
rect 19705 6817 19717 6851
rect 19751 6848 19763 6851
rect 20070 6848 20076 6860
rect 19751 6820 20076 6848
rect 19751 6817 19763 6820
rect 19705 6811 19763 6817
rect 20070 6808 20076 6820
rect 20128 6808 20134 6860
rect 23658 6848 23664 6860
rect 23619 6820 23664 6848
rect 23658 6808 23664 6820
rect 23716 6808 23722 6860
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6749 16267 6783
rect 17678 6780 17684 6792
rect 17639 6752 17684 6780
rect 16209 6743 16267 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 15565 6715 15623 6721
rect 15565 6681 15577 6715
rect 15611 6712 15623 6715
rect 16850 6712 16856 6724
rect 15611 6684 16856 6712
rect 15611 6681 15623 6684
rect 15565 6675 15623 6681
rect 16850 6672 16856 6684
rect 16908 6712 16914 6724
rect 16945 6715 17003 6721
rect 16945 6712 16957 6715
rect 16908 6684 16957 6712
rect 16908 6672 16914 6684
rect 16945 6681 16957 6684
rect 16991 6681 17003 6715
rect 16945 6675 17003 6681
rect 23845 6715 23903 6721
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 25866 6712 25872 6724
rect 23891 6684 25872 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 25866 6672 25872 6684
rect 25924 6672 25930 6724
rect 16666 6604 16672 6656
rect 16724 6644 16730 6656
rect 17129 6647 17187 6653
rect 17129 6644 17141 6647
rect 16724 6616 17141 6644
rect 16724 6604 16730 6616
rect 17129 6613 17141 6616
rect 17175 6613 17187 6647
rect 18230 6644 18236 6656
rect 18191 6616 18236 6644
rect 17129 6607 17187 6613
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15436 6412 15577 6440
rect 15436 6400 15442 6412
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15930 6440 15936 6452
rect 15891 6412 15936 6440
rect 15565 6403 15623 6409
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16390 6440 16396 6452
rect 16351 6412 16396 6440
rect 16390 6400 16396 6412
rect 16448 6440 16454 6452
rect 16761 6443 16819 6449
rect 16761 6440 16773 6443
rect 16448 6412 16773 6440
rect 16448 6400 16454 6412
rect 16761 6409 16773 6412
rect 16807 6409 16819 6443
rect 17494 6440 17500 6452
rect 17455 6412 17500 6440
rect 16761 6403 16819 6409
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 23658 6400 23664 6452
rect 23716 6440 23722 6452
rect 23845 6443 23903 6449
rect 23845 6440 23857 6443
rect 23716 6412 23857 6440
rect 23716 6400 23722 6412
rect 23845 6409 23857 6412
rect 23891 6409 23903 6443
rect 23845 6403 23903 6409
rect 17126 6100 17132 6112
rect 17087 6072 17132 6100
rect 17126 6060 17132 6072
rect 17184 6100 17190 6112
rect 17586 6100 17592 6112
rect 17184 6072 17592 6100
rect 17184 6060 17190 6072
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 12483 2536 13124 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 13096 2496 13124 2536
rect 13164 2499 13222 2505
rect 13164 2496 13176 2499
rect 13096 2468 13176 2496
rect 13164 2465 13176 2468
rect 13210 2496 13222 2499
rect 13722 2496 13728 2508
rect 13210 2468 13728 2496
rect 13210 2465 13222 2468
rect 13164 2459 13222 2465
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2428 12038 2440
rect 12894 2428 12900 2440
rect 12032 2400 12900 2428
rect 12032 2388 12038 2400
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 13452 27004 13504 27056
rect 15384 27004 15436 27056
rect 10048 26188 10100 26240
rect 14832 26188 14884 26240
rect 11612 26120 11664 26172
rect 19984 26120 20036 26172
rect 12072 26052 12124 26104
rect 9588 25984 9640 26036
rect 18144 25984 18196 26036
rect 2688 25916 2740 25968
rect 17500 25916 17552 25968
rect 2228 25848 2280 25900
rect 6276 25848 6328 25900
rect 10968 25848 11020 25900
rect 20904 25848 20956 25900
rect 3792 25780 3844 25832
rect 6460 25780 6512 25832
rect 8668 25780 8720 25832
rect 11980 25780 12032 25832
rect 12808 25780 12860 25832
rect 22652 25780 22704 25832
rect 1952 25712 2004 25764
rect 3148 25644 3200 25696
rect 12440 25644 12492 25696
rect 19064 25712 19116 25764
rect 17224 25644 17276 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 1952 25483 2004 25492
rect 1952 25449 1961 25483
rect 1961 25449 1995 25483
rect 1995 25449 2004 25483
rect 1952 25440 2004 25449
rect 3608 25440 3660 25492
rect 4804 25483 4856 25492
rect 4804 25449 4813 25483
rect 4813 25449 4847 25483
rect 4847 25449 4856 25483
rect 4804 25440 4856 25449
rect 3056 25372 3108 25424
rect 7288 25440 7340 25492
rect 10968 25483 11020 25492
rect 10968 25449 10977 25483
rect 10977 25449 11011 25483
rect 11011 25449 11020 25483
rect 10968 25440 11020 25449
rect 12072 25483 12124 25492
rect 12072 25449 12081 25483
rect 12081 25449 12115 25483
rect 12115 25449 12124 25483
rect 12072 25440 12124 25449
rect 17776 25440 17828 25492
rect 20076 25440 20128 25492
rect 21824 25440 21876 25492
rect 22652 25483 22704 25492
rect 22652 25449 22661 25483
rect 22661 25449 22695 25483
rect 22695 25449 22704 25483
rect 22652 25440 22704 25449
rect 23756 25483 23808 25492
rect 11704 25372 11756 25424
rect 2504 25304 2556 25356
rect 2780 25347 2832 25356
rect 2780 25313 2789 25347
rect 2789 25313 2823 25347
rect 2823 25313 2832 25347
rect 2780 25304 2832 25313
rect 5448 25304 5500 25356
rect 6552 25304 6604 25356
rect 8484 25347 8536 25356
rect 8484 25313 8493 25347
rect 8493 25313 8527 25347
rect 8527 25313 8536 25347
rect 8484 25304 8536 25313
rect 9588 25304 9640 25356
rect 2964 25279 3016 25288
rect 2964 25245 2973 25279
rect 2973 25245 3007 25279
rect 3007 25245 3016 25279
rect 2964 25236 3016 25245
rect 8300 25236 8352 25288
rect 8760 25279 8812 25288
rect 8760 25245 8769 25279
rect 8769 25245 8803 25279
rect 8803 25245 8812 25279
rect 8760 25236 8812 25245
rect 1952 25100 2004 25152
rect 2504 25100 2556 25152
rect 3424 25143 3476 25152
rect 3424 25109 3433 25143
rect 3433 25109 3467 25143
rect 3467 25109 3476 25143
rect 3424 25100 3476 25109
rect 3700 25100 3752 25152
rect 5172 25168 5224 25220
rect 5908 25168 5960 25220
rect 8024 25168 8076 25220
rect 10416 25168 10468 25220
rect 5540 25100 5592 25152
rect 6644 25100 6696 25152
rect 7012 25100 7064 25152
rect 7656 25100 7708 25152
rect 8944 25100 8996 25152
rect 10692 25236 10744 25288
rect 11520 25279 11572 25288
rect 11520 25245 11529 25279
rect 11529 25245 11563 25279
rect 11563 25245 11572 25279
rect 11520 25236 11572 25245
rect 11980 25100 12032 25152
rect 13268 25372 13320 25424
rect 12808 25304 12860 25356
rect 14464 25304 14516 25356
rect 15476 25372 15528 25424
rect 16948 25372 17000 25424
rect 17684 25304 17736 25356
rect 18328 25347 18380 25356
rect 18328 25313 18337 25347
rect 18337 25313 18371 25347
rect 18371 25313 18380 25347
rect 18328 25304 18380 25313
rect 19984 25347 20036 25356
rect 19984 25313 19993 25347
rect 19993 25313 20027 25347
rect 20027 25313 20036 25347
rect 19984 25304 20036 25313
rect 23756 25449 23765 25483
rect 23765 25449 23799 25483
rect 23799 25449 23808 25483
rect 23756 25440 23808 25449
rect 25872 25440 25924 25492
rect 25320 25372 25372 25424
rect 23848 25304 23900 25356
rect 25136 25347 25188 25356
rect 25136 25313 25145 25347
rect 25145 25313 25179 25347
rect 25179 25313 25188 25347
rect 25136 25304 25188 25313
rect 12900 25236 12952 25288
rect 13176 25236 13228 25288
rect 15936 25279 15988 25288
rect 15292 25168 15344 25220
rect 15936 25245 15945 25279
rect 15945 25245 15979 25279
rect 15979 25245 15988 25279
rect 15936 25236 15988 25245
rect 16120 25279 16172 25288
rect 16120 25245 16129 25279
rect 16129 25245 16163 25279
rect 16163 25245 16172 25279
rect 16120 25236 16172 25245
rect 19524 25168 19576 25220
rect 24768 25168 24820 25220
rect 16580 25143 16632 25152
rect 16580 25109 16589 25143
rect 16589 25109 16623 25143
rect 16623 25109 16632 25143
rect 16580 25100 16632 25109
rect 18052 25143 18104 25152
rect 18052 25109 18061 25143
rect 18061 25109 18095 25143
rect 18095 25109 18104 25143
rect 18052 25100 18104 25109
rect 22928 25100 22980 25152
rect 24676 25100 24728 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 1584 24896 1636 24948
rect 18328 24896 18380 24948
rect 18880 24939 18932 24948
rect 18880 24905 18889 24939
rect 18889 24905 18923 24939
rect 18923 24905 18932 24939
rect 18880 24896 18932 24905
rect 1492 24828 1544 24880
rect 2504 24828 2556 24880
rect 2780 24828 2832 24880
rect 4804 24828 4856 24880
rect 5448 24871 5500 24880
rect 5448 24837 5457 24871
rect 5457 24837 5491 24871
rect 5491 24837 5500 24871
rect 5448 24828 5500 24837
rect 10692 24871 10744 24880
rect 10692 24837 10701 24871
rect 10701 24837 10735 24871
rect 10735 24837 10744 24871
rect 10692 24828 10744 24837
rect 11612 24828 11664 24880
rect 12900 24828 12952 24880
rect 16120 24871 16172 24880
rect 2044 24803 2096 24812
rect 2044 24769 2053 24803
rect 2053 24769 2087 24803
rect 2087 24769 2096 24803
rect 2044 24760 2096 24769
rect 2228 24803 2280 24812
rect 2228 24769 2237 24803
rect 2237 24769 2271 24803
rect 2271 24769 2280 24803
rect 2228 24760 2280 24769
rect 7472 24803 7524 24812
rect 7472 24769 7481 24803
rect 7481 24769 7515 24803
rect 7515 24769 7524 24803
rect 7472 24760 7524 24769
rect 13176 24760 13228 24812
rect 16120 24837 16129 24871
rect 16129 24837 16163 24871
rect 16163 24837 16172 24871
rect 16120 24828 16172 24837
rect 16856 24828 16908 24880
rect 25136 24828 25188 24880
rect 1952 24735 2004 24744
rect 1952 24701 1961 24735
rect 1961 24701 1995 24735
rect 1995 24701 2004 24735
rect 1952 24692 2004 24701
rect 3240 24692 3292 24744
rect 3424 24735 3476 24744
rect 3424 24701 3458 24735
rect 3458 24701 3476 24735
rect 3424 24692 3476 24701
rect 5540 24692 5592 24744
rect 7288 24692 7340 24744
rect 8576 24735 8628 24744
rect 8576 24701 8585 24735
rect 8585 24701 8619 24735
rect 8619 24701 8628 24735
rect 8576 24692 8628 24701
rect 12072 24692 12124 24744
rect 12992 24692 13044 24744
rect 13452 24735 13504 24744
rect 13452 24701 13461 24735
rect 13461 24701 13495 24735
rect 13495 24701 13504 24735
rect 13452 24692 13504 24701
rect 2872 24624 2924 24676
rect 6092 24624 6144 24676
rect 7932 24624 7984 24676
rect 8760 24624 8812 24676
rect 9864 24624 9916 24676
rect 14372 24624 14424 24676
rect 15200 24760 15252 24812
rect 18328 24760 18380 24812
rect 20996 24760 21048 24812
rect 21548 24803 21600 24812
rect 21548 24769 21557 24803
rect 21557 24769 21591 24803
rect 21591 24769 21600 24803
rect 21548 24760 21600 24769
rect 16580 24735 16632 24744
rect 14556 24624 14608 24676
rect 15384 24667 15436 24676
rect 1860 24556 1912 24608
rect 1952 24556 2004 24608
rect 2780 24556 2832 24608
rect 3608 24556 3660 24608
rect 3884 24556 3936 24608
rect 6000 24556 6052 24608
rect 6552 24599 6604 24608
rect 6552 24565 6561 24599
rect 6561 24565 6595 24599
rect 6595 24565 6604 24599
rect 6552 24556 6604 24565
rect 7196 24556 7248 24608
rect 7288 24599 7340 24608
rect 7288 24565 7297 24599
rect 7297 24565 7331 24599
rect 7331 24565 7340 24599
rect 8116 24599 8168 24608
rect 7288 24556 7340 24565
rect 8116 24565 8125 24599
rect 8125 24565 8159 24599
rect 8159 24565 8168 24599
rect 8116 24556 8168 24565
rect 9956 24599 10008 24608
rect 9956 24565 9965 24599
rect 9965 24565 9999 24599
rect 9999 24565 10008 24599
rect 9956 24556 10008 24565
rect 11428 24556 11480 24608
rect 12808 24556 12860 24608
rect 13360 24599 13412 24608
rect 13360 24565 13369 24599
rect 13369 24565 13403 24599
rect 13403 24565 13412 24599
rect 13360 24556 13412 24565
rect 14004 24599 14056 24608
rect 14004 24565 14013 24599
rect 14013 24565 14047 24599
rect 14047 24565 14056 24599
rect 14004 24556 14056 24565
rect 15384 24633 15393 24667
rect 15393 24633 15427 24667
rect 15427 24633 15436 24667
rect 15384 24624 15436 24633
rect 16580 24701 16589 24735
rect 16589 24701 16623 24735
rect 16623 24701 16632 24735
rect 16580 24692 16632 24701
rect 16948 24692 17000 24744
rect 18052 24735 18104 24744
rect 18052 24701 18061 24735
rect 18061 24701 18095 24735
rect 18095 24701 18104 24735
rect 18052 24692 18104 24701
rect 18880 24692 18932 24744
rect 15476 24599 15528 24608
rect 15476 24565 15485 24599
rect 15485 24565 15519 24599
rect 15519 24565 15528 24599
rect 15476 24556 15528 24565
rect 15936 24556 15988 24608
rect 16764 24599 16816 24608
rect 16764 24565 16773 24599
rect 16773 24565 16807 24599
rect 16807 24565 16816 24599
rect 16764 24556 16816 24565
rect 17684 24556 17736 24608
rect 19248 24599 19300 24608
rect 19248 24565 19257 24599
rect 19257 24565 19291 24599
rect 19291 24565 19300 24599
rect 19248 24556 19300 24565
rect 19524 24556 19576 24608
rect 20812 24624 20864 24676
rect 20168 24599 20220 24608
rect 20168 24565 20177 24599
rect 20177 24565 20211 24599
rect 20211 24565 20220 24599
rect 20168 24556 20220 24565
rect 20536 24599 20588 24608
rect 20536 24565 20545 24599
rect 20545 24565 20579 24599
rect 20579 24565 20588 24599
rect 20536 24556 20588 24565
rect 21916 24556 21968 24608
rect 22928 24760 22980 24812
rect 23480 24803 23532 24812
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 24308 24803 24360 24812
rect 23480 24760 23532 24769
rect 24308 24769 24317 24803
rect 24317 24769 24351 24803
rect 24351 24769 24360 24803
rect 24308 24760 24360 24769
rect 23756 24692 23808 24744
rect 24124 24692 24176 24744
rect 25780 24692 25832 24744
rect 22652 24624 22704 24676
rect 23204 24624 23256 24676
rect 23848 24624 23900 24676
rect 22468 24599 22520 24608
rect 22468 24565 22477 24599
rect 22477 24565 22511 24599
rect 22511 24565 22520 24599
rect 22468 24556 22520 24565
rect 22928 24556 22980 24608
rect 23756 24556 23808 24608
rect 24216 24556 24268 24608
rect 25412 24599 25464 24608
rect 25412 24565 25421 24599
rect 25421 24565 25455 24599
rect 25455 24565 25464 24599
rect 25412 24556 25464 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 2044 24352 2096 24404
rect 2320 24395 2372 24404
rect 2320 24361 2329 24395
rect 2329 24361 2363 24395
rect 2363 24361 2372 24395
rect 2320 24352 2372 24361
rect 2872 24395 2924 24404
rect 2872 24361 2881 24395
rect 2881 24361 2915 24395
rect 2915 24361 2924 24395
rect 2872 24352 2924 24361
rect 3240 24352 3292 24404
rect 3884 24395 3936 24404
rect 3884 24361 3893 24395
rect 3893 24361 3927 24395
rect 3927 24361 3936 24395
rect 3884 24352 3936 24361
rect 4436 24395 4488 24404
rect 4436 24361 4445 24395
rect 4445 24361 4479 24395
rect 4479 24361 4488 24395
rect 4436 24352 4488 24361
rect 2136 24284 2188 24336
rect 7012 24352 7064 24404
rect 8484 24352 8536 24404
rect 9956 24352 10008 24404
rect 10692 24395 10744 24404
rect 10692 24361 10701 24395
rect 10701 24361 10735 24395
rect 10735 24361 10744 24395
rect 10692 24352 10744 24361
rect 11152 24395 11204 24404
rect 11152 24361 11161 24395
rect 11161 24361 11195 24395
rect 11195 24361 11204 24395
rect 11152 24352 11204 24361
rect 11704 24395 11756 24404
rect 11704 24361 11713 24395
rect 11713 24361 11747 24395
rect 11747 24361 11756 24395
rect 11704 24352 11756 24361
rect 13452 24352 13504 24404
rect 16856 24352 16908 24404
rect 17040 24395 17092 24404
rect 17040 24361 17049 24395
rect 17049 24361 17083 24395
rect 17083 24361 17092 24395
rect 17040 24352 17092 24361
rect 17224 24395 17276 24404
rect 17224 24361 17233 24395
rect 17233 24361 17267 24395
rect 17267 24361 17276 24395
rect 17224 24352 17276 24361
rect 18144 24352 18196 24404
rect 20536 24352 20588 24404
rect 23112 24352 23164 24404
rect 23940 24352 23992 24404
rect 25228 24395 25280 24404
rect 25228 24361 25237 24395
rect 25237 24361 25271 24395
rect 25271 24361 25280 24395
rect 25228 24352 25280 24361
rect 25504 24352 25556 24404
rect 2044 24216 2096 24268
rect 2320 24216 2372 24268
rect 2596 24216 2648 24268
rect 3332 24216 3384 24268
rect 4528 24259 4580 24268
rect 4528 24225 4537 24259
rect 4537 24225 4571 24259
rect 4571 24225 4580 24259
rect 4528 24216 4580 24225
rect 6092 24284 6144 24336
rect 8576 24284 8628 24336
rect 9588 24284 9640 24336
rect 10968 24284 11020 24336
rect 11244 24284 11296 24336
rect 12072 24284 12124 24336
rect 4620 24191 4672 24200
rect 4620 24157 4629 24191
rect 4629 24157 4663 24191
rect 4663 24157 4672 24191
rect 4620 24148 4672 24157
rect 5172 24191 5224 24200
rect 5172 24157 5181 24191
rect 5181 24157 5215 24191
rect 5215 24157 5224 24191
rect 6368 24216 6420 24268
rect 8208 24216 8260 24268
rect 12716 24259 12768 24268
rect 12716 24225 12725 24259
rect 12725 24225 12759 24259
rect 12759 24225 12768 24259
rect 12716 24216 12768 24225
rect 14648 24216 14700 24268
rect 15292 24216 15344 24268
rect 17592 24259 17644 24268
rect 17592 24225 17601 24259
rect 17601 24225 17635 24259
rect 17635 24225 17644 24259
rect 17592 24216 17644 24225
rect 5172 24148 5224 24157
rect 9312 24148 9364 24200
rect 11704 24148 11756 24200
rect 12808 24191 12860 24200
rect 12808 24157 12817 24191
rect 12817 24157 12851 24191
rect 12851 24157 12860 24191
rect 12808 24148 12860 24157
rect 14740 24148 14792 24200
rect 16304 24191 16356 24200
rect 16304 24157 16313 24191
rect 16313 24157 16347 24191
rect 16347 24157 16356 24191
rect 16304 24148 16356 24157
rect 20168 24284 20220 24336
rect 20352 24216 20404 24268
rect 21824 24216 21876 24268
rect 22836 24216 22888 24268
rect 3516 24080 3568 24132
rect 7932 24123 7984 24132
rect 7932 24089 7941 24123
rect 7941 24089 7975 24123
rect 7975 24089 7984 24123
rect 7932 24080 7984 24089
rect 14280 24123 14332 24132
rect 14280 24089 14289 24123
rect 14289 24089 14323 24123
rect 14323 24089 14332 24123
rect 14280 24080 14332 24089
rect 2412 24055 2464 24064
rect 2412 24021 2421 24055
rect 2421 24021 2455 24055
rect 2455 24021 2464 24055
rect 2412 24012 2464 24021
rect 4068 24055 4120 24064
rect 4068 24021 4077 24055
rect 4077 24021 4111 24055
rect 4111 24021 4120 24055
rect 4068 24012 4120 24021
rect 5540 24055 5592 24064
rect 5540 24021 5549 24055
rect 5549 24021 5583 24055
rect 5583 24021 5592 24055
rect 5540 24012 5592 24021
rect 6920 24012 6972 24064
rect 7104 24012 7156 24064
rect 7472 24012 7524 24064
rect 8300 24055 8352 24064
rect 8300 24021 8309 24055
rect 8309 24021 8343 24055
rect 8343 24021 8352 24055
rect 8300 24012 8352 24021
rect 9496 24055 9548 24064
rect 9496 24021 9505 24055
rect 9505 24021 9539 24055
rect 9539 24021 9548 24055
rect 9496 24012 9548 24021
rect 12256 24055 12308 24064
rect 12256 24021 12265 24055
rect 12265 24021 12299 24055
rect 12299 24021 12308 24055
rect 12256 24012 12308 24021
rect 12992 24012 13044 24064
rect 13912 24012 13964 24064
rect 15384 24080 15436 24132
rect 15752 24080 15804 24132
rect 19340 24148 19392 24200
rect 17868 24080 17920 24132
rect 18788 24080 18840 24132
rect 19984 24148 20036 24200
rect 21732 24148 21784 24200
rect 22928 24148 22980 24200
rect 24216 24148 24268 24200
rect 25688 24148 25740 24200
rect 21824 24080 21876 24132
rect 23388 24080 23440 24132
rect 14464 24012 14516 24064
rect 16212 24012 16264 24064
rect 22008 24012 22060 24064
rect 23296 24055 23348 24064
rect 23296 24021 23305 24055
rect 23305 24021 23339 24055
rect 23339 24021 23348 24055
rect 23296 24012 23348 24021
rect 24860 24055 24912 24064
rect 24860 24021 24869 24055
rect 24869 24021 24903 24055
rect 24903 24021 24912 24055
rect 24860 24012 24912 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2688 23808 2740 23860
rect 3332 23808 3384 23860
rect 4620 23808 4672 23860
rect 5356 23851 5408 23860
rect 5356 23817 5365 23851
rect 5365 23817 5399 23851
rect 5399 23817 5408 23851
rect 5356 23808 5408 23817
rect 9312 23851 9364 23860
rect 9312 23817 9321 23851
rect 9321 23817 9355 23851
rect 9355 23817 9364 23851
rect 9312 23808 9364 23817
rect 9588 23851 9640 23860
rect 9588 23817 9597 23851
rect 9597 23817 9631 23851
rect 9631 23817 9640 23851
rect 9588 23808 9640 23817
rect 12072 23808 12124 23860
rect 12716 23851 12768 23860
rect 12716 23817 12725 23851
rect 12725 23817 12759 23851
rect 12759 23817 12768 23851
rect 12716 23808 12768 23817
rect 14740 23808 14792 23860
rect 19524 23808 19576 23860
rect 19892 23851 19944 23860
rect 19892 23817 19901 23851
rect 19901 23817 19935 23851
rect 19935 23817 19944 23851
rect 19892 23808 19944 23817
rect 25412 23851 25464 23860
rect 25412 23817 25421 23851
rect 25421 23817 25455 23851
rect 25455 23817 25464 23851
rect 25412 23808 25464 23817
rect 25688 23808 25740 23860
rect 2872 23740 2924 23792
rect 1860 23672 1912 23724
rect 2504 23672 2556 23724
rect 3516 23740 3568 23792
rect 6368 23783 6420 23792
rect 6368 23749 6377 23783
rect 6377 23749 6411 23783
rect 6411 23749 6420 23783
rect 6368 23740 6420 23749
rect 9128 23740 9180 23792
rect 3240 23672 3292 23724
rect 8852 23715 8904 23724
rect 8852 23681 8861 23715
rect 8861 23681 8895 23715
rect 8895 23681 8904 23715
rect 8852 23672 8904 23681
rect 16856 23783 16908 23792
rect 16856 23749 16865 23783
rect 16865 23749 16899 23783
rect 16899 23749 16908 23783
rect 16856 23740 16908 23749
rect 20352 23783 20404 23792
rect 20352 23749 20361 23783
rect 20361 23749 20395 23783
rect 20395 23749 20404 23783
rect 20352 23740 20404 23749
rect 24952 23783 25004 23792
rect 24952 23749 24961 23783
rect 24961 23749 24995 23783
rect 24995 23749 25004 23783
rect 24952 23740 25004 23749
rect 25504 23740 25556 23792
rect 2136 23604 2188 23656
rect 1308 23536 1360 23588
rect 3608 23604 3660 23656
rect 2688 23468 2740 23520
rect 3884 23536 3936 23588
rect 6552 23536 6604 23588
rect 5632 23468 5684 23520
rect 6092 23468 6144 23520
rect 7012 23511 7064 23520
rect 7012 23477 7021 23511
rect 7021 23477 7055 23511
rect 7055 23477 7064 23511
rect 7012 23468 7064 23477
rect 8208 23604 8260 23656
rect 9312 23604 9364 23656
rect 15384 23672 15436 23724
rect 18788 23715 18840 23724
rect 18788 23681 18797 23715
rect 18797 23681 18831 23715
rect 18831 23681 18840 23715
rect 18788 23672 18840 23681
rect 24216 23715 24268 23724
rect 24216 23681 24225 23715
rect 24225 23681 24259 23715
rect 24259 23681 24268 23715
rect 24216 23672 24268 23681
rect 11520 23604 11572 23656
rect 12992 23647 13044 23656
rect 12992 23613 13001 23647
rect 13001 23613 13035 23647
rect 13035 23613 13044 23647
rect 12992 23604 13044 23613
rect 9956 23536 10008 23588
rect 17592 23604 17644 23656
rect 18144 23604 18196 23656
rect 19432 23604 19484 23656
rect 13544 23536 13596 23588
rect 14096 23536 14148 23588
rect 15292 23579 15344 23588
rect 15292 23545 15301 23579
rect 15301 23545 15335 23579
rect 15335 23545 15344 23579
rect 15292 23536 15344 23545
rect 15752 23579 15804 23588
rect 15752 23545 15786 23579
rect 15786 23545 15804 23579
rect 17776 23579 17828 23588
rect 15752 23536 15804 23545
rect 17776 23545 17785 23579
rect 17785 23545 17819 23579
rect 17819 23545 17828 23579
rect 17776 23536 17828 23545
rect 7932 23468 7984 23520
rect 8116 23468 8168 23520
rect 8668 23511 8720 23520
rect 8668 23477 8677 23511
rect 8677 23477 8711 23511
rect 8711 23477 8720 23511
rect 8668 23468 8720 23477
rect 9772 23468 9824 23520
rect 10784 23468 10836 23520
rect 11060 23468 11112 23520
rect 11796 23511 11848 23520
rect 11796 23477 11805 23511
rect 11805 23477 11839 23511
rect 11839 23477 11848 23511
rect 11796 23468 11848 23477
rect 14004 23468 14056 23520
rect 19340 23511 19392 23520
rect 19340 23477 19349 23511
rect 19349 23477 19383 23511
rect 19383 23477 19392 23511
rect 19340 23468 19392 23477
rect 20996 23604 21048 23656
rect 25688 23604 25740 23656
rect 21456 23468 21508 23520
rect 21732 23468 21784 23520
rect 22836 23468 22888 23520
rect 23572 23468 23624 23520
rect 23940 23468 23992 23520
rect 24124 23511 24176 23520
rect 24124 23477 24133 23511
rect 24133 23477 24167 23511
rect 24167 23477 24176 23511
rect 24124 23468 24176 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2780 23264 2832 23316
rect 1400 23196 1452 23248
rect 1768 23196 1820 23248
rect 3240 23264 3292 23316
rect 3516 23239 3568 23248
rect 3516 23205 3525 23239
rect 3525 23205 3559 23239
rect 3559 23205 3568 23239
rect 3516 23196 3568 23205
rect 1584 23060 1636 23112
rect 3240 23128 3292 23180
rect 4436 23264 4488 23316
rect 8116 23264 8168 23316
rect 8668 23264 8720 23316
rect 10968 23264 11020 23316
rect 11152 23307 11204 23316
rect 11152 23273 11161 23307
rect 11161 23273 11195 23307
rect 11195 23273 11204 23307
rect 11152 23264 11204 23273
rect 12900 23307 12952 23316
rect 12900 23273 12909 23307
rect 12909 23273 12943 23307
rect 12943 23273 12952 23307
rect 12900 23264 12952 23273
rect 13176 23264 13228 23316
rect 18788 23264 18840 23316
rect 20996 23264 21048 23316
rect 23388 23264 23440 23316
rect 24768 23264 24820 23316
rect 24952 23307 25004 23316
rect 24952 23273 24961 23307
rect 24961 23273 24995 23307
rect 24995 23273 25004 23307
rect 24952 23264 25004 23273
rect 25228 23264 25280 23316
rect 5632 23196 5684 23248
rect 7840 23239 7892 23248
rect 7840 23205 7849 23239
rect 7849 23205 7883 23239
rect 7883 23205 7892 23239
rect 7840 23196 7892 23205
rect 8852 23196 8904 23248
rect 9404 23196 9456 23248
rect 9956 23196 10008 23248
rect 4988 23128 5040 23180
rect 5448 23128 5500 23180
rect 6920 23171 6972 23180
rect 6920 23137 6929 23171
rect 6929 23137 6963 23171
rect 6963 23137 6972 23171
rect 6920 23128 6972 23137
rect 10048 23171 10100 23180
rect 10048 23137 10057 23171
rect 10057 23137 10091 23171
rect 10091 23137 10100 23171
rect 10048 23128 10100 23137
rect 3056 23103 3108 23112
rect 1676 22992 1728 23044
rect 3056 23069 3065 23103
rect 3065 23069 3099 23103
rect 3099 23069 3108 23103
rect 3056 23060 3108 23069
rect 3424 23060 3476 23112
rect 6552 23060 6604 23112
rect 8116 23060 8168 23112
rect 8760 23060 8812 23112
rect 8944 23060 8996 23112
rect 11980 23196 12032 23248
rect 11520 23171 11572 23180
rect 11520 23137 11529 23171
rect 11529 23137 11563 23171
rect 11563 23137 11572 23171
rect 11520 23128 11572 23137
rect 11796 23171 11848 23180
rect 11796 23137 11830 23171
rect 11830 23137 11848 23171
rect 11796 23128 11848 23137
rect 14740 23128 14792 23180
rect 16396 23196 16448 23248
rect 17960 23239 18012 23248
rect 17960 23205 17969 23239
rect 17969 23205 18003 23239
rect 18003 23205 18012 23239
rect 17960 23196 18012 23205
rect 18328 23196 18380 23248
rect 24400 23239 24452 23248
rect 16856 23128 16908 23180
rect 19524 23128 19576 23180
rect 24400 23205 24409 23239
rect 24409 23205 24443 23239
rect 24443 23205 24452 23239
rect 24400 23196 24452 23205
rect 25044 23196 25096 23248
rect 21732 23171 21784 23180
rect 21732 23137 21766 23171
rect 21766 23137 21784 23171
rect 21732 23128 21784 23137
rect 12992 23060 13044 23112
rect 15384 23060 15436 23112
rect 16028 23103 16080 23112
rect 16028 23069 16037 23103
rect 16037 23069 16071 23103
rect 16071 23069 16080 23103
rect 16028 23060 16080 23069
rect 19708 23103 19760 23112
rect 19708 23069 19717 23103
rect 19717 23069 19751 23103
rect 19751 23069 19760 23103
rect 19708 23060 19760 23069
rect 19892 23103 19944 23112
rect 19892 23069 19901 23103
rect 19901 23069 19935 23103
rect 19935 23069 19944 23103
rect 19892 23060 19944 23069
rect 21456 23103 21508 23112
rect 21456 23069 21465 23103
rect 21465 23069 21499 23103
rect 21499 23069 21508 23103
rect 21456 23060 21508 23069
rect 24216 23060 24268 23112
rect 1952 22967 2004 22976
rect 1952 22933 1961 22967
rect 1961 22933 1995 22967
rect 1995 22933 2004 22967
rect 1952 22924 2004 22933
rect 2320 22967 2372 22976
rect 2320 22933 2329 22967
rect 2329 22933 2363 22967
rect 2363 22933 2372 22967
rect 2320 22924 2372 22933
rect 2596 22924 2648 22976
rect 3700 22992 3752 23044
rect 8024 23035 8076 23044
rect 8024 23001 8033 23035
rect 8033 23001 8067 23035
rect 8067 23001 8076 23035
rect 8024 22992 8076 23001
rect 13544 23035 13596 23044
rect 13544 23001 13553 23035
rect 13553 23001 13587 23035
rect 13587 23001 13596 23035
rect 13544 22992 13596 23001
rect 14832 22992 14884 23044
rect 17408 23035 17460 23044
rect 17408 23001 17417 23035
rect 17417 23001 17451 23035
rect 17451 23001 17460 23035
rect 17408 22992 17460 23001
rect 18972 22992 19024 23044
rect 19432 22992 19484 23044
rect 4528 22924 4580 22976
rect 6368 22924 6420 22976
rect 7104 22924 7156 22976
rect 13820 22967 13872 22976
rect 13820 22933 13829 22967
rect 13829 22933 13863 22967
rect 13863 22933 13872 22967
rect 13820 22924 13872 22933
rect 14004 22924 14056 22976
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 16304 22924 16356 22976
rect 19248 22967 19300 22976
rect 19248 22933 19257 22967
rect 19257 22933 19291 22967
rect 19291 22933 19300 22967
rect 19248 22924 19300 22933
rect 20720 22967 20772 22976
rect 20720 22933 20729 22967
rect 20729 22933 20763 22967
rect 20763 22933 20772 22967
rect 20720 22924 20772 22933
rect 22560 22924 22612 22976
rect 23020 22924 23072 22976
rect 24124 22924 24176 22976
rect 25136 22924 25188 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2320 22584 2372 22636
rect 3516 22720 3568 22772
rect 4988 22763 5040 22772
rect 4988 22729 4997 22763
rect 4997 22729 5031 22763
rect 5031 22729 5040 22763
rect 4988 22720 5040 22729
rect 4620 22652 4672 22704
rect 3884 22627 3936 22636
rect 3884 22593 3893 22627
rect 3893 22593 3927 22627
rect 3927 22593 3936 22627
rect 3884 22584 3936 22593
rect 4804 22584 4856 22636
rect 4988 22584 5040 22636
rect 1952 22516 2004 22568
rect 1400 22380 1452 22432
rect 2596 22448 2648 22500
rect 1768 22423 1820 22432
rect 1768 22389 1777 22423
rect 1777 22389 1811 22423
rect 1811 22389 1820 22423
rect 1768 22380 1820 22389
rect 2504 22380 2556 22432
rect 5540 22720 5592 22772
rect 7472 22763 7524 22772
rect 7472 22729 7481 22763
rect 7481 22729 7515 22763
rect 7515 22729 7524 22763
rect 7472 22720 7524 22729
rect 8760 22720 8812 22772
rect 9128 22720 9180 22772
rect 11520 22763 11572 22772
rect 11520 22729 11529 22763
rect 11529 22729 11563 22763
rect 11563 22729 11572 22763
rect 11520 22720 11572 22729
rect 14648 22720 14700 22772
rect 15292 22763 15344 22772
rect 15292 22729 15301 22763
rect 15301 22729 15335 22763
rect 15335 22729 15344 22763
rect 15292 22720 15344 22729
rect 16028 22763 16080 22772
rect 16028 22729 16037 22763
rect 16037 22729 16071 22763
rect 16071 22729 16080 22763
rect 16028 22720 16080 22729
rect 17500 22720 17552 22772
rect 18512 22763 18564 22772
rect 5356 22584 5408 22636
rect 6828 22652 6880 22704
rect 9680 22652 9732 22704
rect 10048 22652 10100 22704
rect 12992 22652 13044 22704
rect 10968 22627 11020 22636
rect 10968 22593 10977 22627
rect 10977 22593 11011 22627
rect 11011 22593 11020 22627
rect 10968 22584 11020 22593
rect 16948 22627 17000 22636
rect 6000 22516 6052 22568
rect 9864 22516 9916 22568
rect 10784 22516 10836 22568
rect 16948 22593 16957 22627
rect 16957 22593 16991 22627
rect 16991 22593 17000 22627
rect 16948 22584 17000 22593
rect 11796 22516 11848 22568
rect 12716 22516 12768 22568
rect 13820 22516 13872 22568
rect 18512 22729 18521 22763
rect 18521 22729 18555 22763
rect 18555 22729 18564 22763
rect 18512 22720 18564 22729
rect 19432 22720 19484 22772
rect 20812 22720 20864 22772
rect 20996 22720 21048 22772
rect 22192 22720 22244 22772
rect 24124 22720 24176 22772
rect 24676 22720 24728 22772
rect 25044 22763 25096 22772
rect 25044 22729 25053 22763
rect 25053 22729 25087 22763
rect 25087 22729 25096 22763
rect 25044 22720 25096 22729
rect 26148 22720 26200 22772
rect 21824 22695 21876 22704
rect 21824 22661 21833 22695
rect 21833 22661 21867 22695
rect 21867 22661 21876 22695
rect 21824 22652 21876 22661
rect 22100 22652 22152 22704
rect 22468 22652 22520 22704
rect 22560 22627 22612 22636
rect 22560 22593 22569 22627
rect 22569 22593 22603 22627
rect 22603 22593 22612 22627
rect 22560 22584 22612 22593
rect 24216 22627 24268 22636
rect 24216 22593 24225 22627
rect 24225 22593 24259 22627
rect 24259 22593 24268 22627
rect 24216 22584 24268 22593
rect 8392 22448 8444 22500
rect 4712 22380 4764 22432
rect 5540 22423 5592 22432
rect 5540 22389 5549 22423
rect 5549 22389 5583 22423
rect 5583 22389 5592 22423
rect 5540 22380 5592 22389
rect 6552 22423 6604 22432
rect 6552 22389 6561 22423
rect 6561 22389 6595 22423
rect 6595 22389 6604 22423
rect 6552 22380 6604 22389
rect 7104 22380 7156 22432
rect 10140 22380 10192 22432
rect 11152 22448 11204 22500
rect 14188 22491 14240 22500
rect 14188 22457 14222 22491
rect 14222 22457 14240 22491
rect 14188 22448 14240 22457
rect 16488 22448 16540 22500
rect 12624 22423 12676 22432
rect 12624 22389 12633 22423
rect 12633 22389 12667 22423
rect 12667 22389 12676 22423
rect 12624 22380 12676 22389
rect 16396 22423 16448 22432
rect 16396 22389 16405 22423
rect 16405 22389 16439 22423
rect 16439 22389 16448 22423
rect 16396 22380 16448 22389
rect 16764 22423 16816 22432
rect 16764 22389 16773 22423
rect 16773 22389 16807 22423
rect 16807 22389 16816 22423
rect 16764 22380 16816 22389
rect 18328 22380 18380 22432
rect 21456 22559 21508 22568
rect 21456 22525 21465 22559
rect 21465 22525 21499 22559
rect 21499 22525 21508 22559
rect 21456 22516 21508 22525
rect 22468 22559 22520 22568
rect 22468 22525 22477 22559
rect 22477 22525 22511 22559
rect 22511 22525 22520 22559
rect 22468 22516 22520 22525
rect 23480 22516 23532 22568
rect 25136 22516 25188 22568
rect 25320 22516 25372 22568
rect 19984 22448 20036 22500
rect 20352 22448 20404 22500
rect 23756 22448 23808 22500
rect 19524 22380 19576 22432
rect 20444 22380 20496 22432
rect 21824 22380 21876 22432
rect 22376 22423 22428 22432
rect 22376 22389 22385 22423
rect 22385 22389 22419 22423
rect 22419 22389 22428 22423
rect 22376 22380 22428 22389
rect 22928 22380 22980 22432
rect 23296 22423 23348 22432
rect 23296 22389 23305 22423
rect 23305 22389 23339 22423
rect 23339 22389 23348 22423
rect 23296 22380 23348 22389
rect 23480 22380 23532 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1216 22176 1268 22228
rect 2596 22176 2648 22228
rect 3056 22219 3108 22228
rect 3056 22185 3065 22219
rect 3065 22185 3099 22219
rect 3099 22185 3108 22219
rect 3056 22176 3108 22185
rect 5540 22176 5592 22228
rect 8668 22219 8720 22228
rect 8668 22185 8677 22219
rect 8677 22185 8711 22219
rect 8711 22185 8720 22219
rect 8668 22176 8720 22185
rect 9404 22219 9456 22228
rect 9404 22185 9413 22219
rect 9413 22185 9447 22219
rect 9447 22185 9456 22219
rect 9404 22176 9456 22185
rect 10048 22176 10100 22228
rect 1676 22108 1728 22160
rect 4620 22108 4672 22160
rect 2228 22015 2280 22024
rect 2228 21981 2237 22015
rect 2237 21981 2271 22015
rect 2271 21981 2280 22015
rect 2228 21972 2280 21981
rect 4528 22015 4580 22024
rect 4528 21981 4537 22015
rect 4537 21981 4571 22015
rect 4571 21981 4580 22015
rect 4528 21972 4580 21981
rect 5448 22040 5500 22092
rect 6368 22040 6420 22092
rect 10784 22176 10836 22228
rect 12440 22176 12492 22228
rect 16304 22219 16356 22228
rect 10692 22108 10744 22160
rect 11520 22108 11572 22160
rect 12256 22108 12308 22160
rect 12900 22108 12952 22160
rect 14188 22108 14240 22160
rect 14464 22108 14516 22160
rect 16304 22185 16313 22219
rect 16313 22185 16347 22219
rect 16347 22185 16356 22219
rect 16304 22176 16356 22185
rect 18696 22176 18748 22228
rect 20720 22176 20772 22228
rect 22376 22176 22428 22228
rect 22468 22176 22520 22228
rect 17132 22151 17184 22160
rect 17132 22117 17141 22151
rect 17141 22117 17175 22151
rect 17175 22117 17184 22151
rect 17132 22108 17184 22117
rect 20812 22108 20864 22160
rect 10324 22040 10376 22092
rect 11336 22083 11388 22092
rect 11336 22049 11345 22083
rect 11345 22049 11379 22083
rect 11379 22049 11388 22083
rect 11336 22040 11388 22049
rect 6092 21972 6144 22024
rect 9588 21972 9640 22024
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 3056 21904 3108 21956
rect 1584 21879 1636 21888
rect 1584 21845 1593 21879
rect 1593 21845 1627 21879
rect 1627 21845 1636 21879
rect 1584 21836 1636 21845
rect 1952 21836 2004 21888
rect 2872 21836 2924 21888
rect 3424 21836 3476 21888
rect 3608 21836 3660 21888
rect 5356 21904 5408 21956
rect 9864 21947 9916 21956
rect 9864 21913 9873 21947
rect 9873 21913 9907 21947
rect 9907 21913 9916 21947
rect 9864 21904 9916 21913
rect 14280 21947 14332 21956
rect 14280 21913 14289 21947
rect 14289 21913 14323 21947
rect 14323 21913 14332 21947
rect 14280 21904 14332 21913
rect 15384 22040 15436 22092
rect 17316 22040 17368 22092
rect 17868 22040 17920 22092
rect 20352 22083 20404 22092
rect 20352 22049 20361 22083
rect 20361 22049 20395 22083
rect 20395 22049 20404 22083
rect 23296 22108 23348 22160
rect 20352 22040 20404 22049
rect 22928 22040 22980 22092
rect 24860 22083 24912 22092
rect 24860 22049 24869 22083
rect 24869 22049 24903 22083
rect 24903 22049 24912 22083
rect 24860 22040 24912 22049
rect 25044 22083 25096 22092
rect 25044 22049 25053 22083
rect 25053 22049 25087 22083
rect 25087 22049 25096 22083
rect 25044 22040 25096 22049
rect 25320 22040 25372 22092
rect 14648 21972 14700 22024
rect 17408 22015 17460 22024
rect 17408 21981 17417 22015
rect 17417 21981 17451 22015
rect 17451 21981 17460 22015
rect 17408 21972 17460 21981
rect 18328 22015 18380 22024
rect 18328 21981 18337 22015
rect 18337 21981 18371 22015
rect 18371 21981 18380 22015
rect 18328 21972 18380 21981
rect 21732 21972 21784 22024
rect 14832 21904 14884 21956
rect 15844 21947 15896 21956
rect 15844 21913 15853 21947
rect 15853 21913 15887 21947
rect 15887 21913 15896 21947
rect 15844 21904 15896 21913
rect 16764 21947 16816 21956
rect 16764 21913 16773 21947
rect 16773 21913 16807 21947
rect 16807 21913 16816 21947
rect 16764 21904 16816 21913
rect 19708 21947 19760 21956
rect 19708 21913 19717 21947
rect 19717 21913 19751 21947
rect 19751 21913 19760 21947
rect 19708 21904 19760 21913
rect 22560 21904 22612 21956
rect 7656 21879 7708 21888
rect 7656 21845 7665 21879
rect 7665 21845 7699 21879
rect 7699 21845 7708 21879
rect 7656 21836 7708 21845
rect 8392 21836 8444 21888
rect 11428 21836 11480 21888
rect 12348 21836 12400 21888
rect 12900 21836 12952 21888
rect 14740 21879 14792 21888
rect 14740 21845 14749 21879
rect 14749 21845 14783 21879
rect 14783 21845 14792 21879
rect 14740 21836 14792 21845
rect 15568 21879 15620 21888
rect 15568 21845 15577 21879
rect 15577 21845 15611 21879
rect 15611 21845 15620 21879
rect 15568 21836 15620 21845
rect 16028 21836 16080 21888
rect 16948 21836 17000 21888
rect 18604 21836 18656 21888
rect 21548 21879 21600 21888
rect 21548 21845 21557 21879
rect 21557 21845 21591 21879
rect 21591 21845 21600 21879
rect 21548 21836 21600 21845
rect 21732 21836 21784 21888
rect 22192 21836 22244 21888
rect 23756 21972 23808 22024
rect 23940 22015 23992 22024
rect 23940 21981 23949 22015
rect 23949 21981 23983 22015
rect 23983 21981 23992 22015
rect 23940 21972 23992 21981
rect 24032 22015 24084 22024
rect 24032 21981 24041 22015
rect 24041 21981 24075 22015
rect 24075 21981 24084 22015
rect 24032 21972 24084 21981
rect 24216 21972 24268 22024
rect 22928 21904 22980 21956
rect 23204 21836 23256 21888
rect 24216 21836 24268 21888
rect 25228 21879 25280 21888
rect 25228 21845 25237 21879
rect 25237 21845 25271 21879
rect 25271 21845 25280 21879
rect 25228 21836 25280 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1584 21632 1636 21684
rect 2044 21632 2096 21684
rect 2596 21675 2648 21684
rect 2596 21641 2605 21675
rect 2605 21641 2639 21675
rect 2639 21641 2648 21675
rect 2596 21632 2648 21641
rect 2872 21632 2924 21684
rect 5448 21632 5500 21684
rect 6368 21632 6420 21684
rect 10324 21675 10376 21684
rect 10324 21641 10333 21675
rect 10333 21641 10367 21675
rect 10367 21641 10376 21675
rect 10324 21632 10376 21641
rect 10692 21675 10744 21684
rect 10692 21641 10701 21675
rect 10701 21641 10735 21675
rect 10735 21641 10744 21675
rect 10692 21632 10744 21641
rect 11428 21632 11480 21684
rect 11612 21632 11664 21684
rect 12256 21675 12308 21684
rect 10048 21564 10100 21616
rect 10508 21564 10560 21616
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 14188 21632 14240 21684
rect 16488 21632 16540 21684
rect 17868 21675 17920 21684
rect 17868 21641 17877 21675
rect 17877 21641 17911 21675
rect 17911 21641 17920 21675
rect 17868 21632 17920 21641
rect 22284 21632 22336 21684
rect 24032 21632 24084 21684
rect 25596 21675 25648 21684
rect 25596 21641 25605 21675
rect 25605 21641 25639 21675
rect 25639 21641 25648 21675
rect 25596 21632 25648 21641
rect 2228 21539 2280 21548
rect 2228 21505 2237 21539
rect 2237 21505 2271 21539
rect 2271 21505 2280 21539
rect 2228 21496 2280 21505
rect 7196 21496 7248 21548
rect 7656 21496 7708 21548
rect 7932 21496 7984 21548
rect 8300 21539 8352 21548
rect 8300 21505 8309 21539
rect 8309 21505 8343 21539
rect 8343 21505 8352 21539
rect 8300 21496 8352 21505
rect 10876 21496 10928 21548
rect 11336 21539 11388 21548
rect 11336 21505 11345 21539
rect 11345 21505 11379 21539
rect 11379 21505 11388 21539
rect 11336 21496 11388 21505
rect 20904 21564 20956 21616
rect 22376 21564 22428 21616
rect 23572 21564 23624 21616
rect 24860 21564 24912 21616
rect 3332 21471 3384 21480
rect 3332 21437 3341 21471
rect 3341 21437 3375 21471
rect 3375 21437 3384 21471
rect 3332 21428 3384 21437
rect 6092 21428 6144 21480
rect 9864 21428 9916 21480
rect 11152 21471 11204 21480
rect 11152 21437 11161 21471
rect 11161 21437 11195 21471
rect 11195 21437 11204 21471
rect 11152 21428 11204 21437
rect 12624 21471 12676 21480
rect 12624 21437 12633 21471
rect 12633 21437 12667 21471
rect 12667 21437 12676 21471
rect 12624 21428 12676 21437
rect 15568 21539 15620 21548
rect 15568 21505 15577 21539
rect 15577 21505 15611 21539
rect 15611 21505 15620 21539
rect 15568 21496 15620 21505
rect 17408 21496 17460 21548
rect 13360 21428 13412 21480
rect 14372 21428 14424 21480
rect 16304 21428 16356 21480
rect 2596 21360 2648 21412
rect 3608 21403 3660 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 1952 21335 2004 21344
rect 1952 21301 1961 21335
rect 1961 21301 1995 21335
rect 1995 21301 2004 21335
rect 1952 21292 2004 21301
rect 3608 21369 3642 21403
rect 3642 21369 3660 21403
rect 3608 21360 3660 21369
rect 3976 21292 4028 21344
rect 4436 21292 4488 21344
rect 6460 21292 6512 21344
rect 7196 21335 7248 21344
rect 7196 21301 7205 21335
rect 7205 21301 7239 21335
rect 7239 21301 7248 21335
rect 7196 21292 7248 21301
rect 8576 21335 8628 21344
rect 8576 21301 8585 21335
rect 8585 21301 8619 21335
rect 8619 21301 8628 21335
rect 8576 21292 8628 21301
rect 12900 21360 12952 21412
rect 16488 21360 16540 21412
rect 17132 21360 17184 21412
rect 9680 21335 9732 21344
rect 9680 21301 9689 21335
rect 9689 21301 9723 21335
rect 9723 21301 9732 21335
rect 9680 21292 9732 21301
rect 9864 21292 9916 21344
rect 10140 21292 10192 21344
rect 10692 21292 10744 21344
rect 15292 21292 15344 21344
rect 16764 21335 16816 21344
rect 16764 21301 16773 21335
rect 16773 21301 16807 21335
rect 16807 21301 16816 21335
rect 16764 21292 16816 21301
rect 17316 21292 17368 21344
rect 17684 21292 17736 21344
rect 18328 21335 18380 21344
rect 18328 21301 18337 21335
rect 18337 21301 18371 21335
rect 18371 21301 18380 21335
rect 18604 21360 18656 21412
rect 19156 21360 19208 21412
rect 18328 21292 18380 21301
rect 20352 21335 20404 21344
rect 20352 21301 20361 21335
rect 20361 21301 20395 21335
rect 20395 21301 20404 21335
rect 20352 21292 20404 21301
rect 20720 21292 20772 21344
rect 24032 21496 24084 21548
rect 24492 21539 24544 21548
rect 24492 21505 24501 21539
rect 24501 21505 24535 21539
rect 24535 21505 24544 21539
rect 24492 21496 24544 21505
rect 21548 21428 21600 21480
rect 23572 21428 23624 21480
rect 24768 21428 24820 21480
rect 25320 21428 25372 21480
rect 24124 21360 24176 21412
rect 21272 21335 21324 21344
rect 21272 21301 21281 21335
rect 21281 21301 21315 21335
rect 21315 21301 21324 21335
rect 21272 21292 21324 21301
rect 21732 21292 21784 21344
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 25044 21335 25096 21344
rect 25044 21301 25053 21335
rect 25053 21301 25087 21335
rect 25087 21301 25096 21335
rect 25044 21292 25096 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1492 21088 1544 21140
rect 1768 21088 1820 21140
rect 2412 21131 2464 21140
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 2412 21097 2421 21131
rect 2421 21097 2455 21131
rect 2455 21097 2464 21131
rect 2412 21088 2464 21097
rect 3332 21088 3384 21140
rect 4436 21088 4488 21140
rect 4712 21088 4764 21140
rect 6368 21131 6420 21140
rect 6368 21097 6377 21131
rect 6377 21097 6411 21131
rect 6411 21097 6420 21131
rect 6368 21088 6420 21097
rect 7656 21088 7708 21140
rect 10048 21088 10100 21140
rect 11152 21088 11204 21140
rect 11520 21131 11572 21140
rect 11520 21097 11529 21131
rect 11529 21097 11563 21131
rect 11563 21097 11572 21131
rect 11520 21088 11572 21097
rect 12164 21088 12216 21140
rect 12348 21088 12400 21140
rect 12532 21088 12584 21140
rect 13360 21131 13412 21140
rect 13360 21097 13369 21131
rect 13369 21097 13403 21131
rect 13403 21097 13412 21131
rect 13360 21088 13412 21097
rect 15660 21131 15712 21140
rect 2596 21020 2648 21072
rect 4068 21020 4120 21072
rect 10968 21063 11020 21072
rect 10968 21029 10977 21063
rect 10977 21029 11011 21063
rect 11011 21029 11020 21063
rect 10968 21020 11020 21029
rect 14280 21020 14332 21072
rect 15660 21097 15669 21131
rect 15669 21097 15703 21131
rect 15703 21097 15712 21131
rect 15660 21088 15712 21097
rect 15936 21088 15988 21140
rect 16304 21088 16356 21140
rect 17868 21088 17920 21140
rect 16948 21063 17000 21072
rect 16948 21029 16982 21063
rect 16982 21029 17000 21063
rect 16948 21020 17000 21029
rect 17408 21020 17460 21072
rect 18604 21063 18656 21072
rect 18604 21029 18613 21063
rect 18613 21029 18647 21063
rect 18647 21029 18656 21063
rect 18604 21020 18656 21029
rect 3332 20952 3384 21004
rect 4160 20952 4212 21004
rect 7012 20952 7064 21004
rect 7472 20995 7524 21004
rect 7472 20961 7481 20995
rect 7481 20961 7515 20995
rect 7515 20961 7524 20995
rect 7472 20952 7524 20961
rect 7748 20952 7800 21004
rect 8300 20952 8352 21004
rect 9588 20952 9640 21004
rect 10876 20995 10928 21004
rect 10876 20961 10885 20995
rect 10885 20961 10919 20995
rect 10919 20961 10928 20995
rect 10876 20952 10928 20961
rect 12440 20995 12492 21004
rect 12440 20961 12449 20995
rect 12449 20961 12483 20995
rect 12483 20961 12492 20995
rect 12440 20952 12492 20961
rect 14832 20952 14884 21004
rect 15844 20952 15896 21004
rect 16120 20952 16172 21004
rect 2780 20884 2832 20936
rect 3516 20884 3568 20936
rect 5356 20884 5408 20936
rect 7564 20927 7616 20936
rect 6920 20859 6972 20868
rect 6920 20825 6929 20859
rect 6929 20825 6963 20859
rect 6963 20825 6972 20859
rect 6920 20816 6972 20825
rect 7564 20893 7573 20927
rect 7573 20893 7607 20927
rect 7607 20893 7616 20927
rect 7564 20884 7616 20893
rect 8944 20884 8996 20936
rect 11060 20927 11112 20936
rect 11060 20893 11069 20927
rect 11069 20893 11103 20927
rect 11103 20893 11112 20927
rect 11060 20884 11112 20893
rect 12348 20884 12400 20936
rect 12716 20927 12768 20936
rect 12716 20893 12725 20927
rect 12725 20893 12759 20927
rect 12759 20893 12768 20927
rect 12716 20884 12768 20893
rect 13452 20816 13504 20868
rect 14924 20816 14976 20868
rect 19064 21088 19116 21140
rect 22744 21131 22796 21140
rect 22744 21097 22753 21131
rect 22753 21097 22787 21131
rect 22787 21097 22796 21131
rect 22744 21088 22796 21097
rect 23940 21088 23992 21140
rect 22192 21020 22244 21072
rect 22928 21020 22980 21072
rect 19340 20952 19392 21004
rect 21180 20952 21232 21004
rect 22560 20995 22612 21004
rect 22560 20961 22569 20995
rect 22569 20961 22603 20995
rect 22603 20961 22612 20995
rect 22560 20952 22612 20961
rect 23940 20952 23992 21004
rect 24676 20952 24728 21004
rect 19616 20927 19668 20936
rect 19616 20893 19625 20927
rect 19625 20893 19659 20927
rect 19659 20893 19668 20927
rect 19616 20884 19668 20893
rect 20352 20884 20404 20936
rect 20720 20927 20772 20936
rect 20720 20893 20729 20927
rect 20729 20893 20763 20927
rect 20763 20893 20772 20927
rect 20720 20884 20772 20893
rect 21364 20927 21416 20936
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 24216 20884 24268 20936
rect 24492 20927 24544 20936
rect 24492 20893 24501 20927
rect 24501 20893 24535 20927
rect 24535 20893 24544 20927
rect 24492 20884 24544 20893
rect 2412 20748 2464 20800
rect 3608 20748 3660 20800
rect 5448 20791 5500 20800
rect 5448 20757 5457 20791
rect 5457 20757 5491 20791
rect 5491 20757 5500 20791
rect 5448 20748 5500 20757
rect 7012 20791 7064 20800
rect 7012 20757 7021 20791
rect 7021 20757 7055 20791
rect 7055 20757 7064 20791
rect 7012 20748 7064 20757
rect 8392 20791 8444 20800
rect 8392 20757 8401 20791
rect 8401 20757 8435 20791
rect 8435 20757 8444 20791
rect 8392 20748 8444 20757
rect 9036 20791 9088 20800
rect 9036 20757 9045 20791
rect 9045 20757 9079 20791
rect 9079 20757 9088 20791
rect 9036 20748 9088 20757
rect 10232 20791 10284 20800
rect 10232 20757 10241 20791
rect 10241 20757 10275 20791
rect 10275 20757 10284 20791
rect 10232 20748 10284 20757
rect 14372 20748 14424 20800
rect 15384 20748 15436 20800
rect 16028 20791 16080 20800
rect 16028 20757 16037 20791
rect 16037 20757 16071 20791
rect 16071 20757 16080 20791
rect 16028 20748 16080 20757
rect 20720 20748 20772 20800
rect 21824 20748 21876 20800
rect 22100 20748 22152 20800
rect 23756 20748 23808 20800
rect 24032 20748 24084 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1860 20544 1912 20596
rect 2228 20544 2280 20596
rect 3332 20544 3384 20596
rect 3516 20544 3568 20596
rect 4528 20544 4580 20596
rect 6828 20587 6880 20596
rect 2320 20408 2372 20460
rect 2688 20408 2740 20460
rect 3332 20451 3384 20460
rect 3332 20417 3341 20451
rect 3341 20417 3375 20451
rect 3375 20417 3384 20451
rect 3332 20408 3384 20417
rect 1860 20340 1912 20392
rect 4160 20408 4212 20460
rect 6828 20553 6837 20587
rect 6837 20553 6871 20587
rect 6871 20553 6880 20587
rect 6828 20544 6880 20553
rect 9588 20544 9640 20596
rect 10968 20544 11020 20596
rect 14280 20544 14332 20596
rect 14832 20587 14884 20596
rect 14832 20553 14841 20587
rect 14841 20553 14875 20587
rect 14875 20553 14884 20587
rect 14832 20544 14884 20553
rect 5448 20476 5500 20528
rect 6276 20519 6328 20528
rect 6276 20485 6285 20519
rect 6285 20485 6319 20519
rect 6319 20485 6328 20519
rect 6276 20476 6328 20485
rect 7564 20476 7616 20528
rect 7012 20408 7064 20460
rect 16120 20544 16172 20596
rect 17684 20544 17736 20596
rect 17868 20587 17920 20596
rect 17868 20553 17877 20587
rect 17877 20553 17911 20587
rect 17911 20553 17920 20587
rect 17868 20544 17920 20553
rect 18972 20544 19024 20596
rect 19248 20544 19300 20596
rect 22192 20544 22244 20596
rect 22560 20544 22612 20596
rect 25412 20587 25464 20596
rect 25412 20553 25421 20587
rect 25421 20553 25455 20587
rect 25455 20553 25464 20587
rect 25412 20544 25464 20553
rect 19340 20408 19392 20460
rect 20352 20408 20404 20460
rect 24676 20451 24728 20460
rect 3240 20315 3292 20324
rect 3240 20281 3249 20315
rect 3249 20281 3283 20315
rect 3283 20281 3292 20315
rect 3240 20272 3292 20281
rect 6920 20272 6972 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 2596 20204 2648 20256
rect 4436 20204 4488 20256
rect 4804 20247 4856 20256
rect 4804 20213 4813 20247
rect 4813 20213 4847 20247
rect 4847 20213 4856 20247
rect 4804 20204 4856 20213
rect 5448 20247 5500 20256
rect 5448 20213 5457 20247
rect 5457 20213 5491 20247
rect 5491 20213 5500 20247
rect 5448 20204 5500 20213
rect 7472 20272 7524 20324
rect 7196 20247 7248 20256
rect 7196 20213 7205 20247
rect 7205 20213 7239 20247
rect 7239 20213 7248 20247
rect 7196 20204 7248 20213
rect 7656 20204 7708 20256
rect 8024 20204 8076 20256
rect 11612 20340 11664 20392
rect 12256 20340 12308 20392
rect 12532 20340 12584 20392
rect 16028 20340 16080 20392
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 20812 20340 20864 20392
rect 24032 20383 24084 20392
rect 24032 20349 24041 20383
rect 24041 20349 24075 20383
rect 24075 20349 24084 20383
rect 24032 20340 24084 20349
rect 8852 20315 8904 20324
rect 8852 20281 8886 20315
rect 8886 20281 8904 20315
rect 8852 20272 8904 20281
rect 9128 20272 9180 20324
rect 12348 20272 12400 20324
rect 17684 20272 17736 20324
rect 20352 20315 20404 20324
rect 20352 20281 20361 20315
rect 20361 20281 20395 20315
rect 20395 20281 20404 20315
rect 20352 20272 20404 20281
rect 23940 20272 23992 20324
rect 24676 20417 24685 20451
rect 24685 20417 24719 20451
rect 24719 20417 24728 20451
rect 24676 20408 24728 20417
rect 8760 20204 8812 20256
rect 9588 20204 9640 20256
rect 10048 20204 10100 20256
rect 11060 20204 11112 20256
rect 11612 20247 11664 20256
rect 11612 20213 11621 20247
rect 11621 20213 11655 20247
rect 11655 20213 11664 20247
rect 11612 20204 11664 20213
rect 13820 20247 13872 20256
rect 13820 20213 13829 20247
rect 13829 20213 13863 20247
rect 13863 20213 13872 20247
rect 13820 20204 13872 20213
rect 16764 20247 16816 20256
rect 16764 20213 16773 20247
rect 16773 20213 16807 20247
rect 16807 20213 16816 20247
rect 16764 20204 16816 20213
rect 18788 20204 18840 20256
rect 20076 20204 20128 20256
rect 20812 20247 20864 20256
rect 20812 20213 20821 20247
rect 20821 20213 20855 20247
rect 20855 20213 20864 20247
rect 20812 20204 20864 20213
rect 20904 20204 20956 20256
rect 23664 20247 23716 20256
rect 23664 20213 23673 20247
rect 23673 20213 23707 20247
rect 23707 20213 23716 20247
rect 23664 20204 23716 20213
rect 24124 20247 24176 20256
rect 24124 20213 24133 20247
rect 24133 20213 24167 20247
rect 24167 20213 24176 20247
rect 24124 20204 24176 20213
rect 25596 20204 25648 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1860 20000 1912 20052
rect 2320 20000 2372 20052
rect 2780 20000 2832 20052
rect 2872 20043 2924 20052
rect 2872 20009 2881 20043
rect 2881 20009 2915 20043
rect 2915 20009 2924 20043
rect 2872 20000 2924 20009
rect 4068 20043 4120 20052
rect 4068 20009 4077 20043
rect 4077 20009 4111 20043
rect 4111 20009 4120 20043
rect 4068 20000 4120 20009
rect 4436 20043 4488 20052
rect 4436 20009 4445 20043
rect 4445 20009 4479 20043
rect 4479 20009 4488 20043
rect 4436 20000 4488 20009
rect 7012 20000 7064 20052
rect 8852 20000 8904 20052
rect 11152 20000 11204 20052
rect 13728 20000 13780 20052
rect 14556 20000 14608 20052
rect 15844 20000 15896 20052
rect 16580 20000 16632 20052
rect 17684 20000 17736 20052
rect 848 19932 900 19984
rect 3332 19932 3384 19984
rect 6276 19932 6328 19984
rect 7196 19932 7248 19984
rect 12716 19932 12768 19984
rect 16948 19932 17000 19984
rect 19340 20000 19392 20052
rect 20812 20000 20864 20052
rect 21364 20000 21416 20052
rect 21916 20043 21968 20052
rect 21916 20009 21925 20043
rect 21925 20009 21959 20043
rect 21959 20009 21968 20043
rect 21916 20000 21968 20009
rect 24124 20000 24176 20052
rect 24860 20000 24912 20052
rect 25412 20000 25464 20052
rect 2596 19864 2648 19916
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 3148 19864 3200 19916
rect 4160 19864 4212 19916
rect 2320 19839 2372 19848
rect 2320 19805 2329 19839
rect 2329 19805 2363 19839
rect 2363 19805 2372 19839
rect 2320 19796 2372 19805
rect 4528 19839 4580 19848
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 5448 19907 5500 19916
rect 5448 19873 5457 19907
rect 5457 19873 5491 19907
rect 5491 19873 5500 19907
rect 5448 19864 5500 19873
rect 6000 19864 6052 19916
rect 8484 19864 8536 19916
rect 9312 19864 9364 19916
rect 6920 19728 6972 19780
rect 3792 19660 3844 19712
rect 4344 19660 4396 19712
rect 9220 19660 9272 19712
rect 12256 19864 12308 19916
rect 9588 19796 9640 19848
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 10048 19660 10100 19712
rect 11704 19728 11756 19780
rect 11520 19660 11572 19712
rect 12440 19728 12492 19780
rect 15292 19864 15344 19916
rect 16580 19864 16632 19916
rect 18052 19864 18104 19916
rect 18604 19907 18656 19916
rect 18604 19873 18638 19907
rect 18638 19873 18656 19907
rect 18604 19864 18656 19873
rect 21548 19864 21600 19916
rect 22652 19907 22704 19916
rect 22652 19873 22686 19907
rect 22686 19873 22704 19907
rect 22652 19864 22704 19873
rect 24216 19864 24268 19916
rect 15476 19796 15528 19848
rect 15752 19839 15804 19848
rect 15752 19805 15761 19839
rect 15761 19805 15795 19839
rect 15795 19805 15804 19839
rect 15752 19796 15804 19805
rect 12348 19660 12400 19712
rect 13360 19660 13412 19712
rect 14832 19660 14884 19712
rect 16764 19796 16816 19848
rect 22284 19796 22336 19848
rect 23756 19796 23808 19848
rect 24124 19796 24176 19848
rect 25320 19839 25372 19848
rect 25320 19805 25329 19839
rect 25329 19805 25363 19839
rect 25363 19805 25372 19839
rect 25320 19796 25372 19805
rect 25596 19796 25648 19848
rect 20904 19660 20956 19712
rect 21180 19703 21232 19712
rect 21180 19669 21189 19703
rect 21189 19669 21223 19703
rect 21223 19669 21232 19703
rect 21180 19660 21232 19669
rect 21456 19703 21508 19712
rect 21456 19669 21465 19703
rect 21465 19669 21499 19703
rect 21499 19669 21508 19703
rect 21456 19660 21508 19669
rect 23756 19703 23808 19712
rect 23756 19669 23765 19703
rect 23765 19669 23799 19703
rect 23799 19669 23808 19703
rect 23756 19660 23808 19669
rect 24860 19703 24912 19712
rect 24860 19669 24869 19703
rect 24869 19669 24903 19703
rect 24903 19669 24912 19703
rect 24860 19660 24912 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2780 19499 2832 19508
rect 2780 19465 2789 19499
rect 2789 19465 2823 19499
rect 2823 19465 2832 19499
rect 2780 19456 2832 19465
rect 4068 19456 4120 19508
rect 4436 19456 4488 19508
rect 4804 19456 4856 19508
rect 6092 19456 6144 19508
rect 9680 19456 9732 19508
rect 15292 19456 15344 19508
rect 16764 19456 16816 19508
rect 17684 19456 17736 19508
rect 2320 19388 2372 19440
rect 3884 19388 3936 19440
rect 1860 19320 1912 19372
rect 3608 19320 3660 19372
rect 3792 19320 3844 19372
rect 1676 19252 1728 19304
rect 2780 19252 2832 19304
rect 3884 19252 3936 19304
rect 3976 19252 4028 19304
rect 1676 19116 1728 19168
rect 2044 19116 2096 19168
rect 3608 19159 3660 19168
rect 3608 19125 3617 19159
rect 3617 19125 3651 19159
rect 3651 19125 3660 19159
rect 3608 19116 3660 19125
rect 4620 19116 4672 19168
rect 11428 19388 11480 19440
rect 5448 19320 5500 19372
rect 7564 19320 7616 19372
rect 9036 19320 9088 19372
rect 10140 19320 10192 19372
rect 10876 19320 10928 19372
rect 13544 19363 13596 19372
rect 13544 19329 13553 19363
rect 13553 19329 13587 19363
rect 13587 19329 13596 19363
rect 13544 19320 13596 19329
rect 6184 19252 6236 19304
rect 5172 19116 5224 19168
rect 9588 19252 9640 19304
rect 9772 19252 9824 19304
rect 11796 19295 11848 19304
rect 11796 19261 11805 19295
rect 11805 19261 11839 19295
rect 11839 19261 11848 19295
rect 11796 19252 11848 19261
rect 12348 19184 12400 19236
rect 6092 19116 6144 19168
rect 6736 19116 6788 19168
rect 6920 19116 6972 19168
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 7840 19159 7892 19168
rect 7288 19116 7340 19125
rect 7840 19125 7849 19159
rect 7849 19125 7883 19159
rect 7883 19125 7892 19159
rect 7840 19116 7892 19125
rect 8576 19116 8628 19168
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 9496 19116 9548 19168
rect 9956 19159 10008 19168
rect 9956 19125 9965 19159
rect 9965 19125 9999 19159
rect 9999 19125 10008 19159
rect 9956 19116 10008 19125
rect 11428 19159 11480 19168
rect 11428 19125 11437 19159
rect 11437 19125 11471 19159
rect 11471 19125 11480 19159
rect 11428 19116 11480 19125
rect 12256 19159 12308 19168
rect 12256 19125 12265 19159
rect 12265 19125 12299 19159
rect 12299 19125 12308 19159
rect 12256 19116 12308 19125
rect 12532 19116 12584 19168
rect 15844 19320 15896 19372
rect 17040 19320 17092 19372
rect 20352 19456 20404 19508
rect 25320 19456 25372 19508
rect 25596 19431 25648 19440
rect 25596 19397 25605 19431
rect 25605 19397 25639 19431
rect 25639 19397 25648 19431
rect 25596 19388 25648 19397
rect 20996 19363 21048 19372
rect 20996 19329 21005 19363
rect 21005 19329 21039 19363
rect 21039 19329 21048 19363
rect 20996 19320 21048 19329
rect 14188 19252 14240 19304
rect 14832 19295 14884 19304
rect 14832 19261 14866 19295
rect 14866 19261 14884 19295
rect 14832 19252 14884 19261
rect 15936 19252 15988 19304
rect 14096 19184 14148 19236
rect 14280 19184 14332 19236
rect 13360 19116 13412 19168
rect 13728 19116 13780 19168
rect 14556 19116 14608 19168
rect 16948 19116 17000 19168
rect 22008 19184 22060 19236
rect 22284 19184 22336 19236
rect 23756 19184 23808 19236
rect 24492 19184 24544 19236
rect 18604 19116 18656 19168
rect 20996 19116 21048 19168
rect 23296 19116 23348 19168
rect 24032 19116 24084 19168
rect 25044 19159 25096 19168
rect 25044 19125 25053 19159
rect 25053 19125 25087 19159
rect 25087 19125 25096 19159
rect 25044 19116 25096 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1952 18912 2004 18964
rect 3976 18912 4028 18964
rect 4988 18912 5040 18964
rect 7196 18912 7248 18964
rect 10876 18955 10928 18964
rect 10876 18921 10885 18955
rect 10885 18921 10919 18955
rect 10919 18921 10928 18955
rect 10876 18912 10928 18921
rect 11060 18912 11112 18964
rect 13820 18955 13872 18964
rect 13820 18921 13829 18955
rect 13829 18921 13863 18955
rect 13863 18921 13872 18955
rect 13820 18912 13872 18921
rect 15292 18912 15344 18964
rect 16856 18912 16908 18964
rect 19064 18955 19116 18964
rect 19064 18921 19073 18955
rect 19073 18921 19107 18955
rect 19107 18921 19116 18955
rect 19064 18912 19116 18921
rect 21824 18955 21876 18964
rect 21824 18921 21833 18955
rect 21833 18921 21867 18955
rect 21867 18921 21876 18955
rect 21824 18912 21876 18921
rect 22284 18912 22336 18964
rect 22836 18912 22888 18964
rect 24860 18955 24912 18964
rect 24860 18921 24869 18955
rect 24869 18921 24903 18955
rect 24903 18921 24912 18955
rect 24860 18912 24912 18921
rect 25504 18912 25556 18964
rect 2964 18844 3016 18896
rect 3424 18844 3476 18896
rect 4804 18844 4856 18896
rect 6920 18887 6972 18896
rect 6920 18853 6929 18887
rect 6929 18853 6963 18887
rect 6963 18853 6972 18887
rect 6920 18844 6972 18853
rect 1492 18776 1544 18828
rect 4712 18776 4764 18828
rect 5080 18776 5132 18828
rect 2872 18751 2924 18760
rect 2872 18717 2881 18751
rect 2881 18717 2915 18751
rect 2915 18717 2924 18751
rect 2872 18708 2924 18717
rect 3608 18708 3660 18760
rect 4436 18708 4488 18760
rect 3240 18640 3292 18692
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 3424 18572 3476 18624
rect 4528 18572 4580 18624
rect 6092 18708 6144 18760
rect 5172 18683 5224 18692
rect 5172 18649 5181 18683
rect 5181 18649 5215 18683
rect 5215 18649 5224 18683
rect 5172 18640 5224 18649
rect 7104 18708 7156 18760
rect 7564 18844 7616 18896
rect 7288 18640 7340 18692
rect 7840 18751 7892 18760
rect 7840 18717 7849 18751
rect 7849 18717 7883 18751
rect 7883 18717 7892 18751
rect 7840 18708 7892 18717
rect 10232 18819 10284 18828
rect 10232 18785 10241 18819
rect 10241 18785 10275 18819
rect 10275 18785 10284 18819
rect 10232 18776 10284 18785
rect 11336 18776 11388 18828
rect 13636 18844 13688 18896
rect 14096 18844 14148 18896
rect 18696 18844 18748 18896
rect 19156 18844 19208 18896
rect 13544 18776 13596 18828
rect 14832 18776 14884 18828
rect 16304 18819 16356 18828
rect 16304 18785 16313 18819
rect 16313 18785 16347 18819
rect 16347 18785 16356 18819
rect 16304 18776 16356 18785
rect 8852 18708 8904 18760
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 10508 18751 10560 18760
rect 10508 18717 10517 18751
rect 10517 18717 10551 18751
rect 10551 18717 10560 18751
rect 10508 18708 10560 18717
rect 11428 18751 11480 18760
rect 11428 18717 11437 18751
rect 11437 18717 11471 18751
rect 11471 18717 11480 18751
rect 11428 18708 11480 18717
rect 16396 18751 16448 18760
rect 16396 18717 16405 18751
rect 16405 18717 16439 18751
rect 16439 18717 16448 18751
rect 16396 18708 16448 18717
rect 16856 18708 16908 18760
rect 9680 18640 9732 18692
rect 19064 18776 19116 18828
rect 21824 18776 21876 18828
rect 18052 18751 18104 18760
rect 18052 18717 18061 18751
rect 18061 18717 18095 18751
rect 18095 18717 18104 18751
rect 18052 18708 18104 18717
rect 18604 18708 18656 18760
rect 22284 18751 22336 18760
rect 19340 18640 19392 18692
rect 22284 18717 22293 18751
rect 22293 18717 22327 18751
rect 22327 18717 22336 18751
rect 22284 18708 22336 18717
rect 22652 18844 22704 18896
rect 24492 18887 24544 18896
rect 24492 18853 24501 18887
rect 24501 18853 24535 18887
rect 24535 18853 24544 18887
rect 24492 18844 24544 18853
rect 25596 18844 25648 18896
rect 23756 18819 23808 18828
rect 23756 18785 23765 18819
rect 23765 18785 23799 18819
rect 23799 18785 23808 18819
rect 23756 18776 23808 18785
rect 23940 18751 23992 18760
rect 23940 18717 23949 18751
rect 23949 18717 23983 18751
rect 23983 18717 23992 18751
rect 23940 18708 23992 18717
rect 25412 18776 25464 18828
rect 25596 18708 25648 18760
rect 6184 18572 6236 18624
rect 8484 18615 8536 18624
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 9036 18572 9088 18624
rect 9864 18615 9916 18624
rect 9864 18581 9873 18615
rect 9873 18581 9907 18615
rect 9907 18581 9916 18615
rect 9864 18572 9916 18581
rect 12164 18572 12216 18624
rect 15476 18615 15528 18624
rect 15476 18581 15485 18615
rect 15485 18581 15519 18615
rect 15519 18581 15528 18615
rect 15476 18572 15528 18581
rect 16580 18572 16632 18624
rect 19524 18572 19576 18624
rect 20628 18572 20680 18624
rect 21548 18572 21600 18624
rect 22836 18615 22888 18624
rect 22836 18581 22845 18615
rect 22845 18581 22879 18615
rect 22879 18581 22888 18615
rect 22836 18572 22888 18581
rect 23572 18572 23624 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2964 18411 3016 18420
rect 2964 18377 2973 18411
rect 2973 18377 3007 18411
rect 3007 18377 3016 18411
rect 2964 18368 3016 18377
rect 3792 18368 3844 18420
rect 5080 18411 5132 18420
rect 5080 18377 5089 18411
rect 5089 18377 5123 18411
rect 5123 18377 5132 18411
rect 5080 18368 5132 18377
rect 7748 18368 7800 18420
rect 8392 18368 8444 18420
rect 4528 18343 4580 18352
rect 4528 18309 4537 18343
rect 4537 18309 4571 18343
rect 4571 18309 4580 18343
rect 4528 18300 4580 18309
rect 6092 18300 6144 18352
rect 7840 18343 7892 18352
rect 7840 18309 7849 18343
rect 7849 18309 7883 18343
rect 7883 18309 7892 18343
rect 7840 18300 7892 18309
rect 1952 18232 2004 18284
rect 8484 18275 8536 18284
rect 2964 18164 3016 18216
rect 8484 18241 8493 18275
rect 8493 18241 8527 18275
rect 8527 18241 8536 18275
rect 8484 18232 8536 18241
rect 3792 18164 3844 18216
rect 4712 18164 4764 18216
rect 1676 18096 1728 18148
rect 1400 18028 1452 18080
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 2872 18096 2924 18148
rect 4252 18096 4304 18148
rect 8208 18164 8260 18216
rect 8760 18164 8812 18216
rect 9680 18207 9732 18216
rect 9680 18173 9714 18207
rect 9714 18173 9732 18207
rect 7196 18096 7248 18148
rect 7748 18096 7800 18148
rect 9680 18164 9732 18173
rect 11060 18096 11112 18148
rect 12624 18368 12676 18420
rect 14188 18411 14240 18420
rect 14188 18377 14197 18411
rect 14197 18377 14231 18411
rect 14231 18377 14240 18411
rect 14188 18368 14240 18377
rect 16304 18368 16356 18420
rect 5172 18028 5224 18080
rect 5816 18071 5868 18080
rect 5816 18037 5825 18071
rect 5825 18037 5859 18071
rect 5859 18037 5868 18071
rect 5816 18028 5868 18037
rect 6644 18028 6696 18080
rect 7288 18028 7340 18080
rect 8760 18028 8812 18080
rect 9680 18028 9732 18080
rect 11428 18028 11480 18080
rect 11796 18028 11848 18080
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 13636 18232 13688 18284
rect 18052 18368 18104 18420
rect 19340 18368 19392 18420
rect 23480 18411 23532 18420
rect 23480 18377 23489 18411
rect 23489 18377 23523 18411
rect 23523 18377 23532 18411
rect 23480 18368 23532 18377
rect 22836 18232 22888 18284
rect 24860 18368 24912 18420
rect 26240 18411 26292 18420
rect 26240 18377 26249 18411
rect 26249 18377 26283 18411
rect 26283 18377 26292 18411
rect 26240 18368 26292 18377
rect 25044 18343 25096 18352
rect 25044 18309 25053 18343
rect 25053 18309 25087 18343
rect 25087 18309 25096 18343
rect 25044 18300 25096 18309
rect 24216 18275 24268 18284
rect 24216 18241 24225 18275
rect 24225 18241 24259 18275
rect 24259 18241 24268 18275
rect 24216 18232 24268 18241
rect 12624 18164 12676 18216
rect 14556 18207 14608 18216
rect 14556 18173 14590 18207
rect 14590 18173 14608 18207
rect 14556 18164 14608 18173
rect 19248 18164 19300 18216
rect 22468 18164 22520 18216
rect 23664 18164 23716 18216
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 15568 18096 15620 18148
rect 16396 18096 16448 18148
rect 22284 18096 22336 18148
rect 12440 18071 12492 18080
rect 12440 18037 12449 18071
rect 12449 18037 12483 18071
rect 12483 18037 12492 18071
rect 12440 18028 12492 18037
rect 15292 18028 15344 18080
rect 18512 18071 18564 18080
rect 18512 18037 18521 18071
rect 18521 18037 18555 18071
rect 18555 18037 18564 18071
rect 18512 18028 18564 18037
rect 19064 18071 19116 18080
rect 19064 18037 19073 18071
rect 19073 18037 19107 18071
rect 19107 18037 19116 18071
rect 19064 18028 19116 18037
rect 19524 18028 19576 18080
rect 21456 18028 21508 18080
rect 21824 18071 21876 18080
rect 21824 18037 21833 18071
rect 21833 18037 21867 18071
rect 21867 18037 21876 18071
rect 21824 18028 21876 18037
rect 22008 18071 22060 18080
rect 22008 18037 22017 18071
rect 22017 18037 22051 18071
rect 22051 18037 22060 18071
rect 22008 18028 22060 18037
rect 23296 18028 23348 18080
rect 23664 18071 23716 18080
rect 23664 18037 23673 18071
rect 23673 18037 23707 18071
rect 23707 18037 23716 18071
rect 23664 18028 23716 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1860 17824 1912 17876
rect 2320 17824 2372 17876
rect 3792 17867 3844 17876
rect 3792 17833 3801 17867
rect 3801 17833 3835 17867
rect 3835 17833 3844 17867
rect 3792 17824 3844 17833
rect 4988 17824 5040 17876
rect 5540 17824 5592 17876
rect 7104 17867 7156 17876
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 9588 17824 9640 17876
rect 10784 17867 10836 17876
rect 10784 17833 10793 17867
rect 10793 17833 10827 17867
rect 10827 17833 10836 17867
rect 10784 17824 10836 17833
rect 10876 17824 10928 17876
rect 11336 17867 11388 17876
rect 11336 17833 11345 17867
rect 11345 17833 11379 17867
rect 11379 17833 11388 17867
rect 11336 17824 11388 17833
rect 12808 17867 12860 17876
rect 12808 17833 12817 17867
rect 12817 17833 12851 17867
rect 12851 17833 12860 17867
rect 12808 17824 12860 17833
rect 13820 17867 13872 17876
rect 13820 17833 13829 17867
rect 13829 17833 13863 17867
rect 13863 17833 13872 17867
rect 13820 17824 13872 17833
rect 14556 17824 14608 17876
rect 19156 17867 19208 17876
rect 19156 17833 19165 17867
rect 19165 17833 19199 17867
rect 19199 17833 19208 17867
rect 19156 17824 19208 17833
rect 19984 17824 20036 17876
rect 22100 17824 22152 17876
rect 22468 17824 22520 17876
rect 2228 17756 2280 17808
rect 6920 17756 6972 17808
rect 7840 17756 7892 17808
rect 9312 17756 9364 17808
rect 13360 17799 13412 17808
rect 13360 17765 13369 17799
rect 13369 17765 13403 17799
rect 13403 17765 13412 17799
rect 13360 17756 13412 17765
rect 2964 17688 3016 17740
rect 3976 17688 4028 17740
rect 4068 17688 4120 17740
rect 6828 17688 6880 17740
rect 7564 17688 7616 17740
rect 9036 17731 9088 17740
rect 9036 17697 9045 17731
rect 9045 17697 9079 17731
rect 9079 17697 9088 17731
rect 9036 17688 9088 17697
rect 12164 17688 12216 17740
rect 15752 17731 15804 17740
rect 15752 17697 15761 17731
rect 15761 17697 15795 17731
rect 15795 17697 15804 17731
rect 15752 17688 15804 17697
rect 1492 17663 1544 17672
rect 1492 17629 1501 17663
rect 1501 17629 1535 17663
rect 1535 17629 1544 17663
rect 1492 17620 1544 17629
rect 17868 17756 17920 17808
rect 23664 17756 23716 17808
rect 17040 17688 17092 17740
rect 19432 17688 19484 17740
rect 21456 17688 21508 17740
rect 25872 17688 25924 17740
rect 7932 17663 7984 17672
rect 7932 17629 7941 17663
rect 7941 17629 7975 17663
rect 7975 17629 7984 17663
rect 7932 17620 7984 17629
rect 9404 17620 9456 17672
rect 10232 17620 10284 17672
rect 11336 17620 11388 17672
rect 6920 17552 6972 17604
rect 9680 17595 9732 17604
rect 9680 17561 9689 17595
rect 9689 17561 9723 17595
rect 9723 17561 9732 17595
rect 9680 17552 9732 17561
rect 2136 17484 2188 17536
rect 2596 17484 2648 17536
rect 4436 17484 4488 17536
rect 6184 17527 6236 17536
rect 6184 17493 6193 17527
rect 6193 17493 6227 17527
rect 6227 17493 6236 17527
rect 6184 17484 6236 17493
rect 7748 17484 7800 17536
rect 8484 17484 8536 17536
rect 9588 17484 9640 17536
rect 14832 17620 14884 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16028 17663 16080 17672
rect 16028 17629 16037 17663
rect 16037 17629 16071 17663
rect 16071 17629 16080 17663
rect 16028 17620 16080 17629
rect 15384 17595 15436 17604
rect 15384 17561 15393 17595
rect 15393 17561 15427 17595
rect 15427 17561 15436 17595
rect 15384 17552 15436 17561
rect 11796 17484 11848 17536
rect 16580 17484 16632 17536
rect 16948 17484 17000 17536
rect 18696 17484 18748 17536
rect 19248 17484 19300 17536
rect 20812 17620 20864 17672
rect 22928 17620 22980 17672
rect 24032 17663 24084 17672
rect 24032 17629 24041 17663
rect 24041 17629 24075 17663
rect 24075 17629 24084 17663
rect 24032 17620 24084 17629
rect 22192 17484 22244 17536
rect 23112 17484 23164 17536
rect 23388 17527 23440 17536
rect 23388 17493 23397 17527
rect 23397 17493 23431 17527
rect 23431 17493 23440 17527
rect 23388 17484 23440 17493
rect 24216 17484 24268 17536
rect 25136 17527 25188 17536
rect 25136 17493 25145 17527
rect 25145 17493 25179 17527
rect 25179 17493 25188 17527
rect 25136 17484 25188 17493
rect 25596 17527 25648 17536
rect 25596 17493 25605 17527
rect 25605 17493 25639 17527
rect 25639 17493 25648 17527
rect 25596 17484 25648 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1584 17280 1636 17332
rect 2780 17280 2832 17332
rect 3792 17280 3844 17332
rect 4068 17323 4120 17332
rect 4068 17289 4077 17323
rect 4077 17289 4111 17323
rect 4111 17289 4120 17323
rect 4068 17280 4120 17289
rect 4160 17280 4212 17332
rect 1492 17212 1544 17264
rect 1952 17212 2004 17264
rect 3976 17212 4028 17264
rect 4344 17255 4396 17264
rect 4344 17221 4353 17255
rect 4353 17221 4387 17255
rect 4387 17221 4396 17255
rect 4344 17212 4396 17221
rect 5448 17280 5500 17332
rect 7840 17323 7892 17332
rect 7840 17289 7849 17323
rect 7849 17289 7883 17323
rect 7883 17289 7892 17323
rect 7840 17280 7892 17289
rect 9680 17280 9732 17332
rect 9956 17280 10008 17332
rect 10232 17280 10284 17332
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 13268 17280 13320 17332
rect 13636 17323 13688 17332
rect 13636 17289 13645 17323
rect 13645 17289 13679 17323
rect 13679 17289 13688 17323
rect 13636 17280 13688 17289
rect 16028 17280 16080 17332
rect 16488 17280 16540 17332
rect 17040 17280 17092 17332
rect 6276 17212 6328 17264
rect 7932 17212 7984 17264
rect 9404 17255 9456 17264
rect 9404 17221 9413 17255
rect 9413 17221 9447 17255
rect 9447 17221 9456 17255
rect 9404 17212 9456 17221
rect 12716 17212 12768 17264
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5540 17187 5592 17196
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 11428 17187 11480 17196
rect 11428 17153 11437 17187
rect 11437 17153 11471 17187
rect 11471 17153 11480 17187
rect 11428 17144 11480 17153
rect 16948 17187 17000 17196
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 22376 17280 22428 17332
rect 23204 17280 23256 17332
rect 20812 17212 20864 17264
rect 23112 17212 23164 17264
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 22468 17187 22520 17196
rect 22468 17153 22477 17187
rect 22477 17153 22511 17187
rect 22511 17153 22520 17187
rect 22468 17144 22520 17153
rect 2320 17119 2372 17128
rect 2320 17085 2354 17119
rect 2354 17085 2372 17119
rect 2320 17076 2372 17085
rect 4988 17076 5040 17128
rect 1768 16940 1820 16992
rect 2596 16940 2648 16992
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 4896 16940 4948 16949
rect 6000 16983 6052 16992
rect 6000 16949 6009 16983
rect 6009 16949 6043 16983
rect 6043 16949 6052 16983
rect 6000 16940 6052 16949
rect 7748 17076 7800 17128
rect 10784 17076 10836 17128
rect 8484 17008 8536 17060
rect 10048 17008 10100 17060
rect 11336 17076 11388 17128
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 13820 17076 13872 17128
rect 15108 17076 15160 17128
rect 16764 17119 16816 17128
rect 16764 17085 16773 17119
rect 16773 17085 16807 17119
rect 16807 17085 16816 17119
rect 16764 17076 16816 17085
rect 22100 17076 22152 17128
rect 16580 17008 16632 17060
rect 21640 17008 21692 17060
rect 24032 17008 24084 17060
rect 7840 16940 7892 16992
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 14556 16940 14608 16992
rect 17868 16983 17920 16992
rect 17868 16949 17877 16983
rect 17877 16949 17911 16983
rect 17911 16949 17920 16983
rect 17868 16940 17920 16949
rect 18696 16940 18748 16992
rect 19524 16940 19576 16992
rect 21456 16940 21508 16992
rect 22928 16940 22980 16992
rect 25044 16983 25096 16992
rect 25044 16949 25053 16983
rect 25053 16949 25087 16983
rect 25087 16949 25096 16983
rect 25044 16940 25096 16949
rect 25872 16940 25924 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 1676 16736 1728 16788
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 2228 16779 2280 16788
rect 2228 16745 2237 16779
rect 2237 16745 2271 16779
rect 2271 16745 2280 16779
rect 2228 16736 2280 16745
rect 2872 16736 2924 16788
rect 3148 16736 3200 16788
rect 4252 16779 4304 16788
rect 2504 16668 2556 16720
rect 1952 16600 2004 16652
rect 2320 16600 2372 16652
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 4988 16779 5040 16788
rect 4988 16745 4997 16779
rect 4997 16745 5031 16779
rect 5031 16745 5040 16779
rect 4988 16736 5040 16745
rect 5172 16736 5224 16788
rect 6828 16779 6880 16788
rect 5540 16668 5592 16720
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 7564 16736 7616 16788
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 8208 16736 8260 16788
rect 8392 16779 8444 16788
rect 8392 16745 8401 16779
rect 8401 16745 8435 16779
rect 8435 16745 8444 16779
rect 8392 16736 8444 16745
rect 11428 16736 11480 16788
rect 12900 16736 12952 16788
rect 13820 16779 13872 16788
rect 13820 16745 13829 16779
rect 13829 16745 13863 16779
rect 13863 16745 13872 16779
rect 13820 16736 13872 16745
rect 15292 16779 15344 16788
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 16948 16736 17000 16788
rect 17868 16736 17920 16788
rect 18696 16779 18748 16788
rect 18696 16745 18705 16779
rect 18705 16745 18739 16779
rect 18739 16745 18748 16779
rect 18696 16736 18748 16745
rect 18880 16779 18932 16788
rect 18880 16745 18889 16779
rect 18889 16745 18923 16779
rect 18923 16745 18932 16779
rect 18880 16736 18932 16745
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 19340 16779 19392 16788
rect 19340 16745 19349 16779
rect 19349 16745 19383 16779
rect 19383 16745 19392 16779
rect 20720 16779 20772 16788
rect 19340 16736 19392 16745
rect 20720 16745 20729 16779
rect 20729 16745 20763 16779
rect 20763 16745 20772 16779
rect 20720 16736 20772 16745
rect 20812 16736 20864 16788
rect 21640 16736 21692 16788
rect 22100 16736 22152 16788
rect 22928 16779 22980 16788
rect 22928 16745 22937 16779
rect 22937 16745 22971 16779
rect 22971 16745 22980 16779
rect 22928 16736 22980 16745
rect 24400 16779 24452 16788
rect 24400 16745 24409 16779
rect 24409 16745 24443 16779
rect 24443 16745 24452 16779
rect 24400 16736 24452 16745
rect 3056 16575 3108 16584
rect 1768 16464 1820 16516
rect 2596 16464 2648 16516
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 4344 16600 4396 16652
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 7564 16600 7616 16652
rect 9312 16668 9364 16720
rect 23296 16711 23348 16720
rect 9036 16600 9088 16652
rect 3056 16532 3108 16541
rect 3700 16464 3752 16516
rect 5172 16532 5224 16584
rect 8852 16532 8904 16584
rect 9496 16532 9548 16584
rect 23296 16677 23330 16711
rect 23330 16677 23348 16711
rect 23296 16668 23348 16677
rect 10968 16600 11020 16652
rect 11336 16600 11388 16652
rect 10140 16532 10192 16584
rect 10876 16532 10928 16584
rect 3976 16464 4028 16516
rect 4252 16464 4304 16516
rect 9588 16464 9640 16516
rect 10968 16464 11020 16516
rect 12992 16532 13044 16584
rect 14372 16643 14424 16652
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 17040 16600 17092 16652
rect 19432 16600 19484 16652
rect 20168 16600 20220 16652
rect 20444 16600 20496 16652
rect 16212 16532 16264 16584
rect 19524 16575 19576 16584
rect 19524 16541 19533 16575
rect 19533 16541 19567 16575
rect 19567 16541 19576 16575
rect 19524 16532 19576 16541
rect 19984 16532 20036 16584
rect 20720 16600 20772 16652
rect 23112 16600 23164 16652
rect 21364 16575 21416 16584
rect 21364 16541 21373 16575
rect 21373 16541 21407 16575
rect 21407 16541 21416 16575
rect 21364 16532 21416 16541
rect 21916 16532 21968 16584
rect 2228 16396 2280 16448
rect 2504 16396 2556 16448
rect 11060 16396 11112 16448
rect 11704 16396 11756 16448
rect 18420 16439 18472 16448
rect 18420 16405 18429 16439
rect 18429 16405 18463 16439
rect 18463 16405 18472 16439
rect 18420 16396 18472 16405
rect 20444 16396 20496 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1676 16192 1728 16244
rect 5172 16235 5224 16244
rect 5172 16201 5181 16235
rect 5181 16201 5215 16235
rect 5215 16201 5224 16235
rect 5172 16192 5224 16201
rect 5448 16192 5500 16244
rect 5080 16167 5132 16176
rect 5080 16133 5089 16167
rect 5089 16133 5123 16167
rect 5123 16133 5132 16167
rect 5080 16124 5132 16133
rect 5908 16124 5960 16176
rect 4712 16099 4764 16108
rect 4712 16065 4721 16099
rect 4721 16065 4755 16099
rect 4755 16065 4764 16099
rect 4712 16056 4764 16065
rect 5540 16056 5592 16108
rect 7748 16192 7800 16244
rect 9312 16235 9364 16244
rect 9312 16201 9321 16235
rect 9321 16201 9355 16235
rect 9355 16201 9364 16235
rect 9312 16192 9364 16201
rect 10140 16192 10192 16244
rect 10968 16192 11020 16244
rect 11796 16235 11848 16244
rect 11796 16201 11805 16235
rect 11805 16201 11839 16235
rect 11839 16201 11848 16235
rect 11796 16192 11848 16201
rect 14004 16235 14056 16244
rect 14004 16201 14013 16235
rect 14013 16201 14047 16235
rect 14047 16201 14056 16235
rect 14004 16192 14056 16201
rect 14832 16192 14884 16244
rect 11060 16124 11112 16176
rect 12808 16124 12860 16176
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 1584 15895 1636 15904
rect 1584 15861 1593 15895
rect 1593 15861 1627 15895
rect 1627 15861 1636 15895
rect 1584 15852 1636 15861
rect 4344 15988 4396 16040
rect 6000 15988 6052 16040
rect 9312 15988 9364 16040
rect 13820 16031 13872 16040
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 14372 16031 14424 16040
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 15752 16192 15804 16244
rect 18052 16235 18104 16244
rect 18052 16201 18061 16235
rect 18061 16201 18095 16235
rect 18095 16201 18104 16235
rect 18052 16192 18104 16201
rect 19340 16192 19392 16244
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 21364 16192 21416 16244
rect 22008 16192 22060 16244
rect 23112 16235 23164 16244
rect 23112 16201 23121 16235
rect 23121 16201 23155 16235
rect 23155 16201 23164 16235
rect 23112 16192 23164 16201
rect 21916 16124 21968 16176
rect 23296 16124 23348 16176
rect 17040 16099 17092 16108
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 18420 16056 18472 16108
rect 21456 16056 21508 16108
rect 18696 15988 18748 16040
rect 20628 15988 20680 16040
rect 21732 15988 21784 16040
rect 3332 15920 3384 15972
rect 3976 15895 4028 15904
rect 3976 15861 3985 15895
rect 3985 15861 4019 15895
rect 4019 15861 4028 15895
rect 3976 15852 4028 15861
rect 5080 15920 5132 15972
rect 7012 15920 7064 15972
rect 11060 15920 11112 15972
rect 12992 15920 13044 15972
rect 7196 15852 7248 15904
rect 7748 15852 7800 15904
rect 9036 15852 9088 15904
rect 11520 15852 11572 15904
rect 12440 15895 12492 15904
rect 12440 15861 12449 15895
rect 12449 15861 12483 15895
rect 12483 15861 12492 15895
rect 12440 15852 12492 15861
rect 13360 15852 13412 15904
rect 14096 15852 14148 15904
rect 14372 15852 14424 15904
rect 14464 15895 14516 15904
rect 14464 15861 14473 15895
rect 14473 15861 14507 15895
rect 14507 15861 14516 15895
rect 14464 15852 14516 15861
rect 16212 15852 16264 15904
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 17684 15852 17736 15904
rect 18880 15920 18932 15972
rect 19524 15920 19576 15972
rect 20536 15920 20588 15972
rect 21272 15920 21324 15972
rect 23480 15920 23532 15972
rect 24216 15920 24268 15972
rect 18604 15852 18656 15904
rect 20444 15895 20496 15904
rect 20444 15861 20453 15895
rect 20453 15861 20487 15895
rect 20487 15861 20496 15895
rect 20444 15852 20496 15861
rect 24032 15852 24084 15904
rect 25228 15852 25280 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1860 15691 1912 15700
rect 1860 15657 1869 15691
rect 1869 15657 1903 15691
rect 1903 15657 1912 15691
rect 1860 15648 1912 15657
rect 2044 15648 2096 15700
rect 3056 15648 3108 15700
rect 3332 15691 3384 15700
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 4344 15691 4396 15700
rect 4344 15657 4353 15691
rect 4353 15657 4387 15691
rect 4387 15657 4396 15691
rect 4344 15648 4396 15657
rect 4804 15648 4856 15700
rect 5540 15691 5592 15700
rect 5540 15657 5549 15691
rect 5549 15657 5583 15691
rect 5583 15657 5592 15691
rect 5540 15648 5592 15657
rect 8208 15648 8260 15700
rect 8668 15648 8720 15700
rect 9496 15691 9548 15700
rect 9496 15657 9505 15691
rect 9505 15657 9539 15691
rect 9539 15657 9548 15691
rect 9496 15648 9548 15657
rect 9772 15648 9824 15700
rect 9956 15648 10008 15700
rect 10876 15691 10928 15700
rect 10876 15657 10885 15691
rect 10885 15657 10919 15691
rect 10919 15657 10928 15691
rect 10876 15648 10928 15657
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 12808 15691 12860 15700
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 17040 15648 17092 15700
rect 18420 15648 18472 15700
rect 18512 15691 18564 15700
rect 18512 15657 18521 15691
rect 18521 15657 18555 15691
rect 18555 15657 18564 15691
rect 19340 15691 19392 15700
rect 18512 15648 18564 15657
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 21272 15648 21324 15700
rect 21732 15648 21784 15700
rect 22468 15648 22520 15700
rect 22928 15691 22980 15700
rect 22928 15657 22937 15691
rect 22937 15657 22971 15691
rect 22971 15657 22980 15691
rect 23480 15691 23532 15700
rect 22928 15648 22980 15657
rect 23480 15657 23489 15691
rect 23489 15657 23523 15691
rect 23523 15657 23532 15691
rect 23480 15648 23532 15657
rect 23848 15691 23900 15700
rect 23848 15657 23857 15691
rect 23857 15657 23891 15691
rect 23891 15657 23900 15691
rect 23848 15648 23900 15657
rect 4528 15580 4580 15632
rect 6276 15580 6328 15632
rect 8852 15580 8904 15632
rect 11704 15623 11756 15632
rect 11704 15589 11738 15623
rect 11738 15589 11756 15623
rect 11704 15580 11756 15589
rect 12440 15580 12492 15632
rect 2044 15512 2096 15564
rect 2320 15555 2372 15564
rect 2320 15521 2329 15555
rect 2329 15521 2363 15555
rect 2363 15521 2372 15555
rect 3700 15555 3752 15564
rect 2320 15512 2372 15521
rect 3700 15521 3709 15555
rect 3709 15521 3743 15555
rect 3743 15521 3752 15555
rect 3700 15512 3752 15521
rect 4988 15512 5040 15564
rect 5908 15555 5960 15564
rect 5908 15521 5917 15555
rect 5917 15521 5951 15555
rect 5951 15521 5960 15555
rect 5908 15512 5960 15521
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 9312 15512 9364 15564
rect 10968 15512 11020 15564
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 3608 15444 3660 15496
rect 4344 15444 4396 15496
rect 5448 15444 5500 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 9496 15376 9548 15428
rect 10784 15444 10836 15496
rect 13268 15512 13320 15564
rect 14004 15512 14056 15564
rect 16764 15555 16816 15564
rect 16764 15521 16798 15555
rect 16798 15521 16816 15555
rect 16764 15512 16816 15521
rect 21088 15512 21140 15564
rect 23848 15512 23900 15564
rect 24768 15512 24820 15564
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 16212 15444 16264 15496
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 14096 15419 14148 15428
rect 14096 15385 14105 15419
rect 14105 15385 14139 15419
rect 14139 15385 14148 15419
rect 14096 15376 14148 15385
rect 19248 15376 19300 15428
rect 21364 15444 21416 15496
rect 25228 15444 25280 15496
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 13820 15308 13872 15360
rect 14464 15308 14516 15360
rect 18972 15351 19024 15360
rect 18972 15317 18981 15351
rect 18981 15317 19015 15351
rect 19015 15317 19024 15351
rect 18972 15308 19024 15317
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 24032 15351 24084 15360
rect 24032 15317 24041 15351
rect 24041 15317 24075 15351
rect 24075 15317 24084 15351
rect 24032 15308 24084 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 4804 15104 4856 15156
rect 6000 15104 6052 15156
rect 2320 15036 2372 15088
rect 6276 15104 6328 15156
rect 7012 15147 7064 15156
rect 7012 15113 7021 15147
rect 7021 15113 7055 15147
rect 7055 15113 7064 15147
rect 7012 15104 7064 15113
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 10784 15147 10836 15156
rect 10784 15113 10793 15147
rect 10793 15113 10827 15147
rect 10827 15113 10836 15147
rect 10784 15104 10836 15113
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 12532 15104 12584 15156
rect 12716 15147 12768 15156
rect 12716 15113 12725 15147
rect 12725 15113 12759 15147
rect 12759 15113 12768 15147
rect 12716 15104 12768 15113
rect 16764 15104 16816 15156
rect 17592 15104 17644 15156
rect 2504 15011 2556 15020
rect 2504 14977 2513 15011
rect 2513 14977 2547 15011
rect 2547 14977 2556 15011
rect 2504 14968 2556 14977
rect 2412 14900 2464 14952
rect 3976 14968 4028 15020
rect 4988 14968 5040 15020
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 5172 14900 5224 14952
rect 4620 14832 4672 14884
rect 4988 14832 5040 14884
rect 5264 14832 5316 14884
rect 6828 14900 6880 14952
rect 11060 14968 11112 15020
rect 11704 14968 11756 15020
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 19064 15104 19116 15156
rect 19340 15104 19392 15156
rect 21088 15104 21140 15156
rect 22100 15104 22152 15156
rect 22652 15147 22704 15156
rect 22652 15113 22661 15147
rect 22661 15113 22695 15147
rect 22695 15113 22704 15147
rect 22652 15104 22704 15113
rect 23480 15147 23532 15156
rect 23480 15113 23489 15147
rect 23489 15113 23523 15147
rect 23523 15113 23532 15147
rect 23480 15104 23532 15113
rect 23848 15147 23900 15156
rect 23848 15113 23857 15147
rect 23857 15113 23891 15147
rect 23891 15113 23900 15147
rect 23848 15104 23900 15113
rect 24676 15104 24728 15156
rect 24216 15036 24268 15088
rect 25228 15079 25280 15088
rect 25228 15045 25237 15079
rect 25237 15045 25271 15079
rect 25271 15045 25280 15079
rect 25228 15036 25280 15045
rect 8852 14900 8904 14952
rect 7840 14832 7892 14884
rect 13176 14875 13228 14884
rect 13176 14841 13185 14875
rect 13185 14841 13219 14875
rect 13219 14841 13228 14875
rect 13176 14832 13228 14841
rect 13452 14832 13504 14884
rect 16212 14900 16264 14952
rect 18236 14900 18288 14952
rect 18972 14900 19024 14952
rect 14556 14832 14608 14884
rect 18696 14832 18748 14884
rect 19064 14875 19116 14884
rect 19064 14841 19073 14875
rect 19073 14841 19107 14875
rect 19107 14841 19116 14875
rect 19064 14832 19116 14841
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 2504 14764 2556 14816
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 4068 14807 4120 14816
rect 4068 14773 4077 14807
rect 4077 14773 4111 14807
rect 4111 14773 4120 14807
rect 4068 14764 4120 14773
rect 5080 14764 5132 14816
rect 6368 14764 6420 14816
rect 6552 14764 6604 14816
rect 9220 14764 9272 14816
rect 10140 14764 10192 14816
rect 12716 14764 12768 14816
rect 14004 14807 14056 14816
rect 14004 14773 14013 14807
rect 14013 14773 14047 14807
rect 14047 14773 14056 14807
rect 14004 14764 14056 14773
rect 16396 14764 16448 14816
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 18328 14764 18380 14816
rect 21272 14900 21324 14952
rect 23940 14900 23992 14952
rect 24400 15011 24452 15020
rect 24400 14977 24409 15011
rect 24409 14977 24443 15011
rect 24443 14977 24452 15011
rect 24400 14968 24452 14977
rect 19984 14832 20036 14884
rect 20904 14764 20956 14816
rect 21364 14764 21416 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2136 14560 2188 14612
rect 2596 14560 2648 14612
rect 3976 14560 4028 14612
rect 4160 14560 4212 14612
rect 6276 14603 6328 14612
rect 6276 14569 6285 14603
rect 6285 14569 6319 14603
rect 6319 14569 6328 14603
rect 6276 14560 6328 14569
rect 7012 14560 7064 14612
rect 9496 14603 9548 14612
rect 9496 14569 9505 14603
rect 9505 14569 9539 14603
rect 9539 14569 9548 14603
rect 9496 14560 9548 14569
rect 11704 14603 11756 14612
rect 11704 14569 11713 14603
rect 11713 14569 11747 14603
rect 11747 14569 11756 14603
rect 11704 14560 11756 14569
rect 12348 14603 12400 14612
rect 12348 14569 12357 14603
rect 12357 14569 12391 14603
rect 12391 14569 12400 14603
rect 12348 14560 12400 14569
rect 13268 14560 13320 14612
rect 13820 14560 13872 14612
rect 17592 14603 17644 14612
rect 17592 14569 17601 14603
rect 17601 14569 17635 14603
rect 17635 14569 17644 14603
rect 17592 14560 17644 14569
rect 18236 14603 18288 14612
rect 18236 14569 18245 14603
rect 18245 14569 18279 14603
rect 18279 14569 18288 14603
rect 18236 14560 18288 14569
rect 18696 14603 18748 14612
rect 18696 14569 18705 14603
rect 18705 14569 18739 14603
rect 18739 14569 18748 14603
rect 18696 14560 18748 14569
rect 20720 14603 20772 14612
rect 20720 14569 20729 14603
rect 20729 14569 20763 14603
rect 20763 14569 20772 14603
rect 20720 14560 20772 14569
rect 24768 14560 24820 14612
rect 25688 14560 25740 14612
rect 4344 14535 4396 14544
rect 4344 14501 4353 14535
rect 4353 14501 4387 14535
rect 4387 14501 4396 14535
rect 4344 14492 4396 14501
rect 3148 14424 3200 14476
rect 4620 14424 4672 14476
rect 5080 14424 5132 14476
rect 6276 14424 6328 14476
rect 7288 14424 7340 14476
rect 8760 14424 8812 14476
rect 11520 14424 11572 14476
rect 12072 14424 12124 14476
rect 13360 14424 13412 14476
rect 14464 14424 14516 14476
rect 16212 14467 16264 14476
rect 16212 14433 16221 14467
rect 16221 14433 16255 14467
rect 16255 14433 16264 14467
rect 16212 14424 16264 14433
rect 16488 14467 16540 14476
rect 16488 14433 16522 14467
rect 16522 14433 16540 14467
rect 16488 14424 16540 14433
rect 19064 14467 19116 14476
rect 19064 14433 19073 14467
rect 19073 14433 19107 14467
rect 19107 14433 19116 14467
rect 19064 14424 19116 14433
rect 2412 14356 2464 14408
rect 3608 14356 3660 14408
rect 1768 14288 1820 14340
rect 5080 14288 5132 14340
rect 5540 14356 5592 14408
rect 6000 14356 6052 14408
rect 6368 14356 6420 14408
rect 8852 14356 8904 14408
rect 12992 14356 13044 14408
rect 13728 14356 13780 14408
rect 14188 14399 14240 14408
rect 14188 14365 14197 14399
rect 14197 14365 14231 14399
rect 14231 14365 14240 14399
rect 14188 14356 14240 14365
rect 18420 14356 18472 14408
rect 19524 14492 19576 14544
rect 21088 14492 21140 14544
rect 23664 14492 23716 14544
rect 22284 14424 22336 14476
rect 23848 14424 23900 14476
rect 25136 14424 25188 14476
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 20904 14399 20956 14408
rect 19248 14356 19300 14365
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 23480 14356 23532 14408
rect 24308 14399 24360 14408
rect 24308 14365 24317 14399
rect 24317 14365 24351 14399
rect 24351 14365 24360 14399
rect 24308 14356 24360 14365
rect 24400 14399 24452 14408
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 5816 14288 5868 14340
rect 6276 14288 6328 14340
rect 7840 14331 7892 14340
rect 7840 14297 7849 14331
rect 7849 14297 7883 14331
rect 7883 14297 7892 14331
rect 7840 14288 7892 14297
rect 22284 14331 22336 14340
rect 22284 14297 22293 14331
rect 22293 14297 22327 14331
rect 22327 14297 22336 14331
rect 22284 14288 22336 14297
rect 1676 14220 1728 14272
rect 2504 14220 2556 14272
rect 6092 14220 6144 14272
rect 7104 14220 7156 14272
rect 9128 14263 9180 14272
rect 9128 14229 9137 14263
rect 9137 14229 9171 14263
rect 9171 14229 9180 14263
rect 9128 14220 9180 14229
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 12716 14263 12768 14272
rect 12716 14229 12725 14263
rect 12725 14229 12759 14263
rect 12759 14229 12768 14263
rect 12716 14220 12768 14229
rect 13452 14263 13504 14272
rect 13452 14229 13461 14263
rect 13461 14229 13495 14263
rect 13495 14229 13504 14263
rect 13452 14220 13504 14229
rect 14556 14220 14608 14272
rect 16028 14263 16080 14272
rect 16028 14229 16037 14263
rect 16037 14229 16071 14263
rect 16071 14229 16080 14263
rect 16028 14220 16080 14229
rect 18696 14220 18748 14272
rect 19708 14263 19760 14272
rect 19708 14229 19717 14263
rect 19717 14229 19751 14263
rect 19751 14229 19760 14263
rect 19708 14220 19760 14229
rect 23112 14220 23164 14272
rect 23756 14263 23808 14272
rect 23756 14229 23765 14263
rect 23765 14229 23799 14263
rect 23799 14229 23808 14263
rect 23756 14220 23808 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 2688 14059 2740 14068
rect 2688 14025 2697 14059
rect 2697 14025 2731 14059
rect 2731 14025 2740 14059
rect 2688 14016 2740 14025
rect 6368 14016 6420 14068
rect 7380 14016 7432 14068
rect 8484 14016 8536 14068
rect 8852 14016 8904 14068
rect 11520 14059 11572 14068
rect 11520 14025 11529 14059
rect 11529 14025 11563 14059
rect 11563 14025 11572 14059
rect 11520 14016 11572 14025
rect 12992 14059 13044 14068
rect 12992 14025 13001 14059
rect 13001 14025 13035 14059
rect 13035 14025 13044 14059
rect 12992 14016 13044 14025
rect 13360 14059 13412 14068
rect 13360 14025 13369 14059
rect 13369 14025 13403 14059
rect 13403 14025 13412 14059
rect 13360 14016 13412 14025
rect 16488 14016 16540 14068
rect 19248 14016 19300 14068
rect 21272 14059 21324 14068
rect 21272 14025 21281 14059
rect 21281 14025 21315 14059
rect 21315 14025 21324 14059
rect 21272 14016 21324 14025
rect 23112 14016 23164 14068
rect 23480 14059 23532 14068
rect 23480 14025 23489 14059
rect 23489 14025 23523 14059
rect 23523 14025 23532 14059
rect 23480 14016 23532 14025
rect 2596 13948 2648 14000
rect 5172 13991 5224 14000
rect 5172 13957 5181 13991
rect 5181 13957 5215 13991
rect 5215 13957 5224 13991
rect 5172 13948 5224 13957
rect 8208 13948 8260 14000
rect 14556 13948 14608 14000
rect 16212 13948 16264 14000
rect 16856 13948 16908 14000
rect 19984 13991 20036 14000
rect 19984 13957 19993 13991
rect 19993 13957 20027 13991
rect 20027 13957 20036 13991
rect 19984 13948 20036 13957
rect 1676 13880 1728 13932
rect 2688 13880 2740 13932
rect 3884 13880 3936 13932
rect 6184 13880 6236 13932
rect 8116 13880 8168 13932
rect 8760 13880 8812 13932
rect 9128 13880 9180 13932
rect 7840 13855 7892 13864
rect 3516 13744 3568 13796
rect 3884 13744 3936 13796
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 8484 13855 8536 13864
rect 7840 13812 7892 13821
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 16028 13880 16080 13932
rect 20904 13923 20956 13932
rect 10140 13812 10192 13864
rect 11060 13812 11112 13864
rect 12532 13812 12584 13864
rect 13452 13855 13504 13864
rect 13452 13821 13461 13855
rect 13461 13821 13495 13855
rect 13495 13821 13504 13855
rect 13452 13812 13504 13821
rect 15384 13855 15436 13864
rect 15384 13821 15393 13855
rect 15393 13821 15427 13855
rect 15427 13821 15436 13855
rect 15384 13812 15436 13821
rect 18328 13812 18380 13864
rect 20904 13889 20913 13923
rect 20913 13889 20947 13923
rect 20947 13889 20956 13923
rect 20904 13880 20956 13889
rect 22928 13948 22980 14000
rect 22836 13880 22888 13932
rect 23388 13880 23440 13932
rect 23756 13880 23808 13932
rect 25136 13880 25188 13932
rect 9956 13744 10008 13796
rect 12164 13787 12216 13796
rect 12164 13753 12173 13787
rect 12173 13753 12207 13787
rect 12207 13753 12216 13787
rect 12164 13744 12216 13753
rect 13820 13744 13872 13796
rect 18420 13787 18472 13796
rect 3608 13719 3660 13728
rect 3608 13685 3617 13719
rect 3617 13685 3651 13719
rect 3651 13685 3660 13719
rect 3608 13676 3660 13685
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 4988 13719 5040 13728
rect 4988 13685 4997 13719
rect 4997 13685 5031 13719
rect 5031 13685 5040 13719
rect 4988 13676 5040 13685
rect 10968 13719 11020 13728
rect 10968 13685 10977 13719
rect 10977 13685 11011 13719
rect 11011 13685 11020 13719
rect 10968 13676 11020 13685
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 12716 13676 12768 13728
rect 18420 13753 18429 13787
rect 18429 13753 18463 13787
rect 18463 13753 18472 13787
rect 18420 13744 18472 13753
rect 18696 13744 18748 13796
rect 23112 13812 23164 13864
rect 24308 13812 24360 13864
rect 25228 13855 25280 13864
rect 25228 13821 25237 13855
rect 25237 13821 25271 13855
rect 25271 13821 25280 13855
rect 25228 13812 25280 13821
rect 15936 13719 15988 13728
rect 15936 13685 15945 13719
rect 15945 13685 15979 13719
rect 15979 13685 15988 13719
rect 15936 13676 15988 13685
rect 16304 13719 16356 13728
rect 16304 13685 16313 13719
rect 16313 13685 16347 13719
rect 16347 13685 16356 13719
rect 16304 13676 16356 13685
rect 22100 13676 22152 13728
rect 22468 13719 22520 13728
rect 22468 13685 22477 13719
rect 22477 13685 22511 13719
rect 22511 13685 22520 13719
rect 22468 13676 22520 13685
rect 23664 13676 23716 13728
rect 25412 13719 25464 13728
rect 25412 13685 25421 13719
rect 25421 13685 25455 13719
rect 25455 13685 25464 13719
rect 25412 13676 25464 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 1952 13515 2004 13524
rect 1952 13481 1961 13515
rect 1961 13481 1995 13515
rect 1995 13481 2004 13515
rect 1952 13472 2004 13481
rect 2320 13515 2372 13524
rect 2320 13481 2329 13515
rect 2329 13481 2363 13515
rect 2363 13481 2372 13515
rect 2320 13472 2372 13481
rect 2872 13472 2924 13524
rect 3884 13472 3936 13524
rect 3976 13472 4028 13524
rect 4896 13515 4948 13524
rect 4896 13481 4905 13515
rect 4905 13481 4939 13515
rect 4939 13481 4948 13515
rect 4896 13472 4948 13481
rect 6460 13515 6512 13524
rect 6460 13481 6469 13515
rect 6469 13481 6503 13515
rect 6503 13481 6512 13515
rect 6460 13472 6512 13481
rect 8116 13472 8168 13524
rect 8484 13515 8536 13524
rect 8484 13481 8493 13515
rect 8493 13481 8527 13515
rect 8527 13481 8536 13515
rect 8484 13472 8536 13481
rect 13820 13515 13872 13524
rect 13820 13481 13829 13515
rect 13829 13481 13863 13515
rect 13863 13481 13872 13515
rect 13820 13472 13872 13481
rect 14188 13472 14240 13524
rect 18328 13472 18380 13524
rect 21088 13515 21140 13524
rect 21088 13481 21097 13515
rect 21097 13481 21131 13515
rect 21131 13481 21140 13515
rect 21088 13472 21140 13481
rect 23388 13472 23440 13524
rect 23756 13515 23808 13524
rect 23756 13481 23765 13515
rect 23765 13481 23799 13515
rect 23799 13481 23808 13515
rect 23756 13472 23808 13481
rect 24032 13472 24084 13524
rect 25780 13472 25832 13524
rect 6184 13404 6236 13456
rect 8300 13404 8352 13456
rect 9588 13404 9640 13456
rect 12900 13404 12952 13456
rect 16396 13404 16448 13456
rect 23296 13404 23348 13456
rect 25044 13404 25096 13456
rect 2320 13336 2372 13388
rect 3056 13336 3108 13388
rect 4804 13379 4856 13388
rect 4804 13345 4813 13379
rect 4813 13345 4847 13379
rect 4847 13345 4856 13379
rect 4804 13336 4856 13345
rect 5632 13336 5684 13388
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 8760 13336 8812 13388
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 10968 13336 11020 13388
rect 12532 13336 12584 13388
rect 16856 13336 16908 13388
rect 20628 13336 20680 13388
rect 20904 13336 20956 13388
rect 22468 13336 22520 13388
rect 25320 13336 25372 13388
rect 4252 13268 4304 13320
rect 6092 13268 6144 13320
rect 6276 13268 6328 13320
rect 2228 13200 2280 13252
rect 8024 13243 8076 13252
rect 8024 13209 8033 13243
rect 8033 13209 8067 13243
rect 8067 13209 8076 13243
rect 8024 13200 8076 13209
rect 8116 13200 8168 13252
rect 9404 13268 9456 13320
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 19064 13311 19116 13320
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 19800 13311 19852 13320
rect 19800 13277 19809 13311
rect 19809 13277 19843 13311
rect 19843 13277 19852 13311
rect 19800 13268 19852 13277
rect 23848 13268 23900 13320
rect 24124 13268 24176 13320
rect 3148 13175 3200 13184
rect 3148 13141 3157 13175
rect 3157 13141 3191 13175
rect 3191 13141 3200 13175
rect 3148 13132 3200 13141
rect 5080 13132 5132 13184
rect 11428 13132 11480 13184
rect 12072 13132 12124 13184
rect 15476 13175 15528 13184
rect 15476 13141 15485 13175
rect 15485 13141 15519 13175
rect 15519 13141 15528 13175
rect 15476 13132 15528 13141
rect 16304 13175 16356 13184
rect 16304 13141 16313 13175
rect 16313 13141 16347 13175
rect 16347 13141 16356 13175
rect 16304 13132 16356 13141
rect 18604 13132 18656 13184
rect 19248 13175 19300 13184
rect 19248 13141 19257 13175
rect 19257 13141 19291 13175
rect 19291 13141 19300 13175
rect 19248 13132 19300 13141
rect 20352 13175 20404 13184
rect 20352 13141 20361 13175
rect 20361 13141 20395 13175
rect 20395 13141 20404 13175
rect 20352 13132 20404 13141
rect 23388 13175 23440 13184
rect 23388 13141 23397 13175
rect 23397 13141 23431 13175
rect 23431 13141 23440 13175
rect 23388 13132 23440 13141
rect 23848 13175 23900 13184
rect 23848 13141 23857 13175
rect 23857 13141 23891 13175
rect 23891 13141 23900 13175
rect 23848 13132 23900 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1492 12928 1544 12980
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 3608 12928 3660 12980
rect 4252 12971 4304 12980
rect 4252 12937 4261 12971
rect 4261 12937 4295 12971
rect 4295 12937 4304 12971
rect 4252 12928 4304 12937
rect 4712 12971 4764 12980
rect 4712 12937 4721 12971
rect 4721 12937 4755 12971
rect 4755 12937 4764 12971
rect 4712 12928 4764 12937
rect 4804 12928 4856 12980
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 6368 12928 6420 12980
rect 6828 12971 6880 12980
rect 6828 12937 6837 12971
rect 6837 12937 6871 12971
rect 6871 12937 6880 12971
rect 6828 12928 6880 12937
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 9956 12928 10008 12980
rect 10968 12928 11020 12980
rect 13544 12971 13596 12980
rect 13544 12937 13553 12971
rect 13553 12937 13587 12971
rect 13587 12937 13596 12971
rect 13544 12928 13596 12937
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 14832 12860 14884 12912
rect 5724 12792 5776 12801
rect 3608 12767 3660 12776
rect 3608 12733 3617 12767
rect 3617 12733 3651 12767
rect 3651 12733 3660 12767
rect 3608 12724 3660 12733
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 6644 12724 6696 12776
rect 9588 12792 9640 12844
rect 13728 12792 13780 12844
rect 14464 12792 14516 12844
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 17132 12971 17184 12980
rect 17132 12937 17141 12971
rect 17141 12937 17175 12971
rect 17175 12937 17184 12971
rect 17132 12928 17184 12937
rect 18052 12971 18104 12980
rect 18052 12937 18061 12971
rect 18061 12937 18095 12971
rect 18095 12937 18104 12971
rect 18052 12928 18104 12937
rect 19432 12928 19484 12980
rect 19800 12928 19852 12980
rect 20444 12928 20496 12980
rect 20904 12928 20956 12980
rect 21916 12971 21968 12980
rect 21916 12937 21925 12971
rect 21925 12937 21959 12971
rect 21959 12937 21968 12971
rect 21916 12928 21968 12937
rect 18328 12860 18380 12912
rect 20536 12860 20588 12912
rect 7656 12724 7708 12776
rect 4712 12656 4764 12708
rect 5724 12656 5776 12708
rect 7288 12699 7340 12708
rect 7288 12665 7297 12699
rect 7297 12665 7331 12699
rect 7331 12665 7340 12699
rect 7288 12656 7340 12665
rect 7932 12656 7984 12708
rect 2136 12588 2188 12640
rect 2688 12631 2740 12640
rect 2688 12597 2697 12631
rect 2697 12597 2731 12631
rect 2731 12597 2740 12631
rect 2688 12588 2740 12597
rect 3424 12588 3476 12640
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 8852 12588 8904 12640
rect 9036 12724 9088 12776
rect 9680 12724 9732 12776
rect 10048 12724 10100 12776
rect 13452 12767 13504 12776
rect 13452 12733 13461 12767
rect 13461 12733 13495 12767
rect 13495 12733 13504 12767
rect 14004 12767 14056 12776
rect 13452 12724 13504 12733
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 15476 12767 15528 12776
rect 15476 12733 15485 12767
rect 15485 12733 15519 12767
rect 15519 12733 15528 12767
rect 15476 12724 15528 12733
rect 16488 12792 16540 12844
rect 18420 12792 18472 12844
rect 23388 12928 23440 12980
rect 24124 12928 24176 12980
rect 25044 12971 25096 12980
rect 25044 12937 25053 12971
rect 25053 12937 25087 12971
rect 25087 12937 25096 12971
rect 25044 12928 25096 12937
rect 23480 12903 23532 12912
rect 23480 12869 23489 12903
rect 23489 12869 23523 12903
rect 23523 12869 23532 12903
rect 23480 12860 23532 12869
rect 24032 12860 24084 12912
rect 24400 12860 24452 12912
rect 25320 12860 25372 12912
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 22560 12792 22612 12801
rect 23112 12835 23164 12844
rect 23112 12801 23121 12835
rect 23121 12801 23155 12835
rect 23155 12801 23164 12835
rect 23112 12792 23164 12801
rect 24308 12792 24360 12844
rect 24676 12792 24728 12844
rect 15936 12724 15988 12776
rect 16212 12724 16264 12776
rect 16948 12767 17000 12776
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 18236 12724 18288 12776
rect 19156 12724 19208 12776
rect 19340 12724 19392 12776
rect 22192 12724 22244 12776
rect 23480 12724 23532 12776
rect 25044 12724 25096 12776
rect 9496 12656 9548 12708
rect 11612 12656 11664 12708
rect 13544 12656 13596 12708
rect 14188 12656 14240 12708
rect 15660 12656 15712 12708
rect 16120 12656 16172 12708
rect 19524 12656 19576 12708
rect 20444 12656 20496 12708
rect 21548 12656 21600 12708
rect 22468 12656 22520 12708
rect 23940 12656 23992 12708
rect 24308 12656 24360 12708
rect 9036 12588 9088 12640
rect 9772 12588 9824 12640
rect 12624 12588 12676 12640
rect 15568 12588 15620 12640
rect 15936 12588 15988 12640
rect 18144 12588 18196 12640
rect 22928 12588 22980 12640
rect 23756 12588 23808 12640
rect 24584 12588 24636 12640
rect 25412 12631 25464 12640
rect 25412 12597 25421 12631
rect 25421 12597 25455 12631
rect 25455 12597 25464 12631
rect 25412 12588 25464 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 2044 12427 2096 12436
rect 2044 12393 2053 12427
rect 2053 12393 2087 12427
rect 2087 12393 2096 12427
rect 2044 12384 2096 12393
rect 2320 12427 2372 12436
rect 2320 12393 2329 12427
rect 2329 12393 2363 12427
rect 2363 12393 2372 12427
rect 2320 12384 2372 12393
rect 2780 12384 2832 12436
rect 4620 12384 4672 12436
rect 4804 12427 4856 12436
rect 4804 12393 4813 12427
rect 4813 12393 4847 12427
rect 4847 12393 4856 12427
rect 4804 12384 4856 12393
rect 5632 12427 5684 12436
rect 5632 12393 5641 12427
rect 5641 12393 5675 12427
rect 5675 12393 5684 12427
rect 5632 12384 5684 12393
rect 7012 12384 7064 12436
rect 8300 12384 8352 12436
rect 4896 12316 4948 12368
rect 7380 12316 7432 12368
rect 9588 12384 9640 12436
rect 11612 12384 11664 12436
rect 12900 12427 12952 12436
rect 12900 12393 12909 12427
rect 12909 12393 12943 12427
rect 12943 12393 12952 12427
rect 12900 12384 12952 12393
rect 13544 12427 13596 12436
rect 13544 12393 13553 12427
rect 13553 12393 13587 12427
rect 13587 12393 13596 12427
rect 13544 12384 13596 12393
rect 20536 12384 20588 12436
rect 1584 12248 1636 12300
rect 2596 12248 2648 12300
rect 2964 12248 3016 12300
rect 5448 12248 5500 12300
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 6276 12248 6328 12300
rect 7196 12248 7248 12300
rect 7840 12248 7892 12300
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 11428 12248 11480 12300
rect 12164 12248 12216 12300
rect 15384 12248 15436 12300
rect 15568 12291 15620 12300
rect 15568 12257 15602 12291
rect 15602 12257 15620 12291
rect 15568 12248 15620 12257
rect 16856 12248 16908 12300
rect 18604 12291 18656 12300
rect 18604 12257 18638 12291
rect 18638 12257 18656 12291
rect 18604 12248 18656 12257
rect 20444 12248 20496 12300
rect 21640 12316 21692 12368
rect 24400 12384 24452 12436
rect 24952 12384 25004 12436
rect 25596 12384 25648 12436
rect 22560 12316 22612 12368
rect 23112 12248 23164 12300
rect 24584 12316 24636 12368
rect 6460 12180 6512 12232
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 10140 12180 10192 12232
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 18328 12223 18380 12232
rect 18328 12189 18337 12223
rect 18337 12189 18371 12223
rect 18371 12189 18380 12223
rect 18328 12180 18380 12189
rect 20720 12223 20772 12232
rect 20720 12189 20729 12223
rect 20729 12189 20763 12223
rect 20763 12189 20772 12223
rect 20720 12180 20772 12189
rect 22192 12180 22244 12232
rect 6920 12112 6972 12164
rect 8576 12112 8628 12164
rect 11428 12112 11480 12164
rect 22008 12112 22060 12164
rect 25044 12180 25096 12232
rect 24308 12155 24360 12164
rect 24308 12121 24317 12155
rect 24317 12121 24351 12155
rect 24351 12121 24360 12155
rect 24308 12112 24360 12121
rect 26148 12112 26200 12164
rect 8300 12087 8352 12096
rect 8300 12053 8309 12087
rect 8309 12053 8343 12087
rect 8343 12053 8352 12087
rect 8300 12044 8352 12053
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 11520 12044 11572 12096
rect 12624 12044 12676 12096
rect 14464 12044 14516 12096
rect 16212 12044 16264 12096
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 16948 12044 17000 12096
rect 17868 12044 17920 12096
rect 18144 12087 18196 12096
rect 18144 12053 18153 12087
rect 18153 12053 18187 12087
rect 18187 12053 18196 12087
rect 18144 12044 18196 12053
rect 19432 12044 19484 12096
rect 20168 12044 20220 12096
rect 20444 12044 20496 12096
rect 24216 12044 24268 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 5264 11840 5316 11892
rect 6092 11883 6144 11892
rect 6092 11849 6101 11883
rect 6101 11849 6135 11883
rect 6135 11849 6144 11883
rect 6092 11840 6144 11849
rect 7196 11883 7248 11892
rect 7196 11849 7205 11883
rect 7205 11849 7239 11883
rect 7239 11849 7248 11883
rect 7196 11840 7248 11849
rect 7564 11883 7616 11892
rect 7564 11849 7573 11883
rect 7573 11849 7607 11883
rect 7607 11849 7616 11883
rect 7564 11840 7616 11849
rect 5080 11772 5132 11824
rect 6276 11772 6328 11824
rect 7748 11704 7800 11756
rect 9128 11840 9180 11892
rect 10048 11840 10100 11892
rect 10784 11883 10836 11892
rect 10784 11849 10793 11883
rect 10793 11849 10827 11883
rect 10827 11849 10836 11883
rect 10784 11840 10836 11849
rect 11520 11840 11572 11892
rect 15476 11840 15528 11892
rect 21640 11840 21692 11892
rect 22836 11840 22888 11892
rect 23020 11883 23072 11892
rect 23020 11849 23029 11883
rect 23029 11849 23063 11883
rect 23063 11849 23072 11883
rect 23020 11840 23072 11849
rect 23664 11883 23716 11892
rect 23664 11849 23673 11883
rect 23673 11849 23707 11883
rect 23707 11849 23716 11883
rect 23664 11840 23716 11849
rect 24860 11840 24912 11892
rect 26148 11883 26200 11892
rect 26148 11849 26157 11883
rect 26157 11849 26191 11883
rect 26191 11849 26200 11883
rect 26148 11840 26200 11849
rect 9312 11772 9364 11824
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 6460 11636 6512 11688
rect 7104 11636 7156 11688
rect 9404 11704 9456 11756
rect 14464 11772 14516 11824
rect 15568 11772 15620 11824
rect 16028 11772 16080 11824
rect 8576 11636 8628 11688
rect 9220 11636 9272 11688
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 11428 11747 11480 11756
rect 11428 11713 11437 11747
rect 11437 11713 11471 11747
rect 11471 11713 11480 11747
rect 11428 11704 11480 11713
rect 16212 11747 16264 11756
rect 16212 11713 16221 11747
rect 16221 11713 16255 11747
rect 16255 11713 16264 11747
rect 16212 11704 16264 11713
rect 25044 11772 25096 11824
rect 16672 11704 16724 11756
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 18420 11704 18472 11756
rect 24216 11747 24268 11756
rect 24216 11713 24225 11747
rect 24225 11713 24259 11747
rect 24259 11713 24268 11747
rect 24216 11704 24268 11713
rect 11152 11679 11204 11688
rect 11152 11645 11161 11679
rect 11161 11645 11195 11679
rect 11195 11645 11204 11679
rect 11152 11636 11204 11645
rect 12624 11636 12676 11688
rect 8300 11568 8352 11620
rect 9680 11611 9732 11620
rect 9680 11577 9689 11611
rect 9689 11577 9723 11611
rect 9723 11577 9732 11611
rect 9680 11568 9732 11577
rect 12164 11611 12216 11620
rect 12164 11577 12173 11611
rect 12173 11577 12207 11611
rect 12207 11577 12216 11611
rect 12164 11568 12216 11577
rect 13176 11568 13228 11620
rect 19524 11636 19576 11688
rect 18328 11568 18380 11620
rect 20720 11636 20772 11688
rect 22284 11636 22336 11688
rect 23020 11636 23072 11688
rect 24032 11679 24084 11688
rect 24032 11645 24041 11679
rect 24041 11645 24075 11679
rect 24075 11645 24084 11679
rect 24032 11636 24084 11645
rect 25688 11636 25740 11688
rect 20168 11611 20220 11620
rect 20168 11577 20202 11611
rect 20202 11577 20220 11611
rect 20168 11568 20220 11577
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 17408 11500 17460 11552
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 18144 11500 18196 11552
rect 21456 11500 21508 11552
rect 22192 11500 22244 11552
rect 22468 11500 22520 11552
rect 23480 11543 23532 11552
rect 23480 11509 23489 11543
rect 23489 11509 23523 11543
rect 23523 11509 23532 11543
rect 23480 11500 23532 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1768 11296 1820 11348
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 6828 11296 6880 11348
rect 7380 11296 7432 11348
rect 8484 11296 8536 11348
rect 8944 11296 8996 11348
rect 9312 11339 9364 11348
rect 9312 11305 9321 11339
rect 9321 11305 9355 11339
rect 9355 11305 9364 11339
rect 9312 11296 9364 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 11244 11296 11296 11348
rect 14280 11296 14332 11348
rect 15660 11296 15712 11348
rect 15936 11296 15988 11348
rect 16580 11296 16632 11348
rect 18052 11296 18104 11348
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 18604 11296 18656 11348
rect 21272 11296 21324 11348
rect 23112 11296 23164 11348
rect 24032 11339 24084 11348
rect 24032 11305 24041 11339
rect 24041 11305 24075 11339
rect 24075 11305 24084 11339
rect 24032 11296 24084 11305
rect 24952 11296 25004 11348
rect 25412 11296 25464 11348
rect 25596 11339 25648 11348
rect 25596 11305 25605 11339
rect 25605 11305 25639 11339
rect 25639 11305 25648 11339
rect 25596 11296 25648 11305
rect 7104 11228 7156 11280
rect 10048 11228 10100 11280
rect 11152 11228 11204 11280
rect 12256 11228 12308 11280
rect 15568 11271 15620 11280
rect 15568 11237 15602 11271
rect 15602 11237 15620 11271
rect 15568 11228 15620 11237
rect 16028 11228 16080 11280
rect 23296 11228 23348 11280
rect 8392 11160 8444 11212
rect 11796 11160 11848 11212
rect 12440 11160 12492 11212
rect 15292 11203 15344 11212
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 11704 11135 11756 11144
rect 8576 11092 8628 11101
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 12900 11092 12952 11144
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 13176 11092 13228 11101
rect 13820 11092 13872 11144
rect 6000 11024 6052 11076
rect 10876 11067 10928 11076
rect 10876 11033 10885 11067
rect 10885 11033 10919 11067
rect 10919 11033 10928 11067
rect 10876 11024 10928 11033
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 15936 11160 15988 11212
rect 18052 11160 18104 11212
rect 19432 11160 19484 11212
rect 24952 11203 25004 11212
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 10784 10956 10836 11008
rect 14188 11024 14240 11076
rect 19340 11024 19392 11076
rect 20168 11024 20220 11076
rect 24952 11169 24961 11203
rect 24961 11169 24995 11203
rect 24995 11169 25004 11203
rect 24952 11160 25004 11169
rect 21732 11024 21784 11076
rect 12532 10999 12584 11008
rect 12532 10965 12541 10999
rect 12541 10965 12575 10999
rect 12575 10965 12584 10999
rect 12532 10956 12584 10965
rect 21916 10956 21968 11008
rect 24860 11092 24912 11144
rect 22468 10956 22520 11008
rect 23020 10956 23072 11008
rect 24124 10956 24176 11008
rect 25044 10956 25096 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 8208 10752 8260 10804
rect 8484 10795 8536 10804
rect 8484 10761 8493 10795
rect 8493 10761 8527 10795
rect 8527 10761 8536 10795
rect 8484 10752 8536 10761
rect 9220 10795 9272 10804
rect 9220 10761 9229 10795
rect 9229 10761 9263 10795
rect 9263 10761 9272 10795
rect 9220 10752 9272 10761
rect 9680 10752 9732 10804
rect 12164 10752 12216 10804
rect 8576 10684 8628 10736
rect 11152 10684 11204 10736
rect 9312 10616 9364 10668
rect 11244 10659 11296 10668
rect 11244 10625 11253 10659
rect 11253 10625 11287 10659
rect 11287 10625 11296 10659
rect 11244 10616 11296 10625
rect 11612 10616 11664 10668
rect 12624 10752 12676 10804
rect 13820 10795 13872 10804
rect 13820 10761 13829 10795
rect 13829 10761 13863 10795
rect 13863 10761 13872 10795
rect 13820 10752 13872 10761
rect 16396 10752 16448 10804
rect 17960 10752 18012 10804
rect 18052 10684 18104 10736
rect 15016 10616 15068 10668
rect 19248 10752 19300 10804
rect 20720 10752 20772 10804
rect 23020 10795 23072 10804
rect 19984 10727 20036 10736
rect 19984 10693 19993 10727
rect 19993 10693 20027 10727
rect 20027 10693 20036 10727
rect 19984 10684 20036 10693
rect 9496 10548 9548 10600
rect 12532 10548 12584 10600
rect 10140 10480 10192 10532
rect 13820 10480 13872 10532
rect 15292 10523 15344 10532
rect 9680 10455 9732 10464
rect 9680 10421 9689 10455
rect 9689 10421 9723 10455
rect 9723 10421 9732 10455
rect 9680 10412 9732 10421
rect 10692 10412 10744 10464
rect 10876 10412 10928 10464
rect 11796 10455 11848 10464
rect 11796 10421 11805 10455
rect 11805 10421 11839 10455
rect 11839 10421 11848 10455
rect 11796 10412 11848 10421
rect 15292 10489 15301 10523
rect 15301 10489 15335 10523
rect 15335 10489 15344 10523
rect 15292 10480 15344 10489
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 16028 10455 16080 10464
rect 15384 10412 15436 10421
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 16580 10412 16632 10464
rect 19340 10616 19392 10668
rect 23020 10761 23029 10795
rect 23029 10761 23063 10795
rect 23063 10761 23072 10795
rect 23020 10752 23072 10761
rect 23572 10752 23624 10804
rect 23848 10752 23900 10804
rect 24032 10752 24084 10804
rect 24952 10752 25004 10804
rect 25504 10752 25556 10804
rect 25320 10684 25372 10736
rect 20260 10548 20312 10600
rect 24124 10548 24176 10600
rect 25228 10591 25280 10600
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25228 10548 25280 10557
rect 21456 10480 21508 10532
rect 18604 10455 18656 10464
rect 18604 10421 18613 10455
rect 18613 10421 18647 10455
rect 18647 10421 18656 10455
rect 18604 10412 18656 10421
rect 18972 10412 19024 10464
rect 22192 10412 22244 10464
rect 23848 10412 23900 10464
rect 24216 10412 24268 10464
rect 24860 10412 24912 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 10692 10208 10744 10260
rect 10968 10208 11020 10260
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 14188 10251 14240 10260
rect 14188 10217 14197 10251
rect 14197 10217 14231 10251
rect 14231 10217 14240 10251
rect 14188 10208 14240 10217
rect 15016 10251 15068 10260
rect 15016 10217 15025 10251
rect 15025 10217 15059 10251
rect 15059 10217 15068 10251
rect 15016 10208 15068 10217
rect 15292 10208 15344 10260
rect 15568 10251 15620 10260
rect 15568 10217 15577 10251
rect 15577 10217 15611 10251
rect 15611 10217 15620 10251
rect 15568 10208 15620 10217
rect 23020 10208 23072 10260
rect 23296 10251 23348 10260
rect 23296 10217 23305 10251
rect 23305 10217 23339 10251
rect 23339 10217 23348 10251
rect 23296 10208 23348 10217
rect 24124 10208 24176 10260
rect 24584 10208 24636 10260
rect 25044 10208 25096 10260
rect 10784 10140 10836 10192
rect 16396 10140 16448 10192
rect 24860 10140 24912 10192
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 11520 10072 11572 10124
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 16028 10115 16080 10124
rect 16028 10081 16037 10115
rect 16037 10081 16071 10115
rect 16071 10081 16080 10115
rect 16028 10072 16080 10081
rect 18972 10072 19024 10124
rect 22192 10115 22244 10124
rect 22192 10081 22226 10115
rect 22226 10081 22244 10115
rect 22192 10072 22244 10081
rect 24124 10072 24176 10124
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 19248 10047 19300 10056
rect 19248 10013 19257 10047
rect 19257 10013 19291 10047
rect 19291 10013 19300 10047
rect 19248 10004 19300 10013
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 20720 10004 20772 10056
rect 21916 10047 21968 10056
rect 21916 10013 21925 10047
rect 21925 10013 21959 10047
rect 21959 10013 21968 10047
rect 21916 10004 21968 10013
rect 9588 9936 9640 9988
rect 18604 9936 18656 9988
rect 23112 9936 23164 9988
rect 12348 9868 12400 9920
rect 12532 9868 12584 9920
rect 13452 9868 13504 9920
rect 17684 9868 17736 9920
rect 18328 9911 18380 9920
rect 18328 9877 18337 9911
rect 18337 9877 18371 9911
rect 18371 9877 18380 9911
rect 18328 9868 18380 9877
rect 20260 9911 20312 9920
rect 20260 9877 20269 9911
rect 20269 9877 20303 9911
rect 20303 9877 20312 9911
rect 20260 9868 20312 9877
rect 23848 9911 23900 9920
rect 23848 9877 23857 9911
rect 23857 9877 23891 9911
rect 23891 9877 23900 9911
rect 23848 9868 23900 9877
rect 24952 9868 25004 9920
rect 25688 9868 25740 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 12164 9707 12216 9716
rect 12164 9673 12173 9707
rect 12173 9673 12207 9707
rect 12207 9673 12216 9707
rect 12164 9664 12216 9673
rect 12808 9664 12860 9716
rect 9680 9596 9732 9648
rect 11244 9596 11296 9648
rect 12532 9596 12584 9648
rect 9956 9528 10008 9580
rect 10140 9528 10192 9580
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 14740 9664 14792 9716
rect 15292 9664 15344 9716
rect 16396 9664 16448 9716
rect 16212 9639 16264 9648
rect 16212 9605 16221 9639
rect 16221 9605 16255 9639
rect 16255 9605 16264 9639
rect 16212 9596 16264 9605
rect 16764 9664 16816 9716
rect 16948 9664 17000 9716
rect 17776 9664 17828 9716
rect 21916 9664 21968 9716
rect 23020 9664 23072 9716
rect 23296 9664 23348 9716
rect 18236 9596 18288 9648
rect 19432 9596 19484 9648
rect 20444 9596 20496 9648
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 10048 9460 10100 9512
rect 9956 9392 10008 9444
rect 17040 9460 17092 9512
rect 18328 9503 18380 9512
rect 14280 9392 14332 9444
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 12348 9324 12400 9376
rect 12532 9367 12584 9376
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 16948 9324 17000 9376
rect 17132 9324 17184 9376
rect 18328 9469 18337 9503
rect 18337 9469 18371 9503
rect 18371 9469 18380 9503
rect 18328 9460 18380 9469
rect 22008 9503 22060 9512
rect 22008 9469 22017 9503
rect 22017 9469 22051 9503
rect 22051 9469 22060 9503
rect 22008 9460 22060 9469
rect 18512 9392 18564 9444
rect 20904 9392 20956 9444
rect 23664 9664 23716 9716
rect 24124 9707 24176 9716
rect 24124 9673 24133 9707
rect 24133 9673 24167 9707
rect 24167 9673 24176 9707
rect 24124 9664 24176 9673
rect 24676 9596 24728 9648
rect 24860 9596 24912 9648
rect 23664 9460 23716 9512
rect 23940 9460 23992 9512
rect 24952 9392 25004 9444
rect 19524 9324 19576 9376
rect 20536 9324 20588 9376
rect 21088 9324 21140 9376
rect 21640 9367 21692 9376
rect 21640 9333 21649 9367
rect 21649 9333 21683 9367
rect 21683 9333 21692 9367
rect 21640 9324 21692 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 10968 9120 11020 9172
rect 12072 9120 12124 9172
rect 13728 9120 13780 9172
rect 14648 9120 14700 9172
rect 16488 9120 16540 9172
rect 16856 9120 16908 9172
rect 19524 9163 19576 9172
rect 19524 9129 19533 9163
rect 19533 9129 19567 9163
rect 19567 9129 19576 9163
rect 19524 9120 19576 9129
rect 20536 9163 20588 9172
rect 20536 9129 20545 9163
rect 20545 9129 20579 9163
rect 20579 9129 20588 9163
rect 20536 9120 20588 9129
rect 20904 9163 20956 9172
rect 20904 9129 20913 9163
rect 20913 9129 20947 9163
rect 20947 9129 20956 9163
rect 20904 9120 20956 9129
rect 21640 9120 21692 9172
rect 22468 9163 22520 9172
rect 14556 9095 14608 9104
rect 14556 9061 14565 9095
rect 14565 9061 14599 9095
rect 14599 9061 14608 9095
rect 14556 9052 14608 9061
rect 22192 9052 22244 9104
rect 22468 9129 22477 9163
rect 22477 9129 22511 9163
rect 22511 9129 22520 9163
rect 22468 9120 22520 9129
rect 23112 9120 23164 9172
rect 24768 9163 24820 9172
rect 24768 9129 24777 9163
rect 24777 9129 24811 9163
rect 24811 9129 24820 9163
rect 24768 9120 24820 9129
rect 22928 9095 22980 9104
rect 22928 9061 22937 9095
rect 22937 9061 22971 9095
rect 22971 9061 22980 9095
rect 22928 9052 22980 9061
rect 9680 8984 9732 9036
rect 12532 8984 12584 9036
rect 13820 8984 13872 9036
rect 13912 8984 13964 9036
rect 15936 9027 15988 9036
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 17776 8984 17828 9036
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 23848 8984 23900 9036
rect 25044 8984 25096 9036
rect 12348 8848 12400 8900
rect 13544 8891 13596 8900
rect 13544 8857 13553 8891
rect 13553 8857 13587 8891
rect 13587 8857 13596 8891
rect 13544 8848 13596 8857
rect 14280 8916 14332 8968
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 17132 8959 17184 8968
rect 16120 8916 16172 8925
rect 14740 8848 14792 8900
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 19616 8959 19668 8968
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 19892 8916 19944 8968
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 23296 8916 23348 8968
rect 18512 8891 18564 8900
rect 18512 8857 18521 8891
rect 18521 8857 18555 8891
rect 18555 8857 18564 8891
rect 18512 8848 18564 8857
rect 13360 8823 13412 8832
rect 13360 8789 13369 8823
rect 13369 8789 13403 8823
rect 13403 8789 13412 8823
rect 13360 8780 13412 8789
rect 16580 8823 16632 8832
rect 16580 8789 16589 8823
rect 16589 8789 16623 8823
rect 16623 8789 16632 8823
rect 16580 8780 16632 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 12532 8576 12584 8628
rect 12900 8619 12952 8628
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 13912 8619 13964 8628
rect 13912 8585 13921 8619
rect 13921 8585 13955 8619
rect 13955 8585 13964 8619
rect 13912 8576 13964 8585
rect 15384 8576 15436 8628
rect 16120 8576 16172 8628
rect 17132 8576 17184 8628
rect 18972 8619 19024 8628
rect 18972 8585 18981 8619
rect 18981 8585 19015 8619
rect 19015 8585 19024 8619
rect 18972 8576 19024 8585
rect 19340 8576 19392 8628
rect 21272 8576 21324 8628
rect 22928 8619 22980 8628
rect 22928 8585 22937 8619
rect 22937 8585 22971 8619
rect 22971 8585 22980 8619
rect 22928 8576 22980 8585
rect 23112 8576 23164 8628
rect 24032 8576 24084 8628
rect 24860 8619 24912 8628
rect 24860 8585 24869 8619
rect 24869 8585 24903 8619
rect 24903 8585 24912 8619
rect 24860 8576 24912 8585
rect 25044 8576 25096 8628
rect 13360 8508 13412 8560
rect 14832 8508 14884 8560
rect 15936 8508 15988 8560
rect 19892 8508 19944 8560
rect 23296 8508 23348 8560
rect 25412 8508 25464 8560
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 14740 8440 14792 8492
rect 16304 8440 16356 8492
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 20628 8440 20680 8492
rect 20904 8440 20956 8492
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 13360 8372 13412 8424
rect 14556 8372 14608 8424
rect 16764 8415 16816 8424
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 19616 8372 19668 8424
rect 11980 8347 12032 8356
rect 11980 8313 11989 8347
rect 11989 8313 12023 8347
rect 12023 8313 12032 8347
rect 11980 8304 12032 8313
rect 11244 8279 11296 8288
rect 11244 8245 11253 8279
rect 11253 8245 11287 8279
rect 11287 8245 11296 8279
rect 11244 8236 11296 8245
rect 13728 8304 13780 8356
rect 14648 8304 14700 8356
rect 16580 8304 16632 8356
rect 17868 8304 17920 8356
rect 18788 8347 18840 8356
rect 18788 8313 18797 8347
rect 18797 8313 18831 8347
rect 18831 8313 18840 8347
rect 18788 8304 18840 8313
rect 21364 8372 21416 8424
rect 24032 8372 24084 8424
rect 24768 8372 24820 8424
rect 20904 8347 20956 8356
rect 20904 8313 20913 8347
rect 20913 8313 20947 8347
rect 20947 8313 20956 8347
rect 20904 8304 20956 8313
rect 16304 8279 16356 8288
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 16304 8236 16356 8245
rect 24032 8236 24084 8288
rect 25780 8236 25832 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 11520 8032 11572 8084
rect 13452 8032 13504 8084
rect 13728 8032 13780 8084
rect 14096 8032 14148 8084
rect 14740 8075 14792 8084
rect 14740 8041 14749 8075
rect 14749 8041 14783 8075
rect 14783 8041 14792 8075
rect 14740 8032 14792 8041
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 16764 8032 16816 8084
rect 20628 8075 20680 8084
rect 20628 8041 20637 8075
rect 20637 8041 20671 8075
rect 20671 8041 20680 8075
rect 20628 8032 20680 8041
rect 21456 8075 21508 8084
rect 21456 8041 21465 8075
rect 21465 8041 21499 8075
rect 21499 8041 21508 8075
rect 21456 8032 21508 8041
rect 22560 8032 22612 8084
rect 23940 8075 23992 8084
rect 23940 8041 23949 8075
rect 23949 8041 23983 8075
rect 23983 8041 23992 8075
rect 23940 8032 23992 8041
rect 25136 8032 25188 8084
rect 11244 7964 11296 8016
rect 12348 7964 12400 8016
rect 16488 7964 16540 8016
rect 19340 8007 19392 8016
rect 19340 7973 19349 8007
rect 19349 7973 19383 8007
rect 19383 7973 19392 8007
rect 19340 7964 19392 7973
rect 11888 7896 11940 7948
rect 12164 7828 12216 7880
rect 17684 7896 17736 7948
rect 20996 7896 21048 7948
rect 23204 7896 23256 7948
rect 23664 7896 23716 7948
rect 24768 7939 24820 7948
rect 24768 7905 24777 7939
rect 24777 7905 24811 7939
rect 24811 7905 24820 7939
rect 24768 7896 24820 7905
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 16488 7871 16540 7880
rect 16488 7837 16497 7871
rect 16497 7837 16531 7871
rect 16531 7837 16540 7871
rect 16488 7828 16540 7837
rect 17500 7828 17552 7880
rect 19064 7828 19116 7880
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 20628 7828 20680 7880
rect 12716 7760 12768 7812
rect 17776 7760 17828 7812
rect 21088 7803 21140 7812
rect 21088 7769 21097 7803
rect 21097 7769 21131 7803
rect 21131 7769 21140 7803
rect 21088 7760 21140 7769
rect 14280 7692 14332 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 11244 7488 11296 7540
rect 14832 7531 14884 7540
rect 14832 7497 14841 7531
rect 14841 7497 14875 7531
rect 14875 7497 14884 7531
rect 14832 7488 14884 7497
rect 15292 7531 15344 7540
rect 15292 7497 15301 7531
rect 15301 7497 15335 7531
rect 15335 7497 15344 7531
rect 15292 7488 15344 7497
rect 15752 7488 15804 7540
rect 16028 7488 16080 7540
rect 17868 7488 17920 7540
rect 19064 7531 19116 7540
rect 19064 7497 19073 7531
rect 19073 7497 19107 7531
rect 19107 7497 19116 7531
rect 19064 7488 19116 7497
rect 19984 7488 20036 7540
rect 20628 7531 20680 7540
rect 20628 7497 20637 7531
rect 20637 7497 20671 7531
rect 20671 7497 20680 7531
rect 20628 7488 20680 7497
rect 20996 7531 21048 7540
rect 20996 7497 21005 7531
rect 21005 7497 21039 7531
rect 21039 7497 21048 7531
rect 20996 7488 21048 7497
rect 23204 7488 23256 7540
rect 23664 7488 23716 7540
rect 24768 7488 24820 7540
rect 16488 7420 16540 7472
rect 24032 7420 24084 7472
rect 16304 7352 16356 7404
rect 17684 7352 17736 7404
rect 19616 7352 19668 7404
rect 20076 7395 20128 7404
rect 20076 7361 20085 7395
rect 20085 7361 20119 7395
rect 20119 7361 20128 7395
rect 20076 7352 20128 7361
rect 20352 7352 20404 7404
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 23756 7352 23808 7404
rect 12716 7327 12768 7336
rect 12716 7293 12725 7327
rect 12725 7293 12759 7327
rect 12759 7293 12768 7327
rect 12716 7284 12768 7293
rect 15292 7284 15344 7336
rect 16764 7327 16816 7336
rect 16764 7293 16773 7327
rect 16773 7293 16807 7327
rect 16807 7293 16816 7327
rect 16764 7284 16816 7293
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 23664 7284 23716 7293
rect 14740 7216 14792 7268
rect 18512 7259 18564 7268
rect 18512 7225 18521 7259
rect 18521 7225 18555 7259
rect 18555 7225 18564 7259
rect 18512 7216 18564 7225
rect 20168 7216 20220 7268
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 18236 7148 18288 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 15476 6944 15528 6996
rect 17500 6987 17552 6996
rect 17500 6953 17509 6987
rect 17509 6953 17543 6987
rect 17543 6953 17552 6987
rect 17500 6944 17552 6953
rect 20352 6944 20404 6996
rect 15936 6919 15988 6928
rect 15936 6885 15945 6919
rect 15945 6885 15979 6919
rect 15979 6885 15988 6919
rect 15936 6876 15988 6885
rect 17592 6919 17644 6928
rect 17592 6885 17601 6919
rect 17601 6885 17635 6919
rect 17635 6885 17644 6919
rect 17592 6876 17644 6885
rect 15384 6808 15436 6860
rect 16396 6808 16448 6860
rect 19248 6808 19300 6860
rect 20076 6808 20128 6860
rect 23664 6851 23716 6860
rect 23664 6817 23673 6851
rect 23673 6817 23707 6851
rect 23707 6817 23716 6851
rect 23664 6808 23716 6817
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 16856 6672 16908 6724
rect 25872 6672 25924 6724
rect 16672 6604 16724 6656
rect 18236 6647 18288 6656
rect 18236 6613 18245 6647
rect 18245 6613 18279 6647
rect 18279 6613 18288 6647
rect 18236 6604 18288 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 15384 6400 15436 6452
rect 15936 6443 15988 6452
rect 15936 6409 15945 6443
rect 15945 6409 15979 6443
rect 15979 6409 15988 6443
rect 15936 6400 15988 6409
rect 16396 6443 16448 6452
rect 16396 6409 16405 6443
rect 16405 6409 16439 6443
rect 16439 6409 16448 6443
rect 16396 6400 16448 6409
rect 17500 6443 17552 6452
rect 17500 6409 17509 6443
rect 17509 6409 17543 6443
rect 17543 6409 17552 6443
rect 17500 6400 17552 6409
rect 23664 6400 23716 6452
rect 17132 6103 17184 6112
rect 17132 6069 17141 6103
rect 17141 6069 17175 6103
rect 17175 6069 17184 6103
rect 17132 6060 17184 6069
rect 17592 6060 17644 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 13728 2456 13780 2508
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 12900 2431 12952 2440
rect 11980 2388 12032 2397
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 2042 27520 2098 28000
rect 2594 27520 2650 28000
rect 3146 27520 3202 28000
rect 3790 27520 3846 28000
rect 4342 27520 4398 28000
rect 4434 27704 4490 27713
rect 4434 27639 4490 27648
rect 308 15473 336 27520
rect 860 19990 888 27520
rect 1214 26616 1270 26625
rect 1214 26551 1270 26560
rect 1228 22234 1256 26551
rect 1306 24848 1362 24857
rect 1306 24783 1362 24792
rect 1320 23594 1348 24783
rect 1308 23588 1360 23594
rect 1308 23530 1360 23536
rect 1412 23338 1440 27520
rect 2056 25922 2084 27520
rect 1780 25894 2084 25922
rect 2228 25900 2280 25906
rect 1674 25392 1730 25401
rect 1674 25327 1730 25336
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1492 24880 1544 24886
rect 1492 24822 1544 24828
rect 1504 23474 1532 24822
rect 1596 24410 1624 24890
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1504 23446 1624 23474
rect 1412 23310 1532 23338
rect 1400 23248 1452 23254
rect 1400 23190 1452 23196
rect 1412 22522 1440 23190
rect 1320 22494 1440 22522
rect 1216 22228 1268 22234
rect 1216 22170 1268 22176
rect 848 19984 900 19990
rect 1320 19972 1348 22494
rect 1400 22432 1452 22438
rect 1400 22374 1452 22380
rect 1412 21026 1440 22374
rect 1504 21146 1532 23310
rect 1596 23118 1624 23446
rect 1584 23112 1636 23118
rect 1584 23054 1636 23060
rect 1688 23050 1716 25327
rect 1780 23254 1808 25894
rect 2228 25842 2280 25848
rect 1952 25764 2004 25770
rect 1952 25706 2004 25712
rect 1964 25498 1992 25706
rect 1952 25492 2004 25498
rect 1952 25434 2004 25440
rect 1964 25242 1992 25434
rect 1964 25214 2084 25242
rect 1952 25152 2004 25158
rect 1952 25094 2004 25100
rect 1964 24750 1992 25094
rect 2056 24818 2084 25214
rect 2240 24818 2268 25842
rect 2504 25356 2556 25362
rect 2504 25298 2556 25304
rect 2516 25265 2544 25298
rect 2502 25256 2558 25265
rect 2502 25191 2558 25200
rect 2504 25152 2556 25158
rect 2504 25094 2556 25100
rect 2516 24886 2544 25094
rect 2504 24880 2556 24886
rect 2318 24848 2374 24857
rect 2044 24812 2096 24818
rect 2044 24754 2096 24760
rect 2228 24812 2280 24818
rect 2504 24822 2556 24828
rect 2318 24783 2374 24792
rect 2228 24754 2280 24760
rect 1952 24744 2004 24750
rect 1952 24686 2004 24692
rect 1860 24608 1912 24614
rect 1860 24550 1912 24556
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 1872 23730 1900 24550
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1768 23248 1820 23254
rect 1768 23190 1820 23196
rect 1964 23066 1992 24550
rect 2240 24426 2268 24754
rect 2056 24410 2268 24426
rect 2332 24410 2360 24783
rect 2044 24404 2268 24410
rect 2096 24398 2268 24404
rect 2320 24404 2372 24410
rect 2044 24346 2096 24352
rect 2320 24346 2372 24352
rect 2136 24336 2188 24342
rect 2136 24278 2188 24284
rect 2044 24268 2096 24274
rect 2044 24210 2096 24216
rect 2056 23769 2084 24210
rect 2042 23760 2098 23769
rect 2042 23695 2098 23704
rect 2148 23662 2176 24278
rect 2608 24274 2636 27520
rect 3054 26072 3110 26081
rect 3054 26007 3110 26016
rect 2688 25968 2740 25974
rect 2688 25910 2740 25916
rect 2320 24268 2372 24274
rect 2320 24210 2372 24216
rect 2596 24268 2648 24274
rect 2596 24210 2648 24216
rect 2136 23656 2188 23662
rect 2136 23598 2188 23604
rect 2332 23474 2360 24210
rect 2412 24064 2464 24070
rect 2412 24006 2464 24012
rect 1676 23044 1728 23050
rect 1676 22986 1728 22992
rect 1872 23038 1992 23066
rect 2148 23446 2360 23474
rect 1688 22166 1716 22986
rect 1768 22432 1820 22438
rect 1766 22400 1768 22409
rect 1820 22400 1822 22409
rect 1766 22335 1822 22344
rect 1676 22160 1728 22166
rect 1728 22120 1808 22148
rect 1676 22102 1728 22108
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1596 21690 1624 21830
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 21185 1624 21286
rect 1582 21176 1638 21185
rect 1492 21140 1544 21146
rect 1638 21134 1716 21162
rect 1780 21146 1808 22120
rect 1582 21111 1638 21120
rect 1492 21082 1544 21088
rect 1412 20998 1624 21026
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 20097 1440 20878
rect 1596 20346 1624 20998
rect 1504 20318 1624 20346
rect 1398 20088 1454 20097
rect 1398 20023 1454 20032
rect 1320 19944 1440 19972
rect 848 19926 900 19932
rect 1412 18578 1440 19944
rect 1504 18834 1532 20318
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1492 18828 1544 18834
rect 1492 18770 1544 18776
rect 1412 18550 1532 18578
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 294 15464 350 15473
rect 294 15399 350 15408
rect 1412 11694 1440 18022
rect 1504 17785 1532 18550
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1504 17270 1532 17614
rect 1596 17513 1624 20198
rect 1688 19310 1716 21134
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1872 20602 1900 23038
rect 1952 22976 2004 22982
rect 1952 22918 2004 22924
rect 1964 22681 1992 22918
rect 1950 22672 2006 22681
rect 1950 22607 2006 22616
rect 1964 22574 1992 22607
rect 1952 22568 2004 22574
rect 1952 22510 2004 22516
rect 1952 21888 2004 21894
rect 1952 21830 2004 21836
rect 1964 21350 1992 21830
rect 2044 21684 2096 21690
rect 2044 21626 2096 21632
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 1860 20596 1912 20602
rect 1860 20538 1912 20544
rect 1872 20398 1900 20538
rect 1860 20392 1912 20398
rect 1780 20340 1860 20346
rect 1780 20334 1912 20340
rect 1780 20318 1900 20334
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1688 18154 1716 19110
rect 1676 18148 1728 18154
rect 1676 18090 1728 18096
rect 1582 17504 1638 17513
rect 1582 17439 1638 17448
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1492 17264 1544 17270
rect 1492 17206 1544 17212
rect 1596 16794 1624 17274
rect 1780 16998 1808 20318
rect 1860 20052 1912 20058
rect 1860 19994 1912 20000
rect 1872 19825 1900 19994
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 19378 1900 19654
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1872 17882 1900 19314
rect 1964 18970 1992 21286
rect 2056 19174 2084 21626
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2056 19009 2084 19110
rect 2042 19000 2098 19009
rect 1952 18964 2004 18970
rect 2042 18935 2098 18944
rect 1952 18906 2004 18912
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1964 18290 1992 18566
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1964 17921 1992 18022
rect 1950 17912 2006 17921
rect 1860 17876 1912 17882
rect 1950 17847 2006 17856
rect 1860 17818 1912 17824
rect 1964 17354 1992 17847
rect 2148 17626 2176 23446
rect 2424 23089 2452 24006
rect 2700 23866 2728 25910
rect 3068 25514 3096 26007
rect 3160 25702 3188 27520
rect 3804 25838 3832 27520
rect 3792 25832 3844 25838
rect 3792 25774 3844 25780
rect 3148 25696 3200 25702
rect 3148 25638 3200 25644
rect 3068 25486 3188 25514
rect 3056 25424 3108 25430
rect 3056 25366 3108 25372
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2792 24886 2820 25298
rect 2964 25288 3016 25294
rect 2964 25230 3016 25236
rect 2976 24993 3004 25230
rect 2962 24984 3018 24993
rect 2962 24919 3018 24928
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 2792 24614 2820 24822
rect 2872 24676 2924 24682
rect 2872 24618 2924 24624
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2884 24410 2912 24618
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 2884 23798 2912 24346
rect 2872 23792 2924 23798
rect 2872 23734 2924 23740
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2410 23080 2466 23089
rect 2410 23015 2466 23024
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2332 22642 2360 22918
rect 2320 22636 2372 22642
rect 2320 22578 2372 22584
rect 2516 22522 2544 23666
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2870 23488 2926 23497
rect 2700 23338 2728 23462
rect 2870 23423 2926 23432
rect 2700 23322 2820 23338
rect 2700 23316 2832 23322
rect 2700 23310 2780 23316
rect 2780 23258 2832 23264
rect 2596 22976 2648 22982
rect 2596 22918 2648 22924
rect 2332 22494 2544 22522
rect 2608 22506 2636 22918
rect 2596 22500 2648 22506
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 2240 21554 2268 21966
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2240 20602 2268 21490
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2240 17814 2268 20538
rect 2332 20466 2360 22494
rect 2596 22442 2648 22448
rect 2504 22432 2556 22438
rect 2504 22374 2556 22380
rect 2410 21312 2466 21321
rect 2410 21247 2466 21256
rect 2424 21146 2452 21247
rect 2412 21140 2464 21146
rect 2412 21082 2464 21088
rect 2412 20800 2464 20806
rect 2412 20742 2464 20748
rect 2320 20460 2372 20466
rect 2320 20402 2372 20408
rect 2318 20224 2374 20233
rect 2318 20159 2374 20168
rect 2332 20058 2360 20159
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2320 19848 2372 19854
rect 2320 19790 2372 19796
rect 2332 19446 2360 19790
rect 2320 19440 2372 19446
rect 2320 19382 2372 19388
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2228 17808 2280 17814
rect 2228 17750 2280 17756
rect 1872 17326 1992 17354
rect 2056 17598 2176 17626
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1688 16250 1716 16730
rect 1768 16516 1820 16522
rect 1768 16458 1820 16464
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1596 15745 1624 15846
rect 1582 15736 1638 15745
rect 1582 15671 1638 15680
rect 1780 15586 1808 16458
rect 1872 15706 1900 17326
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 1964 16794 1992 17206
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1780 15558 1900 15586
rect 1582 14648 1638 14657
rect 1582 14583 1638 14592
rect 1596 14074 1624 14583
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1490 13968 1546 13977
rect 1688 13938 1716 14214
rect 1490 13903 1546 13912
rect 1676 13932 1728 13938
rect 1504 12986 1532 13903
rect 1676 13874 1728 13880
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1596 13433 1624 13466
rect 1582 13424 1638 13433
rect 1582 13359 1638 13368
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1582 12880 1638 12889
rect 1582 12815 1638 12824
rect 1596 12442 1624 12815
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1596 11898 1624 12242
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1780 11354 1808 14282
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1872 9081 1900 15558
rect 1964 13530 1992 16594
rect 2056 15706 2084 17598
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2056 14822 2084 15506
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2056 12442 2084 14758
rect 2148 14618 2176 17478
rect 2240 16794 2268 17750
rect 2332 17134 2360 17818
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2240 16454 2268 16730
rect 2332 16658 2360 17070
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2226 16280 2282 16289
rect 2226 16215 2282 16224
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2240 13258 2268 16215
rect 2332 15858 2360 16594
rect 2424 16561 2452 20742
rect 2516 16726 2544 22374
rect 2596 22228 2648 22234
rect 2596 22170 2648 22176
rect 2608 21690 2636 22170
rect 2884 21894 2912 23423
rect 2962 23352 3018 23361
rect 2962 23287 3018 23296
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2596 21412 2648 21418
rect 2596 21354 2648 21360
rect 2608 21078 2636 21354
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 2608 19922 2636 20198
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2608 17542 2636 19858
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2504 16720 2556 16726
rect 2504 16662 2556 16668
rect 2410 16552 2466 16561
rect 2608 16522 2636 16934
rect 2410 16487 2466 16496
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2332 15830 2452 15858
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2332 15094 2360 15506
rect 2424 15502 2452 15830
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2516 15144 2544 16390
rect 2700 15314 2728 20402
rect 2792 20058 2820 20878
rect 2884 20448 2912 21626
rect 2976 21457 3004 23287
rect 3068 23225 3096 25366
rect 3054 23216 3110 23225
rect 3054 23151 3110 23160
rect 3056 23112 3108 23118
rect 3056 23054 3108 23060
rect 3068 22234 3096 23054
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 3056 21956 3108 21962
rect 3056 21898 3108 21904
rect 2962 21448 3018 21457
rect 2962 21383 3018 21392
rect 2884 20420 3004 20448
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19514 2820 19858
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2884 19394 2912 19994
rect 2976 19553 3004 20420
rect 2962 19544 3018 19553
rect 2962 19479 3018 19488
rect 2792 19366 2912 19394
rect 2792 19310 2820 19366
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2976 18902 3004 18933
rect 2964 18896 3016 18902
rect 2962 18864 2964 18873
rect 3016 18864 3018 18873
rect 2962 18799 3018 18808
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2778 18184 2834 18193
rect 2884 18154 2912 18702
rect 2976 18426 3004 18799
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2778 18119 2834 18128
rect 2872 18148 2924 18154
rect 2792 17338 2820 18119
rect 2872 18090 2924 18096
rect 2976 17746 3004 18158
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 3068 17116 3096 21898
rect 3160 19922 3188 25486
rect 3608 25492 3660 25498
rect 3608 25434 3660 25440
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3436 24750 3464 25094
rect 3240 24744 3292 24750
rect 3240 24686 3292 24692
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 3252 24410 3280 24686
rect 3330 24576 3386 24585
rect 3330 24511 3386 24520
rect 3240 24404 3292 24410
rect 3240 24346 3292 24352
rect 3252 23730 3280 24346
rect 3344 24274 3372 24511
rect 3332 24268 3384 24274
rect 3332 24210 3384 24216
rect 3344 23866 3372 24210
rect 3332 23860 3384 23866
rect 3332 23802 3384 23808
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 3252 23322 3280 23666
rect 3240 23316 3292 23322
rect 3240 23258 3292 23264
rect 3238 23216 3294 23225
rect 3238 23151 3240 23160
rect 3292 23151 3294 23160
rect 3240 23122 3292 23128
rect 3436 23118 3464 24686
rect 3620 24614 3648 25434
rect 3700 25152 3752 25158
rect 3700 25094 3752 25100
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3620 24177 3648 24550
rect 3606 24168 3662 24177
rect 3516 24132 3568 24138
rect 3606 24103 3662 24112
rect 3516 24074 3568 24080
rect 3528 23798 3556 24074
rect 3516 23792 3568 23798
rect 3516 23734 3568 23740
rect 3528 23254 3556 23734
rect 3608 23656 3660 23662
rect 3608 23598 3660 23604
rect 3516 23248 3568 23254
rect 3516 23190 3568 23196
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3528 22778 3556 23190
rect 3620 22794 3648 23598
rect 3712 23050 3740 25094
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3896 24410 3924 24550
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3790 24304 3846 24313
rect 3790 24239 3846 24248
rect 3700 23044 3752 23050
rect 3700 22986 3752 22992
rect 3516 22772 3568 22778
rect 3620 22766 3740 22794
rect 3516 22714 3568 22720
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 3344 21146 3372 21422
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3330 21040 3386 21049
rect 3330 20975 3332 20984
rect 3384 20975 3386 20984
rect 3332 20946 3384 20952
rect 3238 20768 3294 20777
rect 3238 20703 3294 20712
rect 3252 20330 3280 20703
rect 3344 20602 3372 20946
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 3330 20496 3386 20505
rect 3330 20431 3332 20440
rect 3384 20431 3386 20440
rect 3332 20402 3384 20408
rect 3240 20324 3292 20330
rect 3240 20266 3292 20272
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3146 19816 3202 19825
rect 3146 19751 3202 19760
rect 2976 17088 3096 17116
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2424 15116 2544 15144
rect 2608 15286 2728 15314
rect 2320 15088 2372 15094
rect 2320 15030 2372 15036
rect 2332 13530 2360 15030
rect 2424 14958 2452 15116
rect 2502 15056 2558 15065
rect 2502 14991 2504 15000
rect 2556 14991 2558 15000
rect 2504 14962 2556 14968
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 14074 2452 14350
rect 2516 14278 2544 14758
rect 2608 14618 2636 15286
rect 2686 15192 2742 15201
rect 2686 15127 2742 15136
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2608 14006 2636 14554
rect 2700 14074 2728 15127
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2596 14000 2648 14006
rect 2596 13942 2648 13948
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2700 13682 2728 13874
rect 2700 13654 2820 13682
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2228 13252 2280 13258
rect 2228 13194 2280 13200
rect 2136 12640 2188 12646
rect 2134 12608 2136 12617
rect 2188 12608 2190 12617
rect 2134 12543 2190 12552
rect 2332 12442 2360 13330
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2700 12345 2728 12582
rect 2792 12442 2820 13654
rect 2884 13530 2912 16730
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2686 12336 2742 12345
rect 2596 12300 2648 12306
rect 2976 12306 3004 17088
rect 3160 16794 3188 19751
rect 3252 18698 3280 20266
rect 3344 20233 3372 20402
rect 3330 20224 3386 20233
rect 3330 20159 3386 20168
rect 3332 19984 3384 19990
rect 3332 19926 3384 19932
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3344 18578 3372 19926
rect 3436 18902 3464 21830
rect 3620 21418 3648 21830
rect 3608 21412 3660 21418
rect 3608 21354 3660 21360
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3528 20602 3556 20878
rect 3620 20806 3648 21354
rect 3608 20800 3660 20806
rect 3608 20742 3660 20748
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3528 19530 3556 20538
rect 3528 19502 3648 19530
rect 3514 19408 3570 19417
rect 3620 19378 3648 19502
rect 3514 19343 3570 19352
rect 3608 19372 3660 19378
rect 3424 18896 3476 18902
rect 3424 18838 3476 18844
rect 3252 18550 3372 18578
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 3068 15706 3096 16526
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3252 15586 3280 18550
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3344 15745 3372 15914
rect 3330 15736 3386 15745
rect 3330 15671 3332 15680
rect 3384 15671 3386 15680
rect 3332 15642 3384 15648
rect 3068 15558 3280 15586
rect 3068 13569 3096 15558
rect 3238 14784 3294 14793
rect 3238 14719 3294 14728
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3054 13560 3110 13569
rect 3054 13495 3110 13504
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3068 12986 3096 13330
rect 3160 13190 3188 14418
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3068 12753 3096 12922
rect 3160 12889 3188 13126
rect 3146 12880 3202 12889
rect 3146 12815 3202 12824
rect 3054 12744 3110 12753
rect 3054 12679 3110 12688
rect 2686 12271 2742 12280
rect 2964 12300 3016 12306
rect 2596 12242 2648 12248
rect 2964 12242 3016 12248
rect 2608 11898 2636 12242
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 3252 11801 3280 14719
rect 3436 14260 3464 18566
rect 3528 15314 3556 19343
rect 3608 19314 3660 19320
rect 3606 19272 3662 19281
rect 3606 19207 3662 19216
rect 3620 19174 3648 19207
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 3620 15502 3648 18702
rect 3712 18408 3740 22766
rect 3804 19802 3832 24239
rect 3896 23594 3924 24346
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 3884 23588 3936 23594
rect 3884 23530 3936 23536
rect 3896 22642 3924 23530
rect 4080 23497 4108 24006
rect 4066 23488 4122 23497
rect 4066 23423 4122 23432
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 3882 21448 3938 21457
rect 3882 21383 3938 21392
rect 3896 20913 3924 21383
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3882 20904 3938 20913
rect 3882 20839 3938 20848
rect 3804 19774 3924 19802
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3804 19378 3832 19654
rect 3896 19446 3924 19774
rect 3884 19440 3936 19446
rect 3884 19382 3936 19388
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3988 19310 4016 21286
rect 4068 21072 4120 21078
rect 4068 21014 4120 21020
rect 4080 20913 4108 21014
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4066 20904 4122 20913
rect 4066 20839 4122 20848
rect 4080 20058 4108 20839
rect 4172 20466 4200 20946
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4172 19922 4200 20402
rect 4356 19961 4384 27520
rect 4448 24410 4476 27639
rect 4894 27520 4950 28000
rect 5538 27520 5594 28000
rect 6090 27520 6146 28000
rect 6642 27520 6698 28000
rect 7286 27520 7342 28000
rect 7838 27520 7894 28000
rect 8390 27520 8446 28000
rect 9034 27520 9090 28000
rect 9586 27520 9642 28000
rect 10138 27520 10194 28000
rect 10782 27520 10838 28000
rect 11334 27520 11390 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 16026 27520 16082 28000
rect 16578 27520 16634 28000
rect 17130 27520 17186 28000
rect 17774 27520 17830 28000
rect 18326 27520 18382 28000
rect 18878 27520 18934 28000
rect 19522 27520 19578 28000
rect 20074 27520 20130 28000
rect 20626 27520 20682 28000
rect 21270 27520 21326 28000
rect 21822 27520 21878 28000
rect 22374 27520 22430 28000
rect 23018 27520 23074 28000
rect 23570 27520 23626 28000
rect 23938 27704 23994 27713
rect 23938 27639 23994 27648
rect 4802 27160 4858 27169
rect 4802 27095 4858 27104
rect 4816 25498 4844 27095
rect 4804 25492 4856 25498
rect 4804 25434 4856 25440
rect 4816 24886 4844 25434
rect 4804 24880 4856 24886
rect 4804 24822 4856 24828
rect 4436 24404 4488 24410
rect 4436 24346 4488 24352
rect 4448 23322 4476 24346
rect 4528 24268 4580 24274
rect 4528 24210 4580 24216
rect 4436 23316 4488 23322
rect 4436 23258 4488 23264
rect 4448 21350 4476 23258
rect 4540 22982 4568 24210
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4632 23866 4660 24142
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 4632 22710 4660 23802
rect 4620 22704 4672 22710
rect 4620 22646 4672 22652
rect 4816 22642 4844 24822
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4620 22160 4672 22166
rect 4620 22102 4672 22108
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4540 21593 4568 21966
rect 4526 21584 4582 21593
rect 4526 21519 4582 21528
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4436 21140 4488 21146
rect 4436 21082 4488 21088
rect 4448 20262 4476 21082
rect 4540 20602 4568 21519
rect 4632 21321 4660 22102
rect 4618 21312 4674 21321
rect 4618 21247 4674 21256
rect 4724 21146 4752 22374
rect 4712 21140 4764 21146
rect 4712 21082 4764 21088
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4436 20256 4488 20262
rect 4804 20256 4856 20262
rect 4436 20198 4488 20204
rect 4802 20224 4804 20233
rect 4856 20224 4858 20233
rect 4802 20159 4858 20168
rect 4434 20088 4490 20097
rect 4434 20023 4436 20032
rect 4488 20023 4490 20032
rect 4436 19994 4488 20000
rect 4342 19952 4398 19961
rect 4160 19916 4212 19922
rect 4342 19887 4398 19896
rect 4160 19858 4212 19864
rect 4344 19712 4396 19718
rect 4342 19680 4344 19689
rect 4396 19680 4398 19689
rect 4342 19615 4398 19624
rect 4342 19544 4398 19553
rect 4068 19508 4120 19514
rect 4448 19514 4476 19994
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4342 19479 4398 19488
rect 4436 19508 4488 19514
rect 4068 19450 4120 19456
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3792 18420 3844 18426
rect 3712 18380 3792 18408
rect 3792 18362 3844 18368
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3804 17882 3832 18158
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 3804 17338 3832 17818
rect 3896 17728 3924 19246
rect 3988 18970 4016 19246
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 4080 17864 4108 19450
rect 4356 19360 4384 19479
rect 4436 19450 4488 19456
rect 4356 19332 4476 19360
rect 4448 18766 4476 19332
rect 4540 19281 4568 19790
rect 4816 19514 4844 20159
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4526 19272 4582 19281
rect 4526 19207 4582 19216
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4080 17836 4200 17864
rect 3976 17740 4028 17746
rect 3896 17700 3976 17728
rect 3976 17682 4028 17688
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3988 17270 4016 17682
rect 4080 17338 4108 17682
rect 4172 17338 4200 17836
rect 4264 17785 4292 18090
rect 4250 17776 4306 17785
rect 4250 17711 4306 17720
rect 4448 17542 4476 18702
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4540 18358 4568 18566
rect 4528 18352 4580 18358
rect 4528 18294 4580 18300
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 4080 16810 4108 17274
rect 4344 17264 4396 17270
rect 4344 17206 4396 17212
rect 3988 16782 4108 16810
rect 4250 16824 4306 16833
rect 3988 16522 4016 16782
rect 4250 16759 4252 16768
rect 4304 16759 4306 16768
rect 4252 16730 4304 16736
rect 4356 16658 4384 17206
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 3712 15609 3740 16458
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3698 15600 3754 15609
rect 3698 15535 3700 15544
rect 3752 15535 3754 15544
rect 3700 15506 3752 15512
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3882 15464 3938 15473
rect 3882 15399 3938 15408
rect 3528 15286 3648 15314
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3344 14232 3464 14260
rect 3344 13569 3372 14232
rect 3528 13802 3556 14758
rect 3620 14414 3648 15286
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3896 13938 3924 15399
rect 3988 15026 4016 15846
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3988 14618 4016 14962
rect 4080 14906 4108 16594
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 4080 14878 4200 14906
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4080 14657 4108 14758
rect 4066 14648 4122 14657
rect 3976 14612 4028 14618
rect 4172 14618 4200 14878
rect 4066 14583 4122 14592
rect 4160 14612 4212 14618
rect 3976 14554 4028 14560
rect 4160 14554 4212 14560
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 3884 13796 3936 13802
rect 3884 13738 3936 13744
rect 3330 13560 3386 13569
rect 3330 13495 3386 13504
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3238 11792 3294 11801
rect 3238 11727 3294 11736
rect 2962 9344 3018 9353
rect 2962 9279 3018 9288
rect 1858 9072 1914 9081
rect 1858 9007 1914 9016
rect 2976 7177 3004 9279
rect 2962 7168 3018 7177
rect 2962 7103 3018 7112
rect 3146 3632 3202 3641
rect 3146 3567 3202 3576
rect 3160 921 3188 3567
rect 3436 2938 3464 12582
rect 3528 9217 3556 13738
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3698 13696 3754 13705
rect 3620 12986 3648 13670
rect 3698 13631 3754 13640
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3620 12782 3648 12922
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3712 9489 3740 13631
rect 3896 13530 3924 13738
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13530 4016 13670
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4264 13326 4292 16458
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4356 15706 4384 15982
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4356 14550 4384 15438
rect 4344 14544 4396 14550
rect 4344 14486 4396 14492
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4264 12986 4292 13262
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4066 11792 4122 11801
rect 4066 11727 4122 11736
rect 3882 10432 3938 10441
rect 3882 10367 3938 10376
rect 3698 9480 3754 9489
rect 3698 9415 3754 9424
rect 3514 9208 3570 9217
rect 3514 9143 3570 9152
rect 3896 4865 3924 10367
rect 4080 10033 4108 11727
rect 4448 11393 4476 17478
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4434 11384 4490 11393
rect 4434 11319 4490 11328
rect 4540 10305 4568 15574
rect 4632 14890 4660 19110
rect 4804 18896 4856 18902
rect 4804 18838 4856 18844
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4724 18222 4752 18770
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4620 14884 4672 14890
rect 4620 14826 4672 14832
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4632 12442 4660 14418
rect 4724 12986 4752 16050
rect 4816 15706 4844 18838
rect 4908 17785 4936 27520
rect 5552 25378 5580 27520
rect 5448 25356 5500 25362
rect 5552 25350 6040 25378
rect 5448 25298 5500 25304
rect 5172 25220 5224 25226
rect 5172 25162 5224 25168
rect 5184 24206 5212 25162
rect 5460 24886 5488 25298
rect 5906 25256 5962 25265
rect 5906 25191 5908 25200
rect 5960 25191 5962 25200
rect 5908 25162 5960 25168
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5448 24880 5500 24886
rect 5448 24822 5500 24828
rect 5552 24750 5580 25094
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5540 24744 5592 24750
rect 6012 24721 6040 25350
rect 6104 24993 6132 27520
rect 6276 25900 6328 25906
rect 6276 25842 6328 25848
rect 6090 24984 6146 24993
rect 6090 24919 6146 24928
rect 5540 24686 5592 24692
rect 5998 24712 6054 24721
rect 6104 24682 6132 24919
rect 5998 24647 6054 24656
rect 6092 24676 6144 24682
rect 6092 24618 6144 24624
rect 6000 24608 6052 24614
rect 6000 24550 6052 24556
rect 5172 24200 5224 24206
rect 5172 24142 5224 24148
rect 5354 24168 5410 24177
rect 5354 24103 5410 24112
rect 5368 23866 5396 24103
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5000 22778 5028 23122
rect 4988 22772 5040 22778
rect 4988 22714 5040 22720
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5000 18970 5028 22578
rect 5368 21962 5396 22578
rect 5460 22098 5488 23122
rect 5552 22778 5580 24006
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5644 23254 5672 23462
rect 6012 23361 6040 24550
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6104 23526 6132 24278
rect 6092 23520 6144 23526
rect 6092 23462 6144 23468
rect 5998 23352 6054 23361
rect 5998 23287 6054 23296
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5998 23080 6054 23089
rect 5998 23015 6054 23024
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 6012 22574 6040 23015
rect 6104 22817 6132 23462
rect 6090 22808 6146 22817
rect 6090 22743 6146 22752
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 5540 22432 5592 22438
rect 5538 22400 5540 22409
rect 5592 22400 5594 22409
rect 5538 22335 5594 22344
rect 5552 22234 5580 22335
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5448 22092 5500 22098
rect 5448 22034 5500 22040
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 5460 21690 5488 22034
rect 6104 22030 6132 22743
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 6104 21486 6132 21966
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5368 20777 5396 20878
rect 5448 20800 5500 20806
rect 5354 20768 5410 20777
rect 5448 20742 5500 20748
rect 5354 20703 5410 20712
rect 5460 20534 5488 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5460 19922 5488 20198
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 6000 19916 6052 19922
rect 6104 19904 6132 21422
rect 6288 20618 6316 25842
rect 6460 25832 6512 25838
rect 6460 25774 6512 25780
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6380 23798 6408 24210
rect 6368 23792 6420 23798
rect 6368 23734 6420 23740
rect 6368 22976 6420 22982
rect 6368 22918 6420 22924
rect 6380 22098 6408 22918
rect 6368 22092 6420 22098
rect 6368 22034 6420 22040
rect 6380 21690 6408 22034
rect 6472 21865 6500 25774
rect 6552 25356 6604 25362
rect 6552 25298 6604 25304
rect 6564 24614 6592 25298
rect 6656 25242 6684 27520
rect 7300 25498 7328 27520
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 6656 25214 6776 25242
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6552 24608 6604 24614
rect 6552 24550 6604 24556
rect 6564 23594 6592 24550
rect 6656 23769 6684 25094
rect 6642 23760 6698 23769
rect 6642 23695 6698 23704
rect 6552 23588 6604 23594
rect 6552 23530 6604 23536
rect 6564 23118 6592 23530
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6458 21856 6514 21865
rect 6458 21791 6514 21800
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6366 21176 6422 21185
rect 6366 21111 6368 21120
rect 6420 21111 6422 21120
rect 6368 21082 6420 21088
rect 6288 20590 6408 20618
rect 6276 20528 6328 20534
rect 6276 20470 6328 20476
rect 6288 19990 6316 20470
rect 6380 20097 6408 20590
rect 6366 20088 6422 20097
rect 6366 20023 6422 20032
rect 6276 19984 6328 19990
rect 6276 19926 6328 19932
rect 6052 19876 6132 19904
rect 6000 19858 6052 19864
rect 5460 19378 5488 19858
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6104 19514 6132 19876
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 6184 19304 6236 19310
rect 6184 19246 6236 19252
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 5000 17882 5028 18906
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 5092 18426 5120 18770
rect 5184 18698 5212 19110
rect 6104 18766 6132 19110
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5446 18456 5502 18465
rect 5080 18420 5132 18426
rect 5622 18448 5918 18468
rect 5446 18391 5502 18400
rect 5080 18362 5132 18368
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 4894 17776 4950 17785
rect 4894 17711 4950 17720
rect 5000 17134 5028 17818
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4816 15162 4844 15642
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4908 13530 4936 16934
rect 5000 16794 5028 17070
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5092 16182 5120 18362
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 16794 5212 18022
rect 5460 17338 5488 18391
rect 6104 18358 6132 18702
rect 6196 18630 6224 19246
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 5816 18080 5868 18086
rect 5814 18048 5816 18057
rect 5868 18048 5870 18057
rect 5814 17983 5870 17992
rect 5538 17912 5594 17921
rect 5538 17847 5540 17856
rect 5592 17847 5594 17856
rect 5540 17818 5592 17824
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5538 17232 5594 17241
rect 5356 17196 5408 17202
rect 5538 17167 5540 17176
rect 5356 17138 5408 17144
rect 5592 17167 5594 17176
rect 5540 17138 5592 17144
rect 5368 17105 5396 17138
rect 5354 17096 5410 17105
rect 5354 17031 5410 17040
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5552 16726 5580 17138
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5184 16250 5212 16526
rect 5460 16250 5488 16594
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5080 16176 5132 16182
rect 5080 16118 5132 16124
rect 5446 16144 5502 16153
rect 5092 15978 5120 16118
rect 5552 16114 5580 16662
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5908 16176 5960 16182
rect 5908 16118 5960 16124
rect 5446 16079 5502 16088
rect 5540 16108 5592 16114
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 4986 15872 5042 15881
rect 4986 15807 5042 15816
rect 5000 15570 5028 15807
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 5000 15026 5028 15506
rect 5460 15502 5488 16079
rect 5540 16050 5592 16056
rect 5552 15706 5580 16050
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5920 15570 5948 16118
rect 6012 16046 6040 16934
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 5908 15564 5960 15570
rect 5960 15524 6040 15552
rect 5908 15506 5960 15512
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5354 15328 5410 15337
rect 5354 15263 5410 15272
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 5000 13734 5028 14826
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5092 14482 5120 14758
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4816 12986 4844 13330
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4724 12714 4752 12922
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4816 12442 4844 12922
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4908 12374 4936 13466
rect 5000 12646 5028 13670
rect 5092 13190 5120 14282
rect 5184 14006 5212 14894
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 5092 11830 5120 13126
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 5184 11354 5212 13942
rect 5276 11898 5304 14826
rect 5368 13977 5396 15263
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 15162 6040 15524
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5540 14408 5592 14414
rect 5538 14376 5540 14385
rect 5592 14376 5594 14385
rect 5828 14346 5856 14962
rect 6012 14414 6040 15098
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5538 14311 5594 14320
rect 5816 14340 5868 14346
rect 5552 14056 5580 14311
rect 5816 14282 5868 14288
rect 6104 14278 6132 18294
rect 6196 17785 6224 18566
rect 6182 17776 6238 17785
rect 6182 17711 6238 17720
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6196 15473 6224 17478
rect 6276 17264 6328 17270
rect 6276 17206 6328 17212
rect 6288 15638 6316 17206
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6182 15464 6238 15473
rect 6182 15399 6238 15408
rect 6288 15162 6316 15574
rect 6276 15156 6328 15162
rect 6196 15116 6276 15144
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5552 14028 5672 14056
rect 5354 13968 5410 13977
rect 5354 13903 5410 13912
rect 5644 13394 5672 14028
rect 6196 13938 6224 15116
rect 6276 15098 6328 15104
rect 6380 14822 6408 20023
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6274 14648 6330 14657
rect 6274 14583 6276 14592
rect 6328 14583 6330 14592
rect 6276 14554 6328 14560
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6288 14346 6316 14418
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6196 13462 6224 13874
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5630 12880 5686 12889
rect 5630 12815 5686 12824
rect 5724 12844 5776 12850
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5448 12300 5500 12306
rect 5552 12288 5580 12718
rect 5644 12442 5672 12815
rect 5724 12786 5776 12792
rect 5736 12714 5764 12786
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5500 12260 5580 12288
rect 6000 12300 6052 12306
rect 5448 12242 5500 12248
rect 6000 12242 6052 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 6012 11082 6040 12242
rect 6104 11898 6132 13262
rect 6196 12986 6224 13398
rect 6288 13326 6316 14282
rect 6380 14074 6408 14350
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6472 13530 6500 21286
rect 6564 18193 6592 22374
rect 6656 18442 6684 23695
rect 6748 22953 6776 25214
rect 7012 25152 7064 25158
rect 7012 25094 7064 25100
rect 6826 24848 6882 24857
rect 6826 24783 6882 24792
rect 6840 23769 6868 24783
rect 7024 24410 7052 25094
rect 7300 24857 7328 25434
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7286 24848 7342 24857
rect 7286 24783 7342 24792
rect 7472 24812 7524 24818
rect 7300 24750 7328 24783
rect 7472 24754 7524 24760
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 6826 23760 6882 23769
rect 6826 23695 6882 23704
rect 6932 23304 6960 24006
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 6840 23276 6960 23304
rect 6734 22944 6790 22953
rect 6734 22879 6790 22888
rect 6840 22710 6868 23276
rect 6918 23216 6974 23225
rect 6918 23151 6920 23160
rect 6972 23151 6974 23160
rect 6920 23122 6972 23128
rect 6828 22704 6880 22710
rect 6828 22646 6880 22652
rect 7024 22001 7052 23462
rect 7116 22982 7144 24006
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7010 21992 7066 22001
rect 7010 21927 7066 21936
rect 7116 21536 7144 22374
rect 7208 21554 7236 24550
rect 7300 24313 7328 24550
rect 7286 24304 7342 24313
rect 7286 24239 7342 24248
rect 7484 24070 7512 24754
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7470 22808 7526 22817
rect 7470 22743 7472 22752
rect 7524 22743 7526 22752
rect 7472 22714 7524 22720
rect 7668 21978 7696 25094
rect 7852 24834 7880 27520
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 7392 21950 7696 21978
rect 7760 24806 7880 24834
rect 7024 21508 7144 21536
rect 7196 21548 7248 21554
rect 6918 21448 6974 21457
rect 6918 21383 6974 21392
rect 6932 21185 6960 21383
rect 6918 21176 6974 21185
rect 6918 21111 6974 21120
rect 7024 21128 7052 21508
rect 7196 21490 7248 21496
rect 7208 21457 7236 21490
rect 7194 21448 7250 21457
rect 7194 21383 7250 21392
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7024 21100 7144 21128
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 7024 20913 7052 20946
rect 7010 20904 7066 20913
rect 6920 20868 6972 20874
rect 7010 20839 7066 20848
rect 6920 20810 6972 20816
rect 6734 20768 6790 20777
rect 6734 20703 6790 20712
rect 6748 19174 6776 20703
rect 6826 20632 6882 20641
rect 6826 20567 6828 20576
rect 6880 20567 6882 20576
rect 6828 20538 6880 20544
rect 6932 20330 6960 20810
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 7024 20466 7052 20742
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 6920 20324 6972 20330
rect 6920 20266 6972 20272
rect 6932 19786 6960 20266
rect 7024 20058 7052 20402
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6920 19168 6972 19174
rect 7116 19145 7144 21100
rect 7208 20913 7236 21286
rect 7194 20904 7250 20913
rect 7194 20839 7250 20848
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7208 19990 7236 20198
rect 7196 19984 7248 19990
rect 7196 19926 7248 19932
rect 6920 19110 6972 19116
rect 7102 19136 7158 19145
rect 6932 18902 6960 19110
rect 7102 19071 7158 19080
rect 7208 18970 7236 19926
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 6920 18896 6972 18902
rect 7300 18873 7328 19110
rect 6920 18838 6972 18844
rect 7286 18864 7342 18873
rect 6656 18414 6776 18442
rect 6550 18184 6606 18193
rect 6550 18119 6606 18128
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6564 13410 6592 14758
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6472 13382 6592 13410
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6380 12986 6408 13330
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6288 11830 6316 12242
rect 6472 12238 6500 13382
rect 6656 12782 6684 18022
rect 6748 14929 6776 18414
rect 6932 17814 6960 18838
rect 7286 18799 7342 18808
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7116 17882 7144 18702
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6840 16794 6868 17682
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6932 15450 6960 17546
rect 7208 16697 7236 18090
rect 7300 18086 7328 18634
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7194 16688 7250 16697
rect 7194 16623 7250 16632
rect 7300 16572 7328 18022
rect 7392 17513 7420 21950
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7668 21554 7696 21830
rect 7656 21548 7708 21554
rect 7656 21490 7708 21496
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7484 20330 7512 20946
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7576 20534 7604 20878
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 7472 20324 7524 20330
rect 7472 20266 7524 20272
rect 7378 17504 7434 17513
rect 7378 17439 7434 17448
rect 7378 16960 7434 16969
rect 7378 16895 7434 16904
rect 7116 16544 7328 16572
rect 7116 16402 7144 16544
rect 7116 16374 7236 16402
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 7024 15473 7052 15914
rect 7208 15910 7236 16374
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 6840 15422 6960 15450
rect 7010 15464 7066 15473
rect 6840 14958 6868 15422
rect 7010 15399 7066 15408
rect 7024 15162 7052 15399
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6828 14952 6880 14958
rect 6734 14920 6790 14929
rect 6828 14894 6880 14900
rect 6734 14855 6790 14864
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7024 13138 7052 14554
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 6932 13110 7052 13138
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6472 11694 6500 12174
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6840 11354 6868 12922
rect 6932 12170 6960 13110
rect 7010 12744 7066 12753
rect 7010 12679 7066 12688
rect 7024 12442 7052 12679
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 7116 11694 7144 14214
rect 7208 13920 7236 15846
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 14482 7328 15302
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7392 14074 7420 16895
rect 7484 15473 7512 20266
rect 7576 19378 7604 20470
rect 7668 20262 7696 21082
rect 7760 21010 7788 24806
rect 7932 24676 7984 24682
rect 7932 24618 7984 24624
rect 7944 24177 7972 24618
rect 7930 24168 7986 24177
rect 7930 24103 7932 24112
rect 7984 24103 7986 24112
rect 7932 24074 7984 24080
rect 7932 23520 7984 23526
rect 7838 23488 7894 23497
rect 7932 23462 7984 23468
rect 7838 23423 7894 23432
rect 7852 23254 7880 23423
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7838 22808 7894 22817
rect 7944 22794 7972 23462
rect 8036 23050 8064 25162
rect 8114 24712 8170 24721
rect 8312 24698 8340 25230
rect 8170 24670 8340 24698
rect 8114 24647 8170 24656
rect 8128 24614 8156 24647
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 23633 8156 24550
rect 8208 24268 8260 24274
rect 8404 24256 8432 27520
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8484 25356 8536 25362
rect 8484 25298 8536 25304
rect 8496 24410 8524 25298
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8588 24342 8616 24686
rect 8576 24336 8628 24342
rect 8576 24278 8628 24284
rect 8404 24228 8524 24256
rect 8208 24210 8260 24216
rect 8220 23662 8248 24210
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 8208 23656 8260 23662
rect 8114 23624 8170 23633
rect 8208 23598 8260 23604
rect 8114 23559 8170 23568
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8128 23322 8156 23462
rect 8116 23316 8168 23322
rect 8116 23258 8168 23264
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8024 23044 8076 23050
rect 8024 22986 8076 22992
rect 7894 22766 7972 22794
rect 7838 22743 7894 22752
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7576 18902 7604 19314
rect 7852 19258 7880 22743
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 7668 19230 7880 19258
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7576 17105 7604 17682
rect 7562 17096 7618 17105
rect 7562 17031 7618 17040
rect 7576 16794 7604 17031
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7470 15464 7526 15473
rect 7470 15399 7526 15408
rect 7470 15328 7526 15337
rect 7576 15314 7604 16594
rect 7526 15286 7604 15314
rect 7470 15263 7526 15272
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7208 13892 7512 13920
rect 7286 12744 7342 12753
rect 7286 12679 7288 12688
rect 7340 12679 7342 12688
rect 7288 12650 7340 12656
rect 7380 12368 7432 12374
rect 7378 12336 7380 12345
rect 7432 12336 7434 12345
rect 7196 12300 7248 12306
rect 7378 12271 7434 12280
rect 7196 12242 7248 12248
rect 7208 11898 7236 12242
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 7116 11286 7144 11630
rect 7392 11354 7420 12271
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 4526 10296 4582 10305
rect 4526 10231 4582 10240
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6550 8256 6606 8265
rect 6550 8191 6606 8200
rect 6564 7721 6592 8191
rect 6550 7712 6606 7721
rect 5622 7644 5918 7664
rect 6550 7647 6606 7656
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 7484 7585 7512 13892
rect 7576 11898 7604 15286
rect 7668 12782 7696 19230
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7852 19009 7880 19110
rect 7838 19000 7894 19009
rect 7838 18935 7894 18944
rect 7840 18760 7892 18766
rect 7838 18728 7840 18737
rect 7892 18728 7894 18737
rect 7760 18686 7838 18714
rect 7760 18426 7788 18686
rect 7838 18663 7894 18672
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 7840 18352 7892 18358
rect 7838 18320 7840 18329
rect 7892 18320 7894 18329
rect 7838 18255 7894 18264
rect 7748 18148 7800 18154
rect 7748 18090 7800 18096
rect 7760 17542 7788 18090
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7760 17134 7788 17478
rect 7852 17338 7880 17750
rect 7944 17678 7972 21490
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 8036 19689 8064 20198
rect 8022 19680 8078 19689
rect 8022 19615 8078 19624
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7944 17270 7972 17614
rect 8022 17368 8078 17377
rect 8022 17303 8078 17312
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 7748 17128 7800 17134
rect 8036 17116 8064 17303
rect 7748 17070 7800 17076
rect 7944 17088 8064 17116
rect 7760 16250 7788 17070
rect 7840 16992 7892 16998
rect 7838 16960 7840 16969
rect 7892 16960 7894 16969
rect 7838 16895 7894 16904
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 15722 7788 15846
rect 7838 15736 7894 15745
rect 7760 15694 7838 15722
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7760 12238 7788 15694
rect 7838 15671 7894 15680
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 7852 14385 7880 14826
rect 7838 14376 7894 14385
rect 7838 14311 7840 14320
rect 7892 14311 7894 14320
rect 7840 14282 7892 14288
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7852 13705 7880 13806
rect 7838 13696 7894 13705
rect 7838 13631 7894 13640
rect 7944 13546 7972 17088
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8036 16697 8064 16730
rect 8022 16688 8078 16697
rect 8022 16623 8078 16632
rect 8022 15600 8078 15609
rect 8022 15535 8078 15544
rect 7852 13518 7972 13546
rect 7852 12306 7880 13518
rect 8036 13258 8064 15535
rect 8128 14113 8156 23054
rect 8220 18306 8248 23598
rect 8312 22409 8340 24006
rect 8392 22500 8444 22506
rect 8392 22442 8444 22448
rect 8298 22400 8354 22409
rect 8298 22335 8354 22344
rect 8404 21894 8432 22442
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8298 21584 8354 21593
rect 8298 21519 8300 21528
rect 8352 21519 8354 21528
rect 8300 21490 8352 21496
rect 8404 21434 8432 21830
rect 8312 21406 8432 21434
rect 8312 21010 8340 21406
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8312 19417 8340 20946
rect 8392 20800 8444 20806
rect 8390 20768 8392 20777
rect 8444 20768 8446 20777
rect 8390 20703 8446 20712
rect 8496 20074 8524 24228
rect 8680 23610 8708 25774
rect 8760 25288 8812 25294
rect 8760 25230 8812 25236
rect 8772 24682 8800 25230
rect 8944 25152 8996 25158
rect 8944 25094 8996 25100
rect 8760 24676 8812 24682
rect 8760 24618 8812 24624
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8588 23582 8708 23610
rect 8588 22114 8616 23582
rect 8668 23520 8720 23526
rect 8666 23488 8668 23497
rect 8720 23488 8722 23497
rect 8666 23423 8722 23432
rect 8668 23316 8720 23322
rect 8668 23258 8720 23264
rect 8680 22234 8708 23258
rect 8864 23254 8892 23666
rect 8852 23248 8904 23254
rect 8852 23190 8904 23196
rect 8956 23118 8984 25094
rect 8760 23112 8812 23118
rect 8758 23080 8760 23089
rect 8944 23112 8996 23118
rect 8812 23080 8814 23089
rect 8944 23054 8996 23060
rect 8758 23015 8814 23024
rect 8772 22778 8800 23015
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8588 22086 8708 22114
rect 8576 21344 8628 21350
rect 8574 21312 8576 21321
rect 8628 21312 8630 21321
rect 8574 21247 8630 21256
rect 8404 20046 8524 20074
rect 8298 19408 8354 19417
rect 8298 19343 8354 19352
rect 8404 18426 8432 20046
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8496 19156 8524 19858
rect 8576 19168 8628 19174
rect 8496 19128 8576 19156
rect 8576 19110 8628 19116
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8220 18278 8340 18306
rect 8208 18216 8260 18222
rect 8206 18184 8208 18193
rect 8260 18184 8262 18193
rect 8206 18119 8262 18128
rect 8312 18068 8340 18278
rect 8220 18040 8340 18068
rect 8220 16794 8248 18040
rect 8404 17649 8432 18362
rect 8496 18290 8524 18566
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8390 17640 8446 17649
rect 8390 17575 8446 17584
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8390 17096 8446 17105
rect 8496 17066 8524 17478
rect 8390 17031 8446 17040
rect 8484 17060 8536 17066
rect 8404 16794 8432 17031
rect 8484 17002 8536 17008
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8404 16674 8432 16730
rect 8220 16646 8432 16674
rect 8220 15706 8248 16646
rect 8496 16153 8524 17002
rect 8298 16144 8354 16153
rect 8298 16079 8354 16088
rect 8482 16144 8538 16153
rect 8482 16079 8538 16088
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8114 14104 8170 14113
rect 8114 14039 8170 14048
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8128 13530 8156 13874
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 8128 12986 8156 13194
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 7932 12708 7984 12714
rect 7984 12668 8064 12696
rect 7932 12650 7984 12656
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7760 11762 7788 12174
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 8036 8945 8064 12668
rect 8220 12424 8248 13942
rect 8312 13462 8340 16079
rect 8588 16017 8616 19110
rect 8574 16008 8630 16017
rect 8574 15943 8630 15952
rect 8680 15706 8708 22086
rect 9048 21876 9076 27520
rect 9600 26042 9628 27520
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 9588 26036 9640 26042
rect 9588 25978 9640 25984
rect 9600 25362 9628 25978
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9864 24676 9916 24682
rect 9864 24618 9916 24624
rect 9588 24336 9640 24342
rect 9588 24278 9640 24284
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9324 23866 9352 24142
rect 9496 24064 9548 24070
rect 9496 24006 9548 24012
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9128 23792 9180 23798
rect 9128 23734 9180 23740
rect 9140 22778 9168 23734
rect 9324 23662 9352 23802
rect 9402 23760 9458 23769
rect 9402 23695 9458 23704
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9416 23508 9444 23695
rect 9324 23480 9444 23508
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 9048 21848 9260 21876
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8772 18222 8800 20198
rect 8864 20097 8892 20266
rect 8850 20088 8906 20097
rect 8850 20023 8852 20032
rect 8904 20023 8906 20032
rect 8852 19994 8904 20000
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8864 18766 8892 19110
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8772 15586 8800 18022
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8864 16425 8892 16526
rect 8850 16416 8906 16425
rect 8850 16351 8906 16360
rect 8864 15638 8892 16351
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8680 15558 8800 15586
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8496 13870 8524 14010
rect 8484 13864 8536 13870
rect 8404 13824 8484 13852
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8404 12889 8432 13824
rect 8484 13806 8536 13812
rect 8482 13560 8538 13569
rect 8482 13495 8484 13504
rect 8536 13495 8538 13504
rect 8484 13466 8536 13472
rect 8496 12986 8524 13466
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8390 12880 8446 12889
rect 8390 12815 8446 12824
rect 8300 12436 8352 12442
rect 8220 12396 8300 12424
rect 8300 12378 8352 12384
rect 8588 12170 8616 15506
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11626 8340 12038
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8390 11384 8446 11393
rect 8390 11319 8446 11328
rect 8484 11348 8536 11354
rect 8404 11218 8432 11319
rect 8484 11290 8536 11296
rect 8392 11212 8444 11218
rect 8220 11172 8392 11200
rect 8220 10810 8248 11172
rect 8392 11154 8444 11160
rect 8496 10810 8524 11290
rect 8588 11150 8616 11630
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8588 10742 8616 11086
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8680 9489 8708 15558
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8772 13938 8800 14418
rect 8864 14414 8892 14894
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8864 14074 8892 14350
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8772 12986 8800 13330
rect 8850 13152 8906 13161
rect 8850 13087 8906 13096
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8864 12730 8892 13087
rect 8772 12702 8892 12730
rect 8772 10713 8800 12702
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8864 11121 8892 12582
rect 8956 11354 8984 20878
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 9048 20505 9076 20742
rect 9034 20496 9090 20505
rect 9034 20431 9090 20440
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9048 18630 9076 19314
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 18465 9076 18566
rect 9034 18456 9090 18465
rect 9034 18391 9090 18400
rect 9034 17776 9090 17785
rect 9034 17711 9036 17720
rect 9088 17711 9090 17720
rect 9036 17682 9088 17688
rect 9140 17626 9168 20266
rect 9232 19802 9260 21848
rect 9324 19922 9352 23480
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9416 22234 9444 23190
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9508 21434 9536 24006
rect 9600 23866 9628 24278
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9588 22024 9640 22030
rect 9692 22012 9720 22646
rect 9640 21984 9720 22012
rect 9588 21966 9640 21972
rect 9508 21406 9720 21434
rect 9692 21350 9720 21406
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9600 20602 9628 20946
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 9600 19854 9628 20198
rect 9588 19848 9640 19854
rect 9232 19774 9352 19802
rect 9588 19790 9640 19796
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 9048 17598 9168 17626
rect 9048 16658 9076 17598
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 9048 15910 9076 16594
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 9048 12782 9076 15846
rect 9232 14822 9260 19654
rect 9324 18601 9352 19774
rect 9692 19514 9720 21286
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9586 19408 9642 19417
rect 9586 19343 9642 19352
rect 9600 19310 9628 19343
rect 9784 19310 9812 23462
rect 9876 22574 9904 24618
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9968 24410 9996 24550
rect 10060 24449 10088 26182
rect 10152 24585 10180 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10692 25288 10744 25294
rect 10414 25256 10470 25265
rect 10692 25230 10744 25236
rect 10414 25191 10416 25200
rect 10468 25191 10470 25200
rect 10416 25162 10468 25168
rect 10704 24886 10732 25230
rect 10692 24880 10744 24886
rect 10692 24822 10744 24828
rect 10690 24712 10746 24721
rect 10690 24647 10746 24656
rect 10138 24576 10194 24585
rect 10138 24511 10194 24520
rect 10046 24440 10102 24449
rect 9956 24404 10008 24410
rect 10046 24375 10102 24384
rect 9956 24346 10008 24352
rect 9968 23594 9996 24346
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 9968 23254 9996 23530
rect 10060 23304 10088 24375
rect 10152 23905 10180 24511
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10704 24410 10732 24647
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10138 23896 10194 23905
rect 10138 23831 10194 23840
rect 10796 23526 10824 27520
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 10980 25498 11008 25842
rect 11348 25514 11376 27520
rect 11612 26172 11664 26178
rect 11612 26114 11664 26120
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 11256 25486 11376 25514
rect 11150 24848 11206 24857
rect 11150 24783 11206 24792
rect 11164 24410 11192 24783
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 10968 24336 11020 24342
rect 10966 24304 10968 24313
rect 11020 24304 11022 24313
rect 10966 24239 11022 24248
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10980 23322 11008 24239
rect 11060 23520 11112 23526
rect 11058 23488 11060 23497
rect 11112 23488 11114 23497
rect 11058 23423 11114 23432
rect 11164 23322 11192 24346
rect 11256 24342 11284 25486
rect 11520 25288 11572 25294
rect 11520 25230 11572 25236
rect 11532 24698 11560 25230
rect 11624 24886 11652 26114
rect 11704 25424 11756 25430
rect 11704 25366 11756 25372
rect 11612 24880 11664 24886
rect 11612 24822 11664 24828
rect 11440 24670 11560 24698
rect 11440 24614 11468 24670
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11244 24336 11296 24342
rect 11244 24278 11296 24284
rect 10968 23316 11020 23322
rect 10060 23276 10272 23304
rect 9956 23248 10008 23254
rect 9956 23190 10008 23196
rect 10138 23216 10194 23225
rect 10048 23180 10100 23186
rect 10138 23151 10194 23160
rect 10048 23122 10100 23128
rect 9954 22944 10010 22953
rect 9954 22879 10010 22888
rect 9864 22568 9916 22574
rect 9864 22510 9916 22516
rect 9862 22128 9918 22137
rect 9862 22063 9918 22072
rect 9876 21962 9904 22063
rect 9864 21956 9916 21962
rect 9864 21898 9916 21904
rect 9876 21486 9904 21898
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9310 18592 9366 18601
rect 9310 18527 9366 18536
rect 9324 17814 9352 18527
rect 9402 17912 9458 17921
rect 9402 17847 9458 17856
rect 9312 17808 9364 17814
rect 9312 17750 9364 17756
rect 9324 16726 9352 17750
rect 9416 17678 9444 17847
rect 9508 17785 9536 19110
rect 9600 18850 9628 19246
rect 9600 18822 9812 18850
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9692 18222 9720 18634
rect 9680 18216 9732 18222
rect 9600 18176 9680 18204
rect 9600 17882 9628 18176
rect 9680 18158 9732 18164
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9494 17776 9550 17785
rect 9692 17762 9720 18022
rect 9494 17711 9550 17720
rect 9600 17734 9720 17762
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9404 17264 9456 17270
rect 9402 17232 9404 17241
rect 9456 17232 9458 17241
rect 9402 17167 9458 17176
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9324 16046 9352 16186
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9324 15570 9352 15982
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 13938 9168 14214
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9126 13424 9182 13433
rect 9126 13359 9182 13368
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9036 12640 9088 12646
rect 9034 12608 9036 12617
rect 9088 12608 9090 12617
rect 9034 12543 9090 12552
rect 9140 11898 9168 13359
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9232 11694 9260 14758
rect 9310 13832 9366 13841
rect 9310 13767 9366 13776
rect 9324 11830 9352 13767
rect 9416 13326 9444 17167
rect 9508 16674 9536 17711
rect 9600 17542 9628 17734
rect 9678 17640 9734 17649
rect 9678 17575 9680 17584
rect 9732 17575 9734 17584
rect 9680 17546 9732 17552
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9692 16969 9720 17274
rect 9678 16960 9734 16969
rect 9678 16895 9734 16904
rect 9508 16646 9628 16674
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9508 15706 9536 16526
rect 9600 16522 9628 16646
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9692 16153 9720 16895
rect 9678 16144 9734 16153
rect 9678 16079 9734 16088
rect 9784 15706 9812 18822
rect 9876 18714 9904 21286
rect 9968 19174 9996 22879
rect 10060 22710 10088 23122
rect 10152 22953 10180 23151
rect 10138 22944 10194 22953
rect 10138 22879 10194 22888
rect 10048 22704 10100 22710
rect 10048 22646 10100 22652
rect 10244 22556 10272 23276
rect 10968 23258 11020 23264
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 10966 22944 11022 22953
rect 10966 22879 11022 22888
rect 10980 22642 11008 22879
rect 11334 22672 11390 22681
rect 10968 22636 11020 22642
rect 11334 22607 11390 22616
rect 10968 22578 11020 22584
rect 10060 22528 10272 22556
rect 10784 22568 10836 22574
rect 10060 22234 10088 22528
rect 10784 22510 10836 22516
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10048 22228 10100 22234
rect 10048 22170 10100 22176
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 10060 21146 10088 21558
rect 10152 21350 10180 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10690 22264 10746 22273
rect 10796 22234 10824 22510
rect 11152 22500 11204 22506
rect 11152 22442 11204 22448
rect 10690 22199 10746 22208
rect 10784 22228 10836 22234
rect 10704 22166 10732 22199
rect 10784 22170 10836 22176
rect 10692 22160 10744 22166
rect 10692 22102 10744 22108
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 10336 21690 10364 22034
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 10520 21622 10548 21966
rect 10704 21690 10732 22102
rect 10966 21720 11022 21729
rect 10692 21684 10744 21690
rect 10744 21644 10824 21672
rect 10692 21626 10744 21632
rect 10508 21616 10560 21622
rect 10508 21558 10560 21564
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10048 21140 10100 21146
rect 10100 21100 10180 21128
rect 10048 21082 10100 21088
rect 10048 20256 10100 20262
rect 10046 20224 10048 20233
rect 10100 20224 10102 20233
rect 10046 20159 10102 20168
rect 10048 19712 10100 19718
rect 10046 19680 10048 19689
rect 10100 19680 10102 19689
rect 10046 19615 10102 19624
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 9876 18686 9996 18714
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9508 14618 9536 15370
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9600 12850 9628 13398
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9680 12776 9732 12782
rect 9402 12744 9458 12753
rect 9600 12724 9680 12730
rect 9600 12718 9732 12724
rect 9402 12679 9458 12688
rect 9496 12708 9548 12714
rect 9312 11824 9364 11830
rect 9312 11766 9364 11772
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9324 11354 9352 11766
rect 9416 11762 9444 12679
rect 9496 12650 9548 12656
rect 9600 12702 9720 12718
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9402 11656 9458 11665
rect 9402 11591 9458 11600
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9218 11248 9274 11257
rect 9416 11234 9444 11591
rect 9218 11183 9274 11192
rect 9324 11206 9444 11234
rect 8850 11112 8906 11121
rect 8850 11047 8906 11056
rect 9232 10810 9260 11183
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 8758 10704 8814 10713
rect 9324 10674 9352 11206
rect 8758 10639 8814 10648
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 10266 9352 10610
rect 9508 10606 9536 12650
rect 9600 12442 9628 12702
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 10810 9720 11562
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9692 10010 9720 10406
rect 9600 9994 9720 10010
rect 9588 9988 9720 9994
rect 9640 9982 9720 9988
rect 9588 9930 9640 9936
rect 9692 9654 9720 9982
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 8666 9480 8722 9489
rect 8666 9415 8722 9424
rect 9678 9480 9734 9489
rect 9678 9415 9734 9424
rect 9692 9042 9720 9415
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 8022 8936 8078 8945
rect 8022 8871 8078 8880
rect 9784 7993 9812 12582
rect 9876 12458 9904 18566
rect 9968 17338 9996 18686
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10060 17218 10088 19615
rect 10152 19378 10180 21100
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10244 20641 10272 20742
rect 10230 20632 10286 20641
rect 10230 20567 10286 20576
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10230 19544 10286 19553
rect 10230 19479 10286 19488
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10244 19156 10272 19479
rect 10152 19128 10272 19156
rect 10152 18737 10180 19128
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10138 18728 10194 18737
rect 10138 18663 10194 18672
rect 9968 17190 10088 17218
rect 9968 15706 9996 17190
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9968 15162 9996 15642
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9968 13394 9996 13738
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 12986 9996 13330
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 10060 12782 10088 17002
rect 10152 16590 10180 18663
rect 10244 18329 10272 18770
rect 10324 18760 10376 18766
rect 10508 18760 10560 18766
rect 10324 18702 10376 18708
rect 10506 18728 10508 18737
rect 10560 18728 10562 18737
rect 10336 18601 10364 18702
rect 10506 18663 10562 18672
rect 10322 18592 10378 18601
rect 10322 18527 10378 18536
rect 10230 18320 10286 18329
rect 10230 18255 10286 18264
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10244 17338 10272 17614
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 16250 10180 16526
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10324 15496 10376 15502
rect 10322 15464 10324 15473
rect 10376 15464 10378 15473
rect 10322 15399 10378 15408
rect 10336 15162 10364 15399
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10140 14816 10192 14822
rect 10138 14784 10140 14793
rect 10192 14784 10194 14793
rect 10138 14719 10194 14728
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9876 12430 9987 12458
rect 9959 12424 9987 12430
rect 9959 12396 9996 12424
rect 9968 9586 9996 12396
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11898 10088 12242
rect 10152 12238 10180 13806
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10060 11286 10088 11834
rect 10152 11354 10180 12174
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10046 10568 10102 10577
rect 10046 10503 10102 10512
rect 10140 10532 10192 10538
rect 10060 10305 10088 10503
rect 10140 10474 10192 10480
rect 10152 10441 10180 10474
rect 10704 10470 10732 21286
rect 10796 17882 10824 21644
rect 10888 21664 10966 21672
rect 11022 21664 11100 21672
rect 10888 21644 11100 21664
rect 10888 21554 10916 21644
rect 10966 21584 11022 21593
rect 10876 21548 10928 21554
rect 10966 21519 11022 21528
rect 10876 21490 10928 21496
rect 10980 21078 11008 21519
rect 10968 21072 11020 21078
rect 10874 21040 10930 21049
rect 10968 21014 11020 21020
rect 10874 20975 10876 20984
rect 10928 20975 10930 20984
rect 10876 20946 10928 20952
rect 11072 20942 11100 21644
rect 11164 21486 11192 22442
rect 11348 22098 11376 22607
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 11348 21554 11376 22034
rect 11440 21894 11468 24550
rect 11716 24410 11744 25366
rect 11794 24848 11850 24857
rect 11794 24783 11850 24792
rect 11704 24404 11756 24410
rect 11704 24346 11756 24352
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11520 23656 11572 23662
rect 11520 23598 11572 23604
rect 11532 23186 11560 23598
rect 11716 23508 11744 24142
rect 11808 23769 11836 24783
rect 11794 23760 11850 23769
rect 11794 23695 11850 23704
rect 11796 23520 11848 23526
rect 11716 23480 11796 23508
rect 11796 23462 11848 23468
rect 11808 23186 11836 23462
rect 11520 23180 11572 23186
rect 11520 23122 11572 23128
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11532 22778 11560 23122
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11532 22166 11560 22714
rect 11808 22574 11836 23122
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11520 22160 11572 22166
rect 11572 22120 11652 22148
rect 11520 22102 11572 22108
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11518 21856 11574 21865
rect 11518 21791 11574 21800
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11164 21146 11192 21422
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11060 20936 11112 20942
rect 10980 20896 11060 20924
rect 10980 20602 11008 20896
rect 11060 20878 11112 20884
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11150 20496 11206 20505
rect 11150 20431 11206 20440
rect 11058 20360 11114 20369
rect 11058 20295 11114 20304
rect 11072 20262 11100 20295
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10874 20088 10930 20097
rect 11164 20058 11192 20431
rect 10874 20023 10930 20032
rect 11152 20052 11204 20058
rect 10888 19553 10916 20023
rect 11152 19994 11204 20000
rect 10966 19816 11022 19825
rect 10966 19751 11022 19760
rect 10874 19544 10930 19553
rect 10874 19479 10930 19488
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10888 18970 10916 19314
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10796 17134 10824 17818
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10784 16992 10836 16998
rect 10782 16960 10784 16969
rect 10836 16960 10838 16969
rect 10782 16895 10838 16904
rect 10888 16590 10916 17818
rect 10980 16658 11008 19751
rect 11150 19680 11206 19689
rect 11150 19615 11206 19624
rect 11058 19272 11114 19281
rect 11058 19207 11114 19216
rect 11072 18970 11100 19207
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11072 17377 11100 18090
rect 11058 17368 11114 17377
rect 11058 17303 11114 17312
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10876 16584 10928 16590
rect 10796 16544 10876 16572
rect 10796 15502 10824 16544
rect 10876 16526 10928 16532
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10874 16280 10930 16289
rect 10980 16250 11008 16458
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11164 16402 11192 19615
rect 11440 19446 11468 21626
rect 11532 21321 11560 21791
rect 11624 21690 11652 22120
rect 11612 21684 11664 21690
rect 11900 21672 11928 27520
rect 12072 26104 12124 26110
rect 12072 26046 12124 26052
rect 11980 25832 12032 25838
rect 11978 25800 11980 25809
rect 12032 25800 12034 25809
rect 11978 25735 12034 25744
rect 12084 25498 12112 26046
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 11992 23254 12020 25094
rect 12084 24750 12112 25434
rect 12162 25392 12218 25401
rect 12162 25327 12218 25336
rect 12072 24744 12124 24750
rect 12072 24686 12124 24692
rect 12072 24336 12124 24342
rect 12072 24278 12124 24284
rect 12084 23905 12112 24278
rect 12070 23896 12126 23905
rect 12070 23831 12072 23840
rect 12124 23831 12126 23840
rect 12072 23802 12124 23808
rect 11980 23248 12032 23254
rect 11980 23190 12032 23196
rect 11612 21626 11664 21632
rect 11716 21644 11928 21672
rect 11518 21312 11574 21321
rect 11518 21247 11574 21256
rect 11518 21176 11574 21185
rect 11518 21111 11520 21120
rect 11572 21111 11574 21120
rect 11520 21082 11572 21088
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11624 20262 11652 20334
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11440 19174 11468 19382
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11348 17882 11376 18770
rect 11440 18766 11468 19110
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11440 18086 11468 18702
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 11336 17672 11388 17678
rect 11388 17620 11468 17626
rect 11336 17614 11468 17620
rect 11348 17598 11468 17614
rect 11334 17368 11390 17377
rect 11334 17303 11390 17312
rect 11348 17134 11376 17303
rect 11440 17202 11468 17598
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11440 16833 11468 17138
rect 11426 16824 11482 16833
rect 11426 16759 11428 16768
rect 11480 16759 11482 16768
rect 11428 16730 11480 16736
rect 11440 16699 11468 16730
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 10874 16215 10930 16224
rect 10968 16244 11020 16250
rect 10888 15706 10916 16215
rect 10968 16186 11020 16192
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10888 15314 10916 15642
rect 10980 15570 11008 16186
rect 11072 16182 11100 16390
rect 11164 16374 11284 16402
rect 11150 16280 11206 16289
rect 11150 16215 11206 16224
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11072 15978 11100 16118
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 11164 15337 11192 16215
rect 11150 15328 11206 15337
rect 10888 15286 11100 15314
rect 10782 15192 10838 15201
rect 10782 15127 10784 15136
rect 10836 15127 10838 15136
rect 10784 15098 10836 15104
rect 11072 15026 11100 15286
rect 11150 15263 11206 15272
rect 11060 15020 11112 15026
rect 11112 14980 11192 15008
rect 11060 14962 11112 14968
rect 11060 14272 11112 14278
rect 11164 14249 11192 14980
rect 11060 14214 11112 14220
rect 11150 14240 11206 14249
rect 11072 13870 11100 14214
rect 11150 14175 11206 14184
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10980 13394 11008 13670
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10980 12986 11008 13330
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10782 12336 10838 12345
rect 10782 12271 10838 12280
rect 10796 11898 10824 12271
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10874 11112 10930 11121
rect 10874 11047 10876 11056
rect 10928 11047 10930 11056
rect 10876 11018 10928 11024
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10692 10464 10744 10470
rect 10138 10432 10194 10441
rect 10692 10406 10744 10412
rect 10138 10367 10194 10376
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10046 10296 10102 10305
rect 10289 10288 10585 10308
rect 10046 10231 10102 10240
rect 10692 10260 10744 10266
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 10060 9518 10088 10231
rect 10692 10202 10744 10208
rect 10704 9586 10732 10202
rect 10796 10198 10824 10950
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10888 10010 10916 10406
rect 10980 10266 11008 12922
rect 11256 12458 11284 16374
rect 11348 16017 11376 16594
rect 11532 16538 11560 19654
rect 11624 17921 11652 20198
rect 11716 19786 11744 21644
rect 11794 21584 11850 21593
rect 11794 21519 11850 21528
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11808 19310 11836 21519
rect 12070 21312 12126 21321
rect 12070 21247 12126 21256
rect 11886 20496 11942 20505
rect 11886 20431 11942 20440
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11610 17912 11666 17921
rect 11610 17847 11666 17856
rect 11440 16510 11560 16538
rect 11334 16008 11390 16017
rect 11334 15943 11390 15952
rect 11348 15706 11376 15943
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11440 15586 11468 16510
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11164 12430 11284 12458
rect 11348 15558 11468 15586
rect 11164 12424 11192 12430
rect 11072 12396 11192 12424
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10796 9982 10916 10010
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9864 9376 9916 9382
rect 9862 9344 9864 9353
rect 9916 9344 9918 9353
rect 9862 9279 9918 9288
rect 9968 9217 9996 9386
rect 9954 9208 10010 9217
rect 10060 9178 10088 9454
rect 9954 9143 10010 9152
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9770 7984 9826 7993
rect 9770 7919 9826 7928
rect 7470 7576 7526 7585
rect 7470 7511 7526 7520
rect 10152 7449 10180 9522
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10138 7440 10194 7449
rect 10138 7375 10194 7384
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10796 6905 10824 9982
rect 10980 9178 11008 10066
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10782 6896 10838 6905
rect 10782 6831 10838 6840
rect 4066 6760 4122 6769
rect 4066 6695 4122 6704
rect 4080 6089 4108 6695
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 4066 6080 4122 6089
rect 4066 6015 4122 6024
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 4066 5400 4122 5409
rect 5622 5392 5918 5412
rect 4066 5335 4122 5344
rect 3974 5264 4030 5273
rect 3974 5199 4030 5208
rect 3882 4856 3938 4865
rect 3882 4791 3938 4800
rect 3988 4321 4016 5199
rect 4080 4729 4108 5335
rect 10690 4992 10746 5001
rect 10289 4924 10585 4944
rect 10690 4927 10746 4936
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 4066 4720 4122 4729
rect 4066 4655 4122 4664
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 3974 4312 4030 4321
rect 5622 4304 5918 4324
rect 3974 4247 4030 4256
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3505 10732 4927
rect 11072 3505 11100 12396
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11150 11792 11206 11801
rect 11256 11762 11284 12038
rect 11150 11727 11206 11736
rect 11244 11756 11296 11762
rect 11164 11694 11192 11727
rect 11244 11698 11296 11704
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11256 11354 11284 11698
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11164 10742 11192 11222
rect 11242 11112 11298 11121
rect 11242 11047 11298 11056
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11256 10674 11284 11047
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9654 11284 9998
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11348 8498 11376 15558
rect 11532 14482 11560 15846
rect 11624 15065 11652 17847
rect 11808 17542 11836 18022
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11808 17338 11836 17478
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 15638 11744 16390
rect 11808 16250 11836 17274
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11610 15056 11666 15065
rect 11716 15026 11744 15574
rect 11808 15162 11836 16186
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11610 14991 11666 15000
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11716 14618 11744 14962
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11532 14074 11560 14418
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11440 12306 11468 13126
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11624 12442 11652 12650
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11520 12232 11572 12238
rect 11426 12200 11482 12209
rect 11520 12174 11572 12180
rect 11426 12135 11428 12144
rect 11480 12135 11482 12144
rect 11428 12106 11480 12112
rect 11440 11762 11468 12106
rect 11532 12102 11560 12174
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11532 11898 11560 12038
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11624 10674 11652 12378
rect 11900 12073 11928 20431
rect 12084 17218 12112 21247
rect 12176 21146 12204 25327
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12268 23905 12296 24006
rect 12254 23896 12310 23905
rect 12254 23831 12310 23840
rect 12452 22234 12480 25638
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12256 22160 12308 22166
rect 12256 22102 12308 22108
rect 12268 21690 12296 22102
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12360 21146 12388 21830
rect 12544 21298 12572 27520
rect 12808 25832 12860 25838
rect 12806 25800 12808 25809
rect 12860 25800 12862 25809
rect 12806 25735 12862 25744
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12820 24614 12848 25298
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 12912 24886 12940 25230
rect 12900 24880 12952 24886
rect 12900 24822 12952 24828
rect 12912 24721 12940 24822
rect 12992 24744 13044 24750
rect 12898 24712 12954 24721
rect 12992 24686 13044 24692
rect 12898 24647 12954 24656
rect 12808 24608 12860 24614
rect 13004 24596 13032 24686
rect 12808 24550 12860 24556
rect 12912 24568 13032 24596
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12728 24177 12756 24210
rect 12808 24200 12860 24206
rect 12714 24168 12770 24177
rect 12808 24142 12860 24148
rect 12714 24103 12770 24112
rect 12728 23866 12756 24103
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12820 23769 12848 24142
rect 12806 23760 12862 23769
rect 12806 23695 12862 23704
rect 12912 23644 12940 24568
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 13004 23662 13032 24006
rect 12820 23616 12940 23644
rect 12992 23656 13044 23662
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12636 22137 12664 22374
rect 12622 22128 12678 22137
rect 12622 22063 12678 22072
rect 12624 21480 12676 21486
rect 12622 21448 12624 21457
rect 12676 21448 12678 21457
rect 12622 21383 12678 21392
rect 12544 21270 12664 21298
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12532 21140 12584 21146
rect 12532 21082 12584 21088
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12268 20210 12296 20334
rect 12360 20330 12388 20878
rect 12348 20324 12400 20330
rect 12348 20266 12400 20272
rect 12268 20182 12388 20210
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12268 19174 12296 19858
rect 12360 19718 12388 20182
rect 12452 19786 12480 20946
rect 12544 20398 12572 21082
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 12360 19242 12388 19654
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12268 18873 12296 19110
rect 12254 18864 12310 18873
rect 12254 18799 12310 18808
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12176 18465 12204 18566
rect 12162 18456 12218 18465
rect 12162 18391 12218 18400
rect 12176 17746 12204 18391
rect 12268 18057 12296 18799
rect 12440 18080 12492 18086
rect 12254 18048 12310 18057
rect 12440 18022 12492 18028
rect 12254 17983 12310 17992
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12176 17338 12204 17682
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12452 17241 12480 18022
rect 12438 17232 12494 17241
rect 12084 17190 12296 17218
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12084 13190 12112 14418
rect 12162 13832 12218 13841
rect 12162 13767 12164 13776
rect 12216 13767 12218 13776
rect 12164 13738 12216 13744
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11886 12064 11942 12073
rect 11886 11999 11942 12008
rect 11702 11928 11758 11937
rect 11702 11863 11758 11872
rect 11716 11150 11744 11863
rect 12084 11257 12112 13126
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12176 11665 12204 12242
rect 12162 11656 12218 11665
rect 12162 11591 12164 11600
rect 12216 11591 12218 11600
rect 12164 11562 12216 11568
rect 12268 11286 12296 17190
rect 12438 17167 12494 17176
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12452 15910 12480 17070
rect 12544 16289 12572 19110
rect 12636 18426 12664 21270
rect 12728 20942 12756 22510
rect 12716 20936 12768 20942
rect 12820 20913 12848 23616
rect 12992 23598 13044 23604
rect 12900 23316 12952 23322
rect 12900 23258 12952 23264
rect 12912 22166 12940 23258
rect 13004 23118 13032 23598
rect 13096 23202 13124 27520
rect 13452 27056 13504 27062
rect 13452 26998 13504 27004
rect 13268 25424 13320 25430
rect 13268 25366 13320 25372
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 13188 24818 13216 25230
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13188 23322 13216 24754
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 13096 23174 13216 23202
rect 12992 23112 13044 23118
rect 12992 23054 13044 23060
rect 13004 22710 13032 23054
rect 12992 22704 13044 22710
rect 12992 22646 13044 22652
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12912 21418 12940 21830
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 12716 20878 12768 20884
rect 12806 20904 12862 20913
rect 12728 19990 12756 20878
rect 12806 20839 12862 20848
rect 12716 19984 12768 19990
rect 12716 19926 12768 19932
rect 12806 18728 12862 18737
rect 12806 18663 12862 18672
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12636 18222 12664 18362
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12714 18184 12770 18193
rect 12714 18119 12770 18128
rect 12728 17270 12756 18119
rect 12820 17882 12848 18663
rect 12898 18320 12954 18329
rect 12898 18255 12954 18264
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 12530 16280 12586 16289
rect 12530 16215 12586 16224
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15638 12480 15846
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12728 15162 12756 17206
rect 12912 16794 12940 18255
rect 13188 17377 13216 23174
rect 13174 17368 13230 17377
rect 13280 17338 13308 25366
rect 13464 24750 13492 26998
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13372 24313 13400 24550
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13358 24304 13414 24313
rect 13358 24239 13414 24248
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 13372 21146 13400 21422
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13464 20874 13492 24346
rect 13544 23588 13596 23594
rect 13544 23530 13596 23536
rect 13556 23089 13584 23530
rect 13542 23080 13598 23089
rect 13542 23015 13544 23024
rect 13596 23015 13598 23024
rect 13544 22986 13596 22992
rect 13556 22681 13584 22986
rect 13648 22953 13676 27520
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13726 23488 13782 23497
rect 13726 23423 13782 23432
rect 13634 22944 13690 22953
rect 13634 22879 13690 22888
rect 13542 22672 13598 22681
rect 13542 22607 13598 22616
rect 13648 22409 13676 22879
rect 13634 22400 13690 22409
rect 13634 22335 13690 22344
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 13740 20058 13768 23423
rect 13820 22976 13872 22982
rect 13820 22918 13872 22924
rect 13832 22574 13860 22918
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13358 19952 13414 19961
rect 13358 19887 13414 19896
rect 13372 19718 13400 19887
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13372 19174 13400 19654
rect 13832 19394 13860 20198
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13648 19366 13860 19394
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13556 18834 13584 19314
rect 13648 18902 13676 19366
rect 13818 19272 13874 19281
rect 13818 19207 13874 19216
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13450 18320 13506 18329
rect 13450 18255 13452 18264
rect 13504 18255 13506 18264
rect 13636 18284 13688 18290
rect 13452 18226 13504 18232
rect 13636 18226 13688 18232
rect 13360 17808 13412 17814
rect 13358 17776 13360 17785
rect 13412 17776 13414 17785
rect 13358 17711 13414 17720
rect 13648 17338 13676 18226
rect 13174 17303 13230 17312
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12820 15706 12848 16118
rect 13004 15978 13032 16526
rect 13634 16280 13690 16289
rect 13634 16215 13690 16224
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12346 14784 12402 14793
rect 12346 14719 12402 14728
rect 12360 14618 12388 14719
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12544 13870 12572 15098
rect 13280 15026 13308 15506
rect 13372 15366 13400 15846
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13372 15201 13400 15302
rect 13358 15192 13414 15201
rect 13358 15127 13414 15136
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 14278 12756 14758
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 12753 12480 13670
rect 12544 13394 12572 13806
rect 12728 13734 12756 14214
rect 13004 14074 13032 14350
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13004 13977 13032 14010
rect 13188 13977 13216 14826
rect 13280 14618 13308 14962
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13372 14113 13400 14418
rect 13464 14278 13492 14826
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13358 14104 13414 14113
rect 13358 14039 13360 14048
rect 13412 14039 13414 14048
rect 13360 14010 13412 14016
rect 13372 13979 13400 14010
rect 12990 13968 13046 13977
rect 12990 13903 13046 13912
rect 13174 13968 13230 13977
rect 13174 13903 13230 13912
rect 13464 13870 13492 14214
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13542 13832 13598 13841
rect 13542 13767 13598 13776
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12544 13274 12572 13330
rect 12544 13246 12664 13274
rect 12438 12744 12494 12753
rect 12438 12679 12494 12688
rect 12636 12646 12664 13246
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12102 12664 12582
rect 12728 12458 12756 13670
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12719 12430 12756 12458
rect 12912 12442 12940 13398
rect 13450 13288 13506 13297
rect 13450 13223 13506 13232
rect 13464 12782 13492 13223
rect 13556 12986 13584 13767
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13542 12880 13598 12889
rect 13542 12815 13598 12824
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13556 12714 13584 12815
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13556 12442 13584 12650
rect 12900 12436 12952 12442
rect 12719 12356 12747 12430
rect 12900 12378 12952 12384
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 12719 12328 12756 12356
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12636 11694 12664 12038
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12256 11280 12308 11286
rect 12070 11248 12126 11257
rect 11796 11212 11848 11218
rect 12256 11222 12308 11228
rect 12070 11183 12126 11192
rect 11796 11154 11848 11160
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 10266 11652 10610
rect 11808 10470 11836 11154
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9382 11560 10066
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 8022 11284 8230
rect 11532 8090 11560 9318
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11256 7546 11284 7958
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 10690 3496 10746 3505
rect 10690 3431 10746 3440
rect 11058 3496 11114 3505
rect 11058 3431 11114 3440
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 3252 2910 3464 2938
rect 3146 912 3202 921
rect 3146 847 3202 856
rect 3252 377 3280 2910
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 3514 2680 3570 2689
rect 10289 2672 10585 2692
rect 3514 2615 3570 2624
rect 3528 1601 3556 2615
rect 4618 2408 4674 2417
rect 4618 2343 4674 2352
rect 3514 1592 3570 1601
rect 3514 1527 3570 1536
rect 4632 480 4660 2343
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 11808 1601 11836 10406
rect 12176 10130 12204 10746
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12176 9722 12204 10066
rect 12268 9761 12296 11222
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12452 10282 12480 11154
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12544 10606 12572 10950
rect 12636 10810 12664 11630
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12360 10254 12480 10282
rect 12360 9926 12388 10254
rect 12544 9926 12572 10542
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12254 9752 12310 9761
rect 12164 9716 12216 9722
rect 12254 9687 12310 9696
rect 12164 9658 12216 9664
rect 12544 9654 12572 9862
rect 12532 9648 12584 9654
rect 12728 9636 12756 12328
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13188 11150 13216 11562
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12532 9590 12584 9596
rect 12636 9608 12756 9636
rect 12348 9376 12400 9382
rect 12070 9344 12126 9353
rect 12348 9318 12400 9324
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12070 9279 12126 9288
rect 12084 9178 12112 9279
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12084 9058 12112 9114
rect 11992 9030 12112 9058
rect 11992 8362 12020 9030
rect 12360 8906 12388 9318
rect 12544 9042 12572 9318
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 7206 11928 7890
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11900 3641 11928 7142
rect 11886 3632 11942 3641
rect 11886 3567 11942 3576
rect 11992 2553 12020 8298
rect 12360 8022 12388 8842
rect 12544 8634 12572 8978
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12348 8016 12400 8022
rect 12162 7984 12218 7993
rect 12348 7958 12400 7964
rect 12162 7919 12218 7928
rect 12176 7886 12204 7919
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12636 6361 12664 9608
rect 12820 8514 12848 9658
rect 12912 8634 12940 11086
rect 13542 10432 13598 10441
rect 13542 10367 13598 10376
rect 13266 10296 13322 10305
rect 13266 10231 13322 10240
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13280 8537 13308 10231
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8566 13400 8774
rect 13360 8560 13412 8566
rect 13266 8528 13322 8537
rect 12820 8486 12940 8514
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12728 7342 12756 7754
rect 12716 7336 12768 7342
rect 12714 7304 12716 7313
rect 12768 7304 12770 7313
rect 12714 7239 12770 7248
rect 12622 6352 12678 6361
rect 12622 6287 12678 6296
rect 11978 2544 12034 2553
rect 11978 2479 12034 2488
rect 12912 2446 12940 8486
rect 13360 8502 13412 8508
rect 13266 8463 13322 8472
rect 13372 8430 13400 8502
rect 13464 8498 13492 9862
rect 13556 8906 13584 10367
rect 13648 10169 13676 16215
rect 13740 15745 13768 19110
rect 13832 18970 13860 19207
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13818 18592 13874 18601
rect 13818 18527 13874 18536
rect 13832 17882 13860 18527
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16794 13860 17070
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13832 16425 13860 16730
rect 13818 16416 13874 16425
rect 13818 16351 13874 16360
rect 13820 16040 13872 16046
rect 13818 16008 13820 16017
rect 13872 16008 13874 16017
rect 13818 15943 13874 15952
rect 13726 15736 13782 15745
rect 13726 15671 13782 15680
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13832 14618 13860 15302
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 13410 13768 14350
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13832 13530 13860 13738
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13740 13382 13860 13410
rect 13726 13288 13782 13297
rect 13726 13223 13782 13232
rect 13740 12850 13768 13223
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13832 11234 13860 13382
rect 13924 11336 13952 24006
rect 14016 23526 14044 24550
rect 14292 24426 14320 27520
rect 14844 26246 14872 27520
rect 15396 27062 15424 27520
rect 15384 27056 15436 27062
rect 15384 26998 15436 27004
rect 14832 26240 14884 26246
rect 14832 26182 14884 26188
rect 15476 25424 15528 25430
rect 15474 25392 15476 25401
rect 15528 25392 15530 25401
rect 16040 25378 16068 27520
rect 14464 25356 14516 25362
rect 15474 25327 15530 25336
rect 15580 25350 16068 25378
rect 14464 25298 14516 25304
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14108 24398 14320 24426
rect 14108 23594 14136 24398
rect 14278 24168 14334 24177
rect 14278 24103 14280 24112
rect 14332 24103 14334 24112
rect 14280 24074 14332 24080
rect 14096 23588 14148 23594
rect 14096 23530 14148 23536
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 14016 16250 14044 22918
rect 14108 22545 14136 23530
rect 14278 23352 14334 23361
rect 14278 23287 14334 23296
rect 14094 22536 14150 22545
rect 14094 22471 14150 22480
rect 14188 22500 14240 22506
rect 14188 22442 14240 22448
rect 14200 22166 14228 22442
rect 14188 22160 14240 22166
rect 14188 22102 14240 22108
rect 14094 21720 14150 21729
rect 14200 21706 14228 22102
rect 14292 21962 14320 23287
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 14150 21690 14228 21706
rect 14150 21684 14240 21690
rect 14150 21678 14188 21684
rect 14094 21655 14150 21664
rect 14188 21626 14240 21632
rect 14384 21486 14412 24618
rect 14476 24070 14504 25298
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15304 24936 15332 25162
rect 15212 24908 15332 24936
rect 15212 24818 15240 24908
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 14556 24676 14608 24682
rect 14556 24618 14608 24624
rect 15384 24676 15436 24682
rect 15384 24618 15436 24624
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14476 22166 14504 24006
rect 14464 22160 14516 22166
rect 14464 22102 14516 22108
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14280 21072 14332 21078
rect 14568 21049 14596 24618
rect 14648 24268 14700 24274
rect 14648 24210 14700 24216
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 14660 22982 14688 24210
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14752 23905 14780 24142
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14738 23896 14794 23905
rect 14956 23888 15252 23908
rect 14738 23831 14740 23840
rect 14792 23831 14794 23840
rect 14740 23802 14792 23808
rect 15304 23594 15332 24210
rect 15396 24138 15424 24618
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15384 24132 15436 24138
rect 15384 24074 15436 24080
rect 15384 23724 15436 23730
rect 15384 23666 15436 23672
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14660 22778 14688 22918
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14280 21014 14332 21020
rect 14554 21040 14610 21049
rect 14292 20602 14320 21014
rect 14554 20975 14610 20984
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14280 20596 14332 20602
rect 14200 20556 14280 20584
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14108 19242 14136 19790
rect 14200 19417 14228 20556
rect 14280 20538 14332 20544
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14186 19408 14242 19417
rect 14186 19343 14242 19352
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14108 18902 14136 19178
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14094 18728 14150 18737
rect 14094 18663 14150 18672
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14108 15910 14136 18663
rect 14200 18426 14228 19246
rect 14292 19242 14320 19790
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14384 19122 14412 20742
rect 14568 20058 14596 20975
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14462 19272 14518 19281
rect 14462 19207 14518 19216
rect 14292 19094 14412 19122
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14186 16416 14242 16425
rect 14186 16351 14242 16360
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 14016 14822 14044 15506
rect 14094 15464 14150 15473
rect 14094 15399 14096 15408
rect 14148 15399 14150 15408
rect 14096 15370 14148 15376
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14016 13433 14044 14758
rect 14200 14414 14228 16351
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14200 13530 14228 14350
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14002 13424 14058 13433
rect 14002 13359 14058 13368
rect 14186 13424 14242 13433
rect 14186 13359 14242 13368
rect 14002 12880 14058 12889
rect 14002 12815 14058 12824
rect 14016 12782 14044 12815
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14200 12714 14228 13359
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14200 11393 14228 12174
rect 14186 11384 14242 11393
rect 13924 11308 14136 11336
rect 14292 11354 14320 19094
rect 14370 16688 14426 16697
rect 14370 16623 14372 16632
rect 14424 16623 14426 16632
rect 14372 16594 14424 16600
rect 14384 16046 14412 16594
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14476 15994 14504 19207
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18222 14596 19110
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14568 17882 14596 18158
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14568 16114 14596 16934
rect 14660 16153 14688 21966
rect 14752 21894 14780 23122
rect 15396 23118 15424 23666
rect 15384 23112 15436 23118
rect 15290 23080 15346 23089
rect 14832 23044 14884 23050
rect 15384 23054 15436 23060
rect 15290 23015 15346 23024
rect 14832 22986 14884 22992
rect 14844 22545 14872 22986
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22778 15332 23015
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 15290 22672 15346 22681
rect 15290 22607 15346 22616
rect 14830 22536 14886 22545
rect 14830 22471 14886 22480
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14646 16144 14702 16153
rect 14556 16108 14608 16114
rect 14646 16079 14702 16088
rect 14556 16050 14608 16056
rect 14476 15966 14596 15994
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14384 15201 14412 15846
rect 14476 15366 14504 15846
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14370 15192 14426 15201
rect 14370 15127 14426 15136
rect 14186 11319 14242 11328
rect 14280 11348 14332 11354
rect 13832 11206 13952 11234
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13832 10810 13860 11086
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13634 10160 13690 10169
rect 13634 10095 13690 10104
rect 13728 9172 13780 9178
rect 13832 9160 13860 10474
rect 13780 9132 13860 9160
rect 13728 9114 13780 9120
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13464 8090 13492 8434
rect 13740 8362 13768 9114
rect 13924 9042 13952 11206
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13832 8129 13860 8978
rect 13924 8634 13952 8978
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13818 8120 13874 8129
rect 13740 8090 13818 8106
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13728 8084 13818 8090
rect 13780 8078 13818 8084
rect 14108 8090 14136 11308
rect 14280 11290 14332 11296
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14200 10266 14228 11018
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14186 10024 14242 10033
rect 14186 9959 14242 9968
rect 13818 8055 13874 8064
rect 14096 8084 14148 8090
rect 13728 8026 13780 8032
rect 13832 7995 13860 8055
rect 14096 8026 14148 8032
rect 14200 7721 14228 9959
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14292 8974 14320 9386
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 7750 14320 8910
rect 14280 7744 14332 7750
rect 14186 7712 14242 7721
rect 14280 7686 14332 7692
rect 14186 7647 14242 7656
rect 14292 2650 14320 7686
rect 14384 6769 14412 15127
rect 14568 15042 14596 15966
rect 14476 15014 14596 15042
rect 14476 14793 14504 15014
rect 14556 14884 14608 14890
rect 14556 14826 14608 14832
rect 14462 14784 14518 14793
rect 14462 14719 14518 14728
rect 14462 14512 14518 14521
rect 14462 14447 14464 14456
rect 14516 14447 14518 14456
rect 14464 14418 14516 14424
rect 14568 14278 14596 14826
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14646 14240 14702 14249
rect 14568 14006 14596 14214
rect 14646 14175 14702 14184
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14476 12102 14504 12786
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11830 14504 12038
rect 14568 11937 14596 13942
rect 14554 11928 14610 11937
rect 14554 11863 14610 11872
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14554 9752 14610 9761
rect 14554 9687 14610 9696
rect 14568 9110 14596 9687
rect 14660 9178 14688 14175
rect 14752 10713 14780 21830
rect 14844 21672 14872 21898
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14844 21644 14964 21672
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14844 20913 14872 20946
rect 14830 20904 14886 20913
rect 14936 20874 14964 21644
rect 15304 21350 15332 22607
rect 15488 22103 15516 24550
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15474 22094 15530 22103
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 14830 20839 14886 20848
rect 14924 20868 14976 20874
rect 14844 20602 14872 20839
rect 14924 20810 14976 20816
rect 15396 20806 15424 22034
rect 15474 22029 15530 22038
rect 15580 21978 15608 25350
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 16592 25242 16620 27520
rect 16948 25424 17000 25430
rect 16948 25366 17000 25372
rect 15658 24848 15714 24857
rect 15658 24783 15714 24792
rect 15488 21950 15608 21978
rect 15384 20800 15436 20806
rect 15382 20768 15384 20777
rect 15436 20768 15438 20777
rect 14956 20700 15252 20720
rect 15382 20703 15438 20712
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 15488 20097 15516 21950
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15580 21554 15608 21830
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15672 21146 15700 24783
rect 15948 24614 15976 25230
rect 16132 24886 16160 25230
rect 16592 25214 16712 25242
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16120 24880 16172 24886
rect 16120 24822 16172 24828
rect 16592 24750 16620 25094
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15842 24440 15898 24449
rect 15842 24375 15898 24384
rect 15752 24132 15804 24138
rect 15752 24074 15804 24080
rect 15764 23594 15792 24074
rect 15752 23588 15804 23594
rect 15752 23530 15804 23536
rect 15764 22681 15792 23530
rect 15750 22672 15806 22681
rect 15750 22607 15806 22616
rect 15750 21992 15806 22001
rect 15856 21962 15884 24375
rect 15750 21927 15806 21936
rect 15844 21956 15896 21962
rect 15764 21457 15792 21927
rect 15844 21898 15896 21904
rect 15750 21448 15806 21457
rect 15750 21383 15806 21392
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15474 20088 15530 20097
rect 15474 20023 15530 20032
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14844 19310 14872 19654
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19514 15332 19858
rect 15764 19854 15792 21383
rect 15948 21146 15976 24550
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 16040 22778 16068 23054
rect 16028 22772 16080 22778
rect 16080 22732 16160 22760
rect 16028 22714 16080 22720
rect 16028 21888 16080 21894
rect 16028 21830 16080 21836
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15856 20058 15884 20946
rect 16040 20806 16068 21830
rect 16132 21010 16160 22732
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 16040 20398 16068 20742
rect 16132 20602 16160 20946
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16028 20392 16080 20398
rect 16028 20334 16080 20340
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 14832 19304 14884 19310
rect 14832 19246 14884 19252
rect 14844 18834 14872 19246
rect 15304 18970 15332 19450
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 15488 18630 15516 19790
rect 15856 19378 15884 19994
rect 16224 19825 16252 24006
rect 16316 22982 16344 24142
rect 16394 23760 16450 23769
rect 16394 23695 16450 23704
rect 16408 23254 16436 23695
rect 16684 23361 16712 25214
rect 16856 24880 16908 24886
rect 16856 24822 16908 24828
rect 16762 24712 16818 24721
rect 16762 24647 16818 24656
rect 16776 24614 16804 24647
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 16868 24410 16896 24822
rect 16960 24750 16988 25366
rect 17144 24857 17172 27520
rect 17500 25968 17552 25974
rect 17500 25910 17552 25916
rect 17224 25696 17276 25702
rect 17224 25638 17276 25644
rect 17130 24848 17186 24857
rect 17130 24783 17186 24792
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 17038 24576 17094 24585
rect 17038 24511 17094 24520
rect 17052 24410 17080 24511
rect 17236 24410 17264 25638
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 17040 24404 17092 24410
rect 17040 24346 17092 24352
rect 17224 24404 17276 24410
rect 17224 24346 17276 24352
rect 16856 23792 16908 23798
rect 16854 23760 16856 23769
rect 16908 23760 16910 23769
rect 16854 23695 16910 23704
rect 16670 23352 16726 23361
rect 16670 23287 16726 23296
rect 16396 23248 16448 23254
rect 16396 23190 16448 23196
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16408 22522 16436 23190
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16316 22494 16436 22522
rect 16488 22500 16540 22506
rect 16316 22234 16344 22494
rect 16488 22442 16540 22448
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16304 21480 16356 21486
rect 16304 21422 16356 21428
rect 16316 21321 16344 21422
rect 16302 21312 16358 21321
rect 16302 21247 16358 21256
rect 16316 21146 16344 21247
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 16408 19904 16436 22374
rect 16500 21690 16528 22442
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16776 21962 16804 22374
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16488 21412 16540 21418
rect 16540 21372 16620 21400
rect 16488 21354 16540 21360
rect 16592 20058 16620 21372
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16776 21049 16804 21286
rect 16762 21040 16818 21049
rect 16762 20975 16818 20984
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16580 19916 16632 19922
rect 16408 19876 16580 19904
rect 16580 19858 16632 19864
rect 16776 19854 16804 20198
rect 16764 19848 16816 19854
rect 16210 19816 16266 19825
rect 16764 19790 16816 19796
rect 16210 19751 16266 19760
rect 16394 19680 16450 19689
rect 16394 19615 16450 19624
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14844 16250 14872 17614
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 17218 15332 18022
rect 15382 17640 15438 17649
rect 15382 17575 15384 17584
rect 15436 17575 15438 17584
rect 15384 17546 15436 17552
rect 15120 17190 15332 17218
rect 15120 17134 15148 17190
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15290 17096 15346 17105
rect 15290 17031 15346 17040
rect 15304 16794 15332 17031
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15106 16688 15162 16697
rect 15106 16623 15108 16632
rect 15160 16623 15162 16632
rect 15108 16594 15160 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14738 10704 14794 10713
rect 14738 10639 14794 10648
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14568 8430 14596 9046
rect 14752 8906 14780 9658
rect 14844 8922 14872 12854
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11801 15332 15438
rect 15384 13864 15436 13870
rect 15382 13832 15384 13841
rect 15436 13832 15438 13841
rect 15382 13767 15438 13776
rect 15488 13682 15516 18566
rect 15568 18148 15620 18154
rect 15568 18090 15620 18096
rect 15396 13654 15516 13682
rect 15396 12753 15424 13654
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15488 12782 15516 13126
rect 15476 12776 15528 12782
rect 15382 12744 15438 12753
rect 15476 12718 15528 12724
rect 15382 12679 15438 12688
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15290 11792 15346 11801
rect 15290 11727 15346 11736
rect 15292 11552 15344 11558
rect 15396 11540 15424 12242
rect 15488 11898 15516 12718
rect 15580 12646 15608 18090
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15764 16250 15792 17682
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 16697 15884 17614
rect 15842 16688 15898 16697
rect 15842 16623 15898 16632
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15658 15328 15714 15337
rect 15658 15263 15714 15272
rect 15672 12714 15700 15263
rect 15948 13818 15976 19246
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16316 18426 16344 18770
rect 16408 18766 16436 19615
rect 16776 19514 16804 19790
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16868 18970 16896 23122
rect 17406 23080 17462 23089
rect 17406 23015 17408 23024
rect 17460 23015 17462 23024
rect 17408 22986 17460 22992
rect 17512 22778 17540 25910
rect 17788 25498 17816 27520
rect 18144 26036 18196 26042
rect 18144 25978 18196 25984
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17684 25356 17736 25362
rect 17684 25298 17736 25304
rect 17696 24614 17724 25298
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18064 24750 18092 25094
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17684 24608 17736 24614
rect 17684 24550 17736 24556
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17604 23662 17632 24210
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 17696 23304 17724 24550
rect 17868 24132 17920 24138
rect 17868 24074 17920 24080
rect 17774 23624 17830 23633
rect 17774 23559 17776 23568
rect 17828 23559 17830 23568
rect 17776 23530 17828 23536
rect 17880 23338 17908 24074
rect 18064 23497 18092 24686
rect 18156 24410 18184 25978
rect 18340 25514 18368 27520
rect 18248 25486 18368 25514
rect 18248 24449 18276 25486
rect 18892 25378 18920 27520
rect 19064 25764 19116 25770
rect 19064 25706 19116 25712
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 18708 25350 18920 25378
rect 18340 24954 18368 25298
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18234 24440 18290 24449
rect 18144 24404 18196 24410
rect 18234 24375 18290 24384
rect 18144 24346 18196 24352
rect 18156 23662 18184 24346
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18050 23488 18106 23497
rect 18050 23423 18106 23432
rect 17880 23310 18000 23338
rect 17696 23276 17816 23304
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 16960 21894 16988 22578
rect 17132 22160 17184 22166
rect 17132 22102 17184 22108
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 17144 21418 17172 22102
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 17328 21350 17356 22034
rect 17408 22024 17460 22030
rect 17406 21992 17408 22001
rect 17460 21992 17462 22001
rect 17406 21927 17462 21936
rect 17420 21554 17448 21927
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16960 19990 16988 21014
rect 17130 20768 17186 20777
rect 17130 20703 17186 20712
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16856 18760 16908 18766
rect 16960 18714 16988 19110
rect 16908 18708 16988 18714
rect 16856 18702 16988 18708
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16408 18154 16436 18702
rect 16868 18686 16988 18702
rect 16580 18624 16632 18630
rect 16500 18584 16580 18612
rect 16396 18148 16448 18154
rect 16396 18090 16448 18096
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 16040 17338 16068 17614
rect 16500 17338 16528 18584
rect 16580 18566 16632 18572
rect 16762 17912 16818 17921
rect 16762 17847 16818 17856
rect 16580 17536 16632 17542
rect 16776 17513 16804 17847
rect 16960 17542 16988 18686
rect 17052 17746 17080 19314
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 16948 17536 17000 17542
rect 16580 17478 16632 17484
rect 16762 17504 16818 17513
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16592 17066 16620 17478
rect 16948 17478 17000 17484
rect 16762 17439 16818 17448
rect 16776 17134 16804 17439
rect 16960 17202 16988 17478
rect 17052 17338 17080 17682
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16118 16144 16174 16153
rect 16118 16079 16174 16088
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 16040 13938 16068 14214
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 15856 13790 15976 13818
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15580 11830 15608 12242
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15344 11512 15424 11540
rect 15292 11494 15344 11500
rect 15304 11218 15332 11494
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 15028 10266 15056 10610
rect 15290 10568 15346 10577
rect 15290 10503 15292 10512
rect 15344 10503 15346 10512
rect 15292 10474 15344 10480
rect 15384 10464 15436 10470
rect 15382 10432 15384 10441
rect 15436 10432 15438 10441
rect 15382 10367 15438 10376
rect 15580 10266 15608 11222
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 10202
rect 15672 10033 15700 11290
rect 15764 11257 15792 13262
rect 15750 11248 15806 11257
rect 15750 11183 15806 11192
rect 15856 11132 15884 13790
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15948 12782 15976 13670
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15948 11354 15976 12582
rect 16040 11830 16068 13874
rect 16132 12866 16160 16079
rect 16224 15910 16252 16526
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 15502 16252 15846
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16224 14958 16252 15438
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16224 14482 16252 14894
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16224 14006 16252 14418
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16316 13190 16344 13670
rect 16408 13462 16436 14758
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16500 14074 16528 14418
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16396 13456 16448 13462
rect 16396 13398 16448 13404
rect 16304 13184 16356 13190
rect 16302 13152 16304 13161
rect 16356 13152 16358 13161
rect 16302 13087 16358 13096
rect 16408 12986 16436 13398
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16132 12838 16436 12866
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16040 11286 16068 11766
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15764 11104 15884 11132
rect 15658 10024 15714 10033
rect 15658 9959 15714 9968
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 14740 8900 14792 8906
rect 14844 8894 15332 8922
rect 14740 8842 14792 8848
rect 14752 8498 14780 8842
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 7993 14596 8366
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14554 7984 14610 7993
rect 14554 7919 14610 7928
rect 14370 6760 14426 6769
rect 14370 6695 14426 6704
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 11980 2440 12032 2446
rect 11978 2408 11980 2417
rect 12900 2440 12952 2446
rect 12032 2408 12034 2417
rect 12900 2382 12952 2388
rect 11978 2343 12034 2352
rect 13740 2258 13768 2450
rect 13740 2230 13952 2258
rect 11794 1592 11850 1601
rect 11794 1527 11850 1536
rect 13924 480 13952 2230
rect 14660 1601 14688 8298
rect 14752 8090 14780 8434
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14738 7576 14794 7585
rect 14844 7546 14872 8502
rect 15106 8256 15162 8265
rect 15106 8191 15162 8200
rect 15120 8090 15148 8191
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7546 15332 8894
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15396 8537 15424 8570
rect 15382 8528 15438 8537
rect 15382 8463 15438 8472
rect 14738 7511 14794 7520
rect 14832 7540 14884 7546
rect 14752 7274 14780 7511
rect 14832 7482 14884 7488
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15304 7342 15332 7482
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 15396 6866 15424 8463
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 7002 15516 7822
rect 15764 7546 15792 11104
rect 15948 10452 15976 11154
rect 16028 10464 16080 10470
rect 15948 10424 16028 10452
rect 16028 10406 16080 10412
rect 16040 10130 16068 10406
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 16132 9058 16160 12650
rect 16224 12209 16252 12718
rect 16210 12200 16266 12209
rect 16210 12135 16266 12144
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16224 11762 16252 12038
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16224 9654 16252 11698
rect 16408 10810 16436 12838
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16500 11336 16528 12786
rect 16592 11506 16620 17002
rect 16960 16794 16988 17138
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17052 16114 17080 16594
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16776 15162 16804 15506
rect 16868 15337 16896 15846
rect 17052 15706 17080 16050
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16854 15328 16910 15337
rect 16854 15263 16910 15272
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16868 13394 16896 13942
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16868 12986 16896 13330
rect 17144 12986 17172 20703
rect 17328 20505 17356 21286
rect 17420 21078 17448 21490
rect 17684 21344 17736 21350
rect 17684 21286 17736 21292
rect 17408 21072 17460 21078
rect 17408 21014 17460 21020
rect 17696 20602 17724 21286
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17314 20496 17370 20505
rect 17314 20431 17370 20440
rect 17696 20330 17724 20538
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17696 20058 17724 20266
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17696 19514 17724 19994
rect 17684 19508 17736 19514
rect 17684 19450 17736 19456
rect 17684 15904 17736 15910
rect 17682 15872 17684 15881
rect 17736 15872 17738 15881
rect 17682 15807 17738 15816
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17604 14618 17632 15098
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11762 16712 12038
rect 16868 11762 16896 12242
rect 16960 12102 16988 12718
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16856 11756 16908 11762
rect 16908 11716 16988 11744
rect 16856 11698 16908 11704
rect 16592 11478 16712 11506
rect 16580 11348 16632 11354
rect 16500 11308 16580 11336
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16500 10554 16528 11308
rect 16580 11290 16632 11296
rect 16408 10526 16528 10554
rect 16408 10198 16436 10526
rect 16580 10464 16632 10470
rect 16500 10424 16580 10452
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16408 9722 16436 10134
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16500 9178 16528 10424
rect 16684 10441 16712 11478
rect 16580 10406 16632 10412
rect 16670 10432 16726 10441
rect 16670 10367 16726 10376
rect 16960 9722 16988 11716
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16776 9568 16804 9658
rect 16856 9580 16908 9586
rect 16776 9540 16856 9568
rect 16856 9522 16908 9528
rect 16868 9178 16896 9522
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 15936 9036 15988 9042
rect 16132 9030 16252 9058
rect 15936 8978 15988 8984
rect 15948 8566 15976 8978
rect 16028 8968 16080 8974
rect 16120 8968 16172 8974
rect 16028 8910 16080 8916
rect 16118 8936 16120 8945
rect 16172 8936 16174 8945
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15934 8120 15990 8129
rect 15934 8055 15990 8064
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15948 6934 15976 8055
rect 16040 7546 16068 8910
rect 16118 8871 16174 8880
rect 16132 8634 16160 8871
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16224 7857 16252 9030
rect 16580 8832 16632 8838
rect 16408 8780 16580 8786
rect 16408 8774 16632 8780
rect 16408 8758 16620 8774
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16316 8294 16344 8434
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16210 7848 16266 7857
rect 16210 7783 16266 7792
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16316 7410 16344 8230
rect 16408 7834 16436 8758
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16488 8016 16540 8022
rect 16592 8004 16620 8298
rect 16776 8265 16804 8366
rect 16762 8256 16818 8265
rect 16540 7976 16620 8004
rect 16684 8214 16762 8242
rect 16488 7958 16540 7964
rect 16488 7880 16540 7886
rect 16408 7828 16488 7834
rect 16408 7822 16540 7828
rect 16408 7806 16528 7822
rect 16500 7478 16528 7806
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15396 6458 15424 6802
rect 15948 6458 15976 6870
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16408 6458 16436 6802
rect 16684 6662 16712 8214
rect 16762 8191 16818 8200
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16776 7342 16804 8026
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 6730 16896 7142
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 16960 4593 16988 9318
rect 16946 4584 17002 4593
rect 16946 4519 17002 4528
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 17052 3097 17080 9454
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17144 8974 17172 9318
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8634 17172 8910
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17144 4049 17172 6054
rect 17420 5001 17448 11494
rect 17498 10568 17554 10577
rect 17498 10503 17554 10512
rect 17512 7886 17540 10503
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17696 7954 17724 9862
rect 17788 9722 17816 23276
rect 17972 23254 18000 23310
rect 18340 23254 18368 24754
rect 17960 23248 18012 23254
rect 17958 23216 17960 23225
rect 18328 23248 18380 23254
rect 18012 23216 18014 23225
rect 18328 23190 18380 23196
rect 17958 23151 18014 23160
rect 18510 22944 18566 22953
rect 18510 22879 18566 22888
rect 18524 22778 18552 22879
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 18708 22545 18736 25350
rect 18878 25256 18934 25265
rect 18878 25191 18934 25200
rect 18892 24954 18920 25191
rect 18880 24948 18932 24954
rect 18880 24890 18932 24896
rect 18892 24750 18920 24890
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18800 23730 18828 24074
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18800 23322 18828 23666
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 18694 22536 18750 22545
rect 18694 22471 18750 22480
rect 18328 22432 18380 22438
rect 18328 22374 18380 22380
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17880 21690 17908 22034
rect 18340 22030 18368 22374
rect 18696 22228 18748 22234
rect 18696 22170 18748 22176
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17880 21146 17908 21626
rect 18340 21350 18368 21966
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18616 21418 18644 21830
rect 18604 21412 18656 21418
rect 18604 21354 18656 21360
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 18616 21078 18644 21354
rect 18604 21072 18656 21078
rect 18604 21014 18656 21020
rect 17866 20632 17922 20641
rect 17866 20567 17868 20576
rect 17920 20567 17922 20576
rect 17868 20538 17920 20544
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 18064 19922 18092 20334
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18616 19174 18644 19858
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18616 18766 18644 19110
rect 18708 18902 18736 22170
rect 18984 20602 19012 22986
rect 19076 21146 19104 25706
rect 19536 25226 19564 27520
rect 19984 26172 20036 26178
rect 19984 26114 20036 26120
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19996 25362 20024 26114
rect 20088 25498 20116 27520
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 19524 25220 19576 25226
rect 19524 25162 19576 25168
rect 19246 24848 19302 24857
rect 19246 24783 19302 24792
rect 19260 24614 19288 24783
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 19352 23526 19380 24142
rect 19536 23866 19564 24550
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20180 24342 20208 24550
rect 20548 24410 20576 24550
rect 20536 24404 20588 24410
rect 20536 24346 20588 24352
rect 20168 24336 20220 24342
rect 20168 24278 20220 24284
rect 20352 24268 20404 24274
rect 20352 24210 20404 24216
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19890 23896 19946 23905
rect 19524 23860 19576 23866
rect 19890 23831 19892 23840
rect 19524 23802 19576 23808
rect 19944 23831 19946 23840
rect 19892 23802 19944 23808
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19260 21593 19288 22918
rect 19352 22409 19380 23462
rect 19444 23050 19472 23598
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19338 22400 19394 22409
rect 19338 22335 19394 22344
rect 19444 22273 19472 22714
rect 19536 22438 19564 23122
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19720 22817 19748 23054
rect 19706 22808 19762 22817
rect 19706 22743 19762 22752
rect 19904 22545 19932 23054
rect 19890 22536 19946 22545
rect 19996 22506 20024 24142
rect 20364 23798 20392 24210
rect 20352 23792 20404 23798
rect 20350 23760 20352 23769
rect 20404 23760 20406 23769
rect 20350 23695 20406 23704
rect 20640 22953 20668 27520
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20812 24676 20864 24682
rect 20812 24618 20864 24624
rect 20720 22976 20772 22982
rect 20626 22944 20682 22953
rect 20720 22918 20772 22924
rect 20626 22879 20682 22888
rect 19890 22471 19946 22480
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 20352 22500 20404 22506
rect 20352 22442 20404 22448
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19430 22264 19486 22273
rect 19622 22256 19918 22276
rect 19430 22199 19486 22208
rect 20364 22098 20392 22442
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 19706 21992 19762 22001
rect 19706 21927 19708 21936
rect 19760 21927 19762 21936
rect 19708 21898 19760 21904
rect 19246 21584 19302 21593
rect 19246 21519 19302 21528
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19062 20632 19118 20641
rect 18972 20596 19024 20602
rect 19062 20567 19118 20576
rect 18972 20538 19024 20544
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18064 18426 18092 18702
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 17880 16998 17908 17750
rect 18524 17377 18552 18022
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18510 17368 18566 17377
rect 18510 17303 18566 17312
rect 18708 17202 18736 17478
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18694 17096 18750 17105
rect 18694 17031 18750 17040
rect 18708 16998 18736 17031
rect 17868 16992 17920 16998
rect 18696 16992 18748 16998
rect 17868 16934 17920 16940
rect 18510 16960 18566 16969
rect 17880 16794 17908 16934
rect 18696 16934 18748 16940
rect 18510 16895 18566 16904
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 18050 16688 18106 16697
rect 18050 16623 18106 16632
rect 18064 16250 18092 16623
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18432 16114 18460 16390
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18142 15736 18198 15745
rect 18432 15706 18460 16050
rect 18524 15706 18552 16895
rect 18708 16833 18736 16934
rect 18694 16824 18750 16833
rect 18694 16759 18696 16768
rect 18748 16759 18750 16768
rect 18696 16730 18748 16736
rect 18696 16040 18748 16046
rect 18616 15988 18696 15994
rect 18616 15982 18748 15988
rect 18616 15966 18736 15982
rect 18616 15910 18644 15966
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18142 15671 18198 15680
rect 18420 15700 18472 15706
rect 18050 14920 18106 14929
rect 18050 14855 18106 14864
rect 18064 14822 18092 14855
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18050 13152 18106 13161
rect 18050 13087 18106 13096
rect 18064 12986 18092 13087
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18156 12646 18184 15671
rect 18420 15642 18472 15648
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18248 14618 18276 14894
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18340 13870 18368 14758
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18340 13530 18368 13806
rect 18432 13802 18460 14350
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18340 12918 18368 13466
rect 18616 13433 18644 15846
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18708 14618 18736 14826
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18708 13802 18736 14214
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18602 13424 18658 13433
rect 18602 13359 18658 13368
rect 18604 13184 18656 13190
rect 18708 13172 18736 13738
rect 18656 13144 18736 13172
rect 18604 13126 18656 13132
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18156 12102 18184 12582
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 17880 11778 17908 12038
rect 18156 11937 18184 12038
rect 18142 11928 18198 11937
rect 18142 11863 18198 11872
rect 17880 11750 18000 11778
rect 17972 10810 18000 11750
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18064 11354 18092 11494
rect 18156 11393 18184 11494
rect 18142 11384 18198 11393
rect 18052 11348 18104 11354
rect 18142 11319 18144 11328
rect 18052 11290 18104 11296
rect 18196 11319 18198 11328
rect 18144 11290 18196 11296
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 18064 10742 18092 11154
rect 18248 11121 18276 12718
rect 18340 12238 18368 12854
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18340 11626 18368 12174
rect 18432 11762 18460 12786
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18616 12209 18644 12242
rect 18602 12200 18658 12209
rect 18602 12135 18658 12144
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18340 11150 18368 11562
rect 18616 11354 18644 12135
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18328 11144 18380 11150
rect 18234 11112 18290 11121
rect 18328 11086 18380 11092
rect 18234 11047 18290 11056
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 18340 9926 18368 11086
rect 18708 10577 18736 13144
rect 18694 10568 18750 10577
rect 18694 10503 18750 10512
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18616 9994 18644 10406
rect 18800 10305 18828 20198
rect 19076 18970 19104 20567
rect 19168 20482 19196 21354
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19248 20596 19300 20602
rect 19352 20584 19380 20946
rect 20364 20942 20392 21286
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 19628 20641 19656 20878
rect 19300 20556 19380 20584
rect 19614 20632 19670 20641
rect 19614 20567 19670 20576
rect 19248 20538 19300 20544
rect 19168 20466 19380 20482
rect 19168 20460 19392 20466
rect 19168 20454 19340 20460
rect 19340 20402 19392 20408
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 19352 20058 19380 20402
rect 20364 20330 20392 20402
rect 20352 20324 20404 20330
rect 20352 20266 20404 20272
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 20088 20097 20116 20198
rect 20074 20088 20130 20097
rect 19340 20052 19392 20058
rect 20074 20023 20130 20032
rect 19340 19994 19392 20000
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19076 18086 19104 18770
rect 19064 18080 19116 18086
rect 19062 18048 19064 18057
rect 19116 18048 19118 18057
rect 19062 17983 19118 17992
rect 19168 17882 19196 18838
rect 19352 18698 19380 19994
rect 20364 19514 20392 20266
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19352 18426 19380 18634
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19156 17876 19208 17882
rect 19156 17818 19208 17824
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18892 16697 18920 16730
rect 18878 16688 18934 16697
rect 18878 16623 18934 16632
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 18786 10296 18842 10305
rect 18786 10231 18842 10240
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17788 8498 17816 8978
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17696 7410 17724 7890
rect 17788 7818 17816 8434
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17880 7546 17908 8298
rect 18248 7857 18276 9590
rect 18340 9518 18368 9862
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 18524 8945 18552 9386
rect 18892 8945 18920 15914
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18984 14958 19012 15302
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 19076 14890 19104 15098
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 19076 14634 19104 14826
rect 18953 14606 19104 14634
rect 18953 14532 18981 14606
rect 18953 14504 19012 14532
rect 18984 12628 19012 14504
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 19076 13326 19104 14418
rect 19064 13320 19116 13326
rect 19062 13288 19064 13297
rect 19116 13288 19118 13297
rect 19062 13223 19118 13232
rect 19168 12782 19196 17818
rect 19260 17542 19288 18158
rect 19536 18086 19564 18566
rect 19982 18320 20038 18329
rect 19982 18255 20038 18264
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19338 17776 19394 17785
rect 19338 17711 19394 17720
rect 19432 17740 19484 17746
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 19246 16960 19302 16969
rect 19246 16895 19302 16904
rect 19260 16794 19288 16895
rect 19352 16794 19380 17711
rect 19432 17682 19484 17688
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19352 16250 19380 16730
rect 19444 16658 19472 17682
rect 19536 16998 19564 18022
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17882 20024 18255
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19338 16008 19394 16017
rect 19338 15943 19394 15952
rect 19352 15706 19380 15943
rect 19444 15858 19472 16594
rect 19536 16590 19564 16934
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20456 16658 20484 22374
rect 20732 22234 20760 22918
rect 20824 22778 20852 24618
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20812 22160 20864 22166
rect 20812 22102 20864 22108
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 20732 20942 20760 21286
rect 20720 20936 20772 20942
rect 20640 20896 20720 20924
rect 20640 18630 20668 20896
rect 20720 20878 20772 20884
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20732 16794 20760 20742
rect 20824 20398 20852 22102
rect 20916 21622 20944 25842
rect 21284 24857 21312 27520
rect 21836 25498 21864 27520
rect 21824 25492 21876 25498
rect 21824 25434 21876 25440
rect 21270 24848 21326 24857
rect 20996 24812 21048 24818
rect 21270 24783 21326 24792
rect 21548 24812 21600 24818
rect 20996 24754 21048 24760
rect 21548 24754 21600 24760
rect 21008 23662 21036 24754
rect 21560 24313 21588 24754
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21546 24304 21602 24313
rect 21546 24239 21602 24248
rect 21824 24268 21876 24274
rect 21824 24210 21876 24216
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 21270 23624 21326 23633
rect 21008 23322 21036 23598
rect 21270 23559 21326 23568
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 21008 22778 21036 23258
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 21284 21350 21312 23559
rect 21744 23526 21772 24142
rect 21836 24138 21864 24210
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21732 23520 21784 23526
rect 21732 23462 21784 23468
rect 21468 23118 21496 23462
rect 21744 23186 21772 23462
rect 21928 23361 21956 24550
rect 22008 24064 22060 24070
rect 22008 24006 22060 24012
rect 21914 23352 21970 23361
rect 21914 23287 21970 23296
rect 21732 23180 21784 23186
rect 21732 23122 21784 23128
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21468 22574 21496 23054
rect 21546 22808 21602 22817
rect 21546 22743 21602 22752
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21560 21894 21588 22743
rect 21744 22030 21772 23122
rect 21824 22704 21876 22710
rect 21822 22672 21824 22681
rect 21876 22672 21878 22681
rect 22020 22658 22048 24006
rect 22388 23905 22416 27520
rect 22652 25832 22704 25838
rect 22652 25774 22704 25780
rect 22664 25498 22692 25774
rect 22652 25492 22704 25498
rect 22652 25434 22704 25440
rect 22928 25152 22980 25158
rect 22928 25094 22980 25100
rect 22742 24848 22798 24857
rect 22940 24818 22968 25094
rect 22742 24783 22798 24792
rect 22928 24812 22980 24818
rect 22652 24676 22704 24682
rect 22652 24618 22704 24624
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22480 24313 22508 24550
rect 22466 24304 22522 24313
rect 22466 24239 22522 24248
rect 22374 23896 22430 23905
rect 22374 23831 22430 23840
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22100 22704 22152 22710
rect 22020 22652 22100 22658
rect 22020 22646 22152 22652
rect 22020 22630 22140 22646
rect 21822 22607 21878 22616
rect 22098 22536 22154 22545
rect 22098 22471 22154 22480
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21744 21894 21772 21966
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21560 21486 21588 21830
rect 21548 21480 21600 21486
rect 21548 21422 21600 21428
rect 21272 21344 21324 21350
rect 21732 21344 21784 21350
rect 21272 21286 21324 21292
rect 21362 21312 21418 21321
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20824 20058 20852 20198
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20824 19689 20852 19994
rect 20916 19718 20944 20198
rect 21192 19718 21220 20946
rect 21284 19961 21312 21286
rect 21732 21286 21784 21292
rect 21362 21247 21418 21256
rect 21376 20942 21404 21247
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21376 20058 21404 20878
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21270 19952 21326 19961
rect 21270 19887 21326 19896
rect 21548 19916 21600 19922
rect 21548 19858 21600 19864
rect 20904 19712 20956 19718
rect 20810 19680 20866 19689
rect 20904 19654 20956 19660
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 20810 19615 20866 19624
rect 20916 18873 20944 19654
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 21008 19174 21036 19314
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20902 18864 20958 18873
rect 20902 18799 20958 18808
rect 20810 18456 20866 18465
rect 20810 18391 20866 18400
rect 20824 18193 20852 18391
rect 20810 18184 20866 18193
rect 20810 18119 20866 18128
rect 21086 18184 21142 18193
rect 21086 18119 21142 18128
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20824 17270 20852 17614
rect 20902 17504 20958 17513
rect 20902 17439 20958 17448
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20720 16788 20772 16794
rect 20640 16748 20720 16776
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19536 15978 19564 16526
rect 19996 16250 20024 16526
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 19444 15830 19564 15858
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19260 14414 19288 15370
rect 19352 15162 19380 15642
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19248 14408 19300 14414
rect 19246 14376 19248 14385
rect 19300 14376 19302 14385
rect 19246 14311 19302 14320
rect 19260 14074 19288 14311
rect 19444 14249 19472 15438
rect 19536 14550 19564 15830
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19996 14890 20024 15302
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19708 14272 19760 14278
rect 19430 14240 19486 14249
rect 19430 14175 19486 14184
rect 19706 14240 19708 14249
rect 19760 14240 19762 14249
rect 19706 14175 19762 14184
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19996 14006 20024 14826
rect 19984 14000 20036 14006
rect 19338 13968 19394 13977
rect 19984 13942 20036 13948
rect 19338 13903 19394 13912
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 18984 12600 19196 12628
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18984 10130 19012 10406
rect 18972 10124 19024 10130
rect 18972 10066 19024 10072
rect 18510 8936 18566 8945
rect 18510 8871 18512 8880
rect 18564 8871 18566 8880
rect 18878 8936 18934 8945
rect 18878 8871 18934 8880
rect 18512 8842 18564 8848
rect 18984 8634 19012 10066
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18234 7848 18290 7857
rect 18234 7783 18290 7792
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17512 6458 17540 6938
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17604 6633 17632 6870
rect 17696 6798 17724 7346
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 18248 6662 18276 7142
rect 18236 6656 18288 6662
rect 17590 6624 17646 6633
rect 18236 6598 18288 6604
rect 17590 6559 17646 6568
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17604 6118 17632 6559
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 18248 5137 18276 6598
rect 18234 5128 18290 5137
rect 18234 5063 18290 5072
rect 17406 4992 17462 5001
rect 17406 4927 17462 4936
rect 17130 4040 17186 4049
rect 17130 3975 17186 3984
rect 18524 3641 18552 7210
rect 18800 5273 18828 8298
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19076 7546 19104 7822
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19168 6905 19196 12600
rect 19260 10810 19288 13126
rect 19352 12782 19380 13903
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19812 12986 19840 13262
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19444 12102 19472 12922
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19444 11218 19472 12038
rect 19536 11694 19564 12650
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19524 11688 19576 11694
rect 19996 11665 20024 13942
rect 20180 12102 20208 16594
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 15910 20484 16390
rect 20640 16046 20668 16748
rect 20720 16730 20772 16736
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20364 12889 20392 13126
rect 20456 12986 20484 15846
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20548 12918 20576 15914
rect 20732 14618 20760 16594
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20536 12912 20588 12918
rect 20350 12880 20406 12889
rect 20536 12854 20588 12860
rect 20350 12815 20406 12824
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20456 12306 20484 12650
rect 20548 12442 20576 12854
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20640 12220 20668 13330
rect 20720 12232 20772 12238
rect 20640 12192 20720 12220
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20444 12096 20496 12102
rect 20640 12073 20668 12192
rect 20720 12174 20772 12180
rect 20444 12038 20496 12044
rect 20626 12064 20682 12073
rect 20074 11928 20130 11937
rect 20074 11863 20130 11872
rect 19524 11630 19576 11636
rect 19982 11656 20038 11665
rect 19982 11591 20038 11600
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19352 10674 19380 11018
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19444 10062 19472 11154
rect 19984 10736 20036 10742
rect 19982 10704 19984 10713
rect 20036 10704 20038 10713
rect 19982 10639 20038 10648
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19248 10056 19300 10062
rect 19432 10056 19484 10062
rect 19300 10016 19380 10044
rect 19248 9998 19300 10004
rect 19352 8634 19380 10016
rect 19432 9998 19484 10004
rect 19444 9654 19472 9998
rect 19982 9888 20038 9897
rect 19982 9823 20038 9832
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19536 9178 19564 9318
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19536 8498 19564 9114
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19628 8430 19656 8910
rect 19904 8566 19932 8910
rect 19892 8560 19944 8566
rect 19890 8528 19892 8537
rect 19944 8528 19946 8537
rect 19890 8463 19946 8472
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19340 8016 19392 8022
rect 19338 7984 19340 7993
rect 19392 7984 19394 7993
rect 19260 7942 19338 7970
rect 19154 6896 19210 6905
rect 19260 6866 19288 7942
rect 19338 7919 19394 7928
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19628 7410 19656 7822
rect 19996 7546 20024 9823
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 20088 7410 20116 11863
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20180 11082 20208 11562
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20272 9926 20300 10542
rect 20350 10296 20406 10305
rect 20350 10231 20406 10240
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20272 9625 20300 9862
rect 20258 9616 20314 9625
rect 20258 9551 20314 9560
rect 20364 7410 20392 10231
rect 20456 9654 20484 12038
rect 20626 11999 20682 12008
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20732 10810 20760 11630
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20732 10062 20760 10746
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20088 6866 20116 7346
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 19154 6831 19210 6840
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 18786 5264 18842 5273
rect 18786 5199 18842 5208
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 20180 3913 20208 7210
rect 20364 7002 20392 7346
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 20456 4729 20484 9590
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 9178 20576 9318
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20640 8090 20668 8434
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20824 7993 20852 16730
rect 20916 15609 20944 17439
rect 20902 15600 20958 15609
rect 21100 15570 21128 18119
rect 20902 15535 20958 15544
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 21100 15162 21128 15506
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20916 14414 20944 14758
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20916 13938 20944 14350
rect 20994 13968 21050 13977
rect 20904 13932 20956 13938
rect 20994 13903 21050 13912
rect 20904 13874 20956 13880
rect 20916 13394 20944 13874
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20916 12986 20944 13330
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20916 9178 20944 9386
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20902 8664 20958 8673
rect 20902 8599 20958 8608
rect 20916 8498 20944 8599
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 20902 8392 20958 8401
rect 20902 8327 20904 8336
rect 20956 8327 20958 8336
rect 20904 8298 20956 8304
rect 20810 7984 20866 7993
rect 21008 7954 21036 13903
rect 21100 13530 21128 14486
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21086 12200 21142 12209
rect 21086 12135 21142 12144
rect 21100 9382 21128 12135
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21100 8498 21128 9318
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 20810 7919 20866 7928
rect 20996 7948 21048 7954
rect 20996 7890 21048 7896
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20640 7546 20668 7822
rect 21008 7546 21036 7890
rect 21086 7848 21142 7857
rect 21086 7783 21088 7792
rect 21140 7783 21142 7792
rect 21088 7754 21140 7760
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 21192 7410 21220 19654
rect 21468 19417 21496 19654
rect 21454 19408 21510 19417
rect 21454 19343 21510 19352
rect 21560 18630 21588 19858
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21468 17746 21496 18022
rect 21456 17740 21508 17746
rect 21456 17682 21508 17688
rect 21468 16998 21496 17682
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21270 16688 21326 16697
rect 21270 16623 21326 16632
rect 21284 15978 21312 16623
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21376 16250 21404 16526
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21468 16114 21496 16934
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21272 15972 21324 15978
rect 21272 15914 21324 15920
rect 21284 15706 21312 15914
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21270 15056 21326 15065
rect 21270 14991 21326 15000
rect 21284 14958 21312 14991
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21284 14074 21312 14894
rect 21376 14822 21404 15438
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21270 13424 21326 13433
rect 21270 13359 21326 13368
rect 21284 11354 21312 13359
rect 21560 12714 21588 18566
rect 21638 17232 21694 17241
rect 21638 17167 21694 17176
rect 21652 17066 21680 17167
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21652 16794 21680 17002
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 21744 16046 21772 21286
rect 21836 20806 21864 22374
rect 21914 21992 21970 22001
rect 21914 21927 21970 21936
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21822 20224 21878 20233
rect 21822 20159 21878 20168
rect 21836 18970 21864 20159
rect 21928 20058 21956 21927
rect 22112 20890 22140 22471
rect 22204 21978 22232 22714
rect 22468 22704 22520 22710
rect 22468 22646 22520 22652
rect 22480 22574 22508 22646
rect 22572 22642 22600 22918
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22468 22568 22520 22574
rect 22468 22510 22520 22516
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 22388 22234 22416 22374
rect 22480 22234 22508 22510
rect 22376 22228 22428 22234
rect 22376 22170 22428 22176
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 22664 22080 22692 24618
rect 22480 22052 22692 22080
rect 22204 21950 22324 21978
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22204 21078 22232 21830
rect 22296 21690 22324 21950
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22376 21616 22428 21622
rect 22376 21558 22428 21564
rect 22192 21072 22244 21078
rect 22192 21014 22244 21020
rect 22112 20862 22232 20890
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 22008 19236 22060 19242
rect 22008 19178 22060 19184
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21836 18086 21864 18770
rect 22020 18170 22048 19178
rect 22112 18465 22140 20742
rect 22204 20602 22232 20862
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22296 19242 22324 19790
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22296 18766 22324 18906
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22098 18456 22154 18465
rect 22098 18391 22154 18400
rect 21928 18142 22140 18170
rect 22296 18154 22324 18702
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21744 15706 21772 15982
rect 21732 15700 21784 15706
rect 21732 15642 21784 15648
rect 21836 15586 21864 18022
rect 21928 16590 21956 18142
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 22020 17116 22048 18022
rect 22112 17882 22140 18142
rect 22284 18148 22336 18154
rect 22284 18090 22336 18096
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22100 17128 22152 17134
rect 22020 17088 22100 17116
rect 22100 17070 22152 17076
rect 22112 16794 22140 17070
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 21916 16584 21968 16590
rect 21916 16526 21968 16532
rect 21928 16182 21956 16526
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 21916 16176 21968 16182
rect 21916 16118 21968 16124
rect 22020 16130 22048 16186
rect 22020 16102 22140 16130
rect 21744 15558 21864 15586
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21640 12368 21692 12374
rect 21640 12310 21692 12316
rect 21744 12322 21772 15558
rect 22112 15162 22140 16102
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22006 15056 22062 15065
rect 22006 14991 22062 15000
rect 21914 13832 21970 13841
rect 21914 13767 21970 13776
rect 21928 12986 21956 13767
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21652 11898 21680 12310
rect 21744 12294 21864 12322
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21362 10704 21418 10713
rect 21362 10639 21418 10648
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 21284 8809 21312 8978
rect 21270 8800 21326 8809
rect 21270 8735 21326 8744
rect 21284 8634 21312 8735
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21284 8537 21312 8570
rect 21270 8528 21326 8537
rect 21270 8463 21326 8472
rect 21376 8430 21404 10639
rect 21468 10538 21496 11494
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 21468 8974 21496 10474
rect 21640 9376 21692 9382
rect 21744 9353 21772 11018
rect 21836 10713 21864 12294
rect 22020 12170 22048 14991
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 21822 10704 21878 10713
rect 21822 10639 21878 10648
rect 21928 10062 21956 10950
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21928 9722 21956 9998
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 22008 9512 22060 9518
rect 22006 9480 22008 9489
rect 22060 9480 22062 9489
rect 22006 9415 22062 9424
rect 21640 9318 21692 9324
rect 21730 9344 21786 9353
rect 21652 9178 21680 9318
rect 21730 9279 21786 9288
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21546 8936 21602 8945
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 21468 8090 21496 8910
rect 21546 8871 21602 8880
rect 21560 8673 21588 8871
rect 21546 8664 21602 8673
rect 21546 8599 21602 8608
rect 22112 8498 22140 13670
rect 22204 12782 22232 17478
rect 22296 14482 22324 18090
rect 22388 17338 22416 21558
rect 22480 18222 22508 22052
rect 22558 21992 22614 22001
rect 22558 21927 22560 21936
rect 22612 21927 22614 21936
rect 22560 21898 22612 21904
rect 22756 21146 22784 24783
rect 22928 24754 22980 24760
rect 22940 24614 22968 24754
rect 23032 24721 23060 27520
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23018 24712 23074 24721
rect 23018 24647 23074 24656
rect 23202 24712 23258 24721
rect 23202 24647 23204 24656
rect 23256 24647 23258 24656
rect 23204 24618 23256 24624
rect 22928 24608 22980 24614
rect 22928 24550 22980 24556
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22848 23526 22876 24210
rect 22940 24206 22968 24550
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22836 23520 22888 23526
rect 22836 23462 22888 23468
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22742 21040 22798 21049
rect 22560 21004 22612 21010
rect 22742 20975 22798 20984
rect 22560 20946 22612 20952
rect 22572 20602 22600 20946
rect 22560 20596 22612 20602
rect 22560 20538 22612 20544
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22480 17882 22508 18158
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22374 16416 22430 16425
rect 22374 16351 22430 16360
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22282 14376 22338 14385
rect 22282 14311 22284 14320
rect 22336 14311 22338 14320
rect 22284 14282 22336 14288
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22204 11558 22232 12174
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 22204 10130 22232 10406
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22204 9586 22232 10066
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22204 9110 22232 9522
rect 22192 9104 22244 9110
rect 22192 9046 22244 9052
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 22296 6633 22324 11630
rect 22388 7410 22416 16351
rect 22480 15706 22508 17138
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22480 13394 22508 13670
rect 22572 13569 22600 20538
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22664 18902 22692 19858
rect 22652 18896 22704 18902
rect 22652 18838 22704 18844
rect 22650 17912 22706 17921
rect 22650 17847 22706 17856
rect 22664 15162 22692 17847
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22650 14920 22706 14929
rect 22650 14855 22706 14864
rect 22558 13560 22614 13569
rect 22558 13495 22614 13504
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22480 12832 22508 13330
rect 22572 13025 22600 13495
rect 22558 13016 22614 13025
rect 22558 12951 22614 12960
rect 22560 12844 22612 12850
rect 22480 12804 22560 12832
rect 22560 12786 22612 12792
rect 22468 12708 22520 12714
rect 22468 12650 22520 12656
rect 22480 12220 22508 12650
rect 22572 12374 22600 12786
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22480 12192 22600 12220
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 11014 22508 11494
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22466 9616 22522 9625
rect 22466 9551 22522 9560
rect 22480 9178 22508 9551
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22572 8090 22600 12192
rect 22664 9081 22692 14855
rect 22756 9761 22784 20975
rect 22848 18970 22876 23462
rect 22940 22438 22968 24142
rect 23020 22976 23072 22982
rect 23020 22918 23072 22924
rect 22928 22432 22980 22438
rect 22928 22374 22980 22380
rect 22928 22092 22980 22098
rect 22928 22034 22980 22040
rect 22940 21962 22968 22034
rect 22928 21956 22980 21962
rect 22928 21898 22980 21904
rect 22940 21078 22968 21898
rect 22928 21072 22980 21078
rect 22928 21014 22980 21020
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 22836 18624 22888 18630
rect 22836 18566 22888 18572
rect 22848 18290 22876 18566
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22848 18193 22876 18226
rect 22834 18184 22890 18193
rect 22834 18119 22890 18128
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22940 16998 22968 17614
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22940 16794 22968 16934
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 22940 14006 22968 15642
rect 22928 14000 22980 14006
rect 22834 13968 22890 13977
rect 22928 13942 22980 13948
rect 22834 13903 22836 13912
rect 22888 13903 22890 13912
rect 22836 13874 22888 13880
rect 22834 13696 22890 13705
rect 22834 13631 22890 13640
rect 22848 11898 22876 13631
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22940 11801 22968 12582
rect 23032 11898 23060 22918
rect 23124 17542 23152 24346
rect 23388 24132 23440 24138
rect 23388 24074 23440 24080
rect 23296 24064 23348 24070
rect 23296 24006 23348 24012
rect 23202 23080 23258 23089
rect 23202 23015 23258 23024
rect 23216 21894 23244 23015
rect 23308 22692 23336 24006
rect 23400 23322 23428 24074
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23492 22817 23520 24754
rect 23584 24177 23612 27520
rect 23754 27160 23810 27169
rect 23754 27095 23810 27104
rect 23768 25498 23796 27095
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 23768 24750 23796 25434
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23756 24744 23808 24750
rect 23676 24692 23756 24698
rect 23676 24686 23808 24692
rect 23676 24670 23796 24686
rect 23860 24682 23888 25298
rect 23848 24676 23900 24682
rect 23570 24168 23626 24177
rect 23570 24103 23626 24112
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23478 22808 23534 22817
rect 23478 22743 23534 22752
rect 23308 22664 23520 22692
rect 23492 22574 23520 22664
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23308 22166 23336 22374
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 23308 19174 23336 22102
rect 23492 22001 23520 22374
rect 23478 21992 23534 22001
rect 23478 21927 23534 21936
rect 23584 21622 23612 23462
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23480 21344 23532 21350
rect 23400 21304 23480 21332
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 23296 18080 23348 18086
rect 23400 18068 23428 21304
rect 23480 21286 23532 21292
rect 23584 20482 23612 21422
rect 23676 20913 23704 24670
rect 23848 24618 23900 24624
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23768 22506 23796 24550
rect 23756 22500 23808 22506
rect 23756 22442 23808 22448
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23662 20904 23718 20913
rect 23662 20839 23718 20848
rect 23492 20454 23612 20482
rect 23492 18426 23520 20454
rect 23676 20346 23704 20839
rect 23768 20806 23796 21966
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23584 20318 23704 20346
rect 23584 18714 23612 20318
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23676 18816 23704 20198
rect 23768 19854 23796 20742
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23768 19242 23796 19654
rect 23860 19281 23888 24618
rect 23952 24410 23980 27639
rect 24122 27520 24178 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25870 27520 25926 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 24136 24857 24164 27520
rect 24214 26616 24270 26625
rect 24214 26551 24270 26560
rect 24122 24848 24178 24857
rect 24122 24783 24178 24792
rect 24124 24744 24176 24750
rect 24228 24698 24256 26551
rect 24780 25226 24808 27520
rect 25226 26072 25282 26081
rect 25226 26007 25282 26016
rect 25136 25356 25188 25362
rect 25136 25298 25188 25304
rect 24768 25220 24820 25226
rect 24768 25162 24820 25168
rect 24676 25152 24728 25158
rect 24676 25094 24728 25100
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24176 24692 24256 24698
rect 24124 24686 24256 24692
rect 24136 24670 24256 24686
rect 24228 24614 24256 24670
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 23940 24404 23992 24410
rect 23940 24346 23992 24352
rect 24216 24200 24268 24206
rect 24320 24188 24348 24754
rect 24268 24160 24348 24188
rect 24216 24142 24268 24148
rect 24228 23730 24256 24142
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24582 23760 24638 23769
rect 24216 23724 24268 23730
rect 24582 23695 24638 23704
rect 24216 23666 24268 23672
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 23952 22030 23980 23462
rect 24136 22982 24164 23462
rect 24398 23352 24454 23361
rect 24398 23287 24454 23296
rect 24412 23254 24440 23287
rect 24400 23248 24452 23254
rect 24400 23190 24452 23196
rect 24216 23112 24268 23118
rect 24216 23054 24268 23060
rect 24596 23066 24624 23695
rect 24688 23225 24716 25094
rect 25148 24886 25176 25298
rect 25136 24880 25188 24886
rect 25136 24822 25188 24828
rect 25240 24410 25268 26007
rect 25332 25430 25360 27520
rect 25884 25498 25912 27520
rect 25872 25492 25924 25498
rect 25872 25434 25924 25440
rect 25320 25424 25372 25430
rect 25320 25366 25372 25372
rect 25502 25392 25558 25401
rect 25502 25327 25558 25336
rect 25410 24848 25466 24857
rect 25410 24783 25466 24792
rect 25424 24614 25452 24783
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25516 24410 25544 25327
rect 25780 24744 25832 24750
rect 25780 24686 25832 24692
rect 25228 24404 25280 24410
rect 25228 24346 25280 24352
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24872 23338 24900 24006
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 24964 23633 24992 23734
rect 24950 23624 25006 23633
rect 24950 23559 25006 23568
rect 24780 23322 24900 23338
rect 25240 23322 25268 24346
rect 25410 24032 25466 24041
rect 25410 23967 25466 23976
rect 25424 23866 25452 23967
rect 25412 23860 25464 23866
rect 25412 23802 25464 23808
rect 25516 23798 25544 24346
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 25700 23866 25728 24142
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25504 23792 25556 23798
rect 25504 23734 25556 23740
rect 25688 23656 25740 23662
rect 25688 23598 25740 23604
rect 24768 23316 24900 23322
rect 24820 23310 24900 23316
rect 24768 23258 24820 23264
rect 24674 23216 24730 23225
rect 24674 23151 24730 23160
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 23952 21146 23980 21966
rect 24044 21690 24072 21966
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 24044 21298 24072 21490
rect 24136 21418 24164 22714
rect 24228 22642 24256 23054
rect 24596 23038 24716 23066
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22778 24716 23038
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 24228 22030 24256 22578
rect 24872 22098 24900 23310
rect 24952 23316 25004 23322
rect 24952 23258 25004 23264
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24124 21412 24176 21418
rect 24124 21354 24176 21360
rect 24044 21270 24164 21298
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 23952 20330 23980 20946
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 24044 20398 24072 20742
rect 24032 20392 24084 20398
rect 24136 20369 24164 21270
rect 24228 20942 24256 21830
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24964 21706 24992 23258
rect 25044 23248 25096 23254
rect 25044 23190 25096 23196
rect 25056 22778 25084 23190
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 25148 22574 25176 22918
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 25320 22568 25372 22574
rect 25320 22510 25372 22516
rect 25594 22536 25650 22545
rect 25332 22114 25360 22510
rect 25594 22471 25650 22480
rect 25148 22098 25360 22114
rect 25044 22092 25096 22098
rect 25044 22034 25096 22040
rect 25148 22092 25372 22098
rect 25148 22086 25320 22092
rect 24780 21678 24992 21706
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24504 20942 24532 21490
rect 24780 21486 24808 21678
rect 24860 21616 24912 21622
rect 24860 21558 24912 21564
rect 24768 21480 24820 21486
rect 24768 21422 24820 21428
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24216 20936 24268 20942
rect 24216 20878 24268 20884
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24032 20334 24084 20340
rect 24122 20360 24178 20369
rect 23940 20324 23992 20330
rect 24122 20295 24178 20304
rect 23940 20266 23992 20272
rect 23846 19272 23902 19281
rect 23756 19236 23808 19242
rect 23846 19207 23902 19216
rect 23756 19178 23808 19184
rect 23952 19009 23980 20266
rect 24124 20256 24176 20262
rect 24122 20224 24124 20233
rect 24176 20224 24178 20233
rect 24122 20159 24178 20168
rect 24136 20058 24164 20159
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24228 19922 24256 20878
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20505 24716 20946
rect 24766 20904 24822 20913
rect 24766 20839 24822 20848
rect 24674 20496 24730 20505
rect 24674 20431 24676 20440
rect 24728 20431 24730 20440
rect 24676 20402 24728 20408
rect 24216 19916 24268 19922
rect 24216 19858 24268 19864
rect 24124 19848 24176 19854
rect 24124 19790 24176 19796
rect 24032 19168 24084 19174
rect 24032 19110 24084 19116
rect 23938 19000 23994 19009
rect 23938 18935 23994 18944
rect 23938 18864 23994 18873
rect 23756 18828 23808 18834
rect 23676 18788 23756 18816
rect 24044 18850 24072 19110
rect 23994 18822 24072 18850
rect 23938 18799 23994 18808
rect 23756 18770 23808 18776
rect 23768 18737 23796 18770
rect 23952 18766 23980 18799
rect 23940 18760 23992 18766
rect 23754 18728 23810 18737
rect 23584 18686 23704 18714
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23348 18040 23428 18068
rect 23296 18022 23348 18028
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 23124 16658 23152 17206
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 23124 16250 23152 16594
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 23124 14074 23152 14214
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23124 13870 23152 14010
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 23216 12866 23244 17274
rect 23294 16960 23350 16969
rect 23294 16895 23350 16904
rect 23308 16726 23336 16895
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23308 16182 23336 16662
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23400 15450 23428 17478
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23492 15706 23520 15914
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23308 15422 23428 15450
rect 23308 13462 23336 15422
rect 23386 15328 23442 15337
rect 23386 15263 23442 15272
rect 23400 15178 23428 15263
rect 23400 15162 23520 15178
rect 23400 15156 23532 15162
rect 23400 15150 23480 15156
rect 23480 15098 23532 15104
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23492 14074 23520 14350
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23400 13530 23428 13874
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23296 13456 23348 13462
rect 23296 13398 23348 13404
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23400 12986 23428 13126
rect 23478 13016 23534 13025
rect 23388 12980 23440 12986
rect 23478 12951 23534 12960
rect 23388 12922 23440 12928
rect 23492 12918 23520 12951
rect 23480 12912 23532 12918
rect 23112 12844 23164 12850
rect 23216 12838 23428 12866
rect 23480 12854 23532 12860
rect 23112 12786 23164 12792
rect 23124 12306 23152 12786
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 22926 11792 22982 11801
rect 22926 11727 22982 11736
rect 23032 11694 23060 11834
rect 23020 11688 23072 11694
rect 23020 11630 23072 11636
rect 23124 11354 23152 12242
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 23020 11008 23072 11014
rect 22834 10976 22890 10985
rect 23020 10950 23072 10956
rect 22834 10911 22890 10920
rect 22742 9752 22798 9761
rect 22742 9687 22798 9696
rect 22650 9072 22706 9081
rect 22650 9007 22706 9016
rect 22848 8945 22876 10911
rect 23032 10810 23060 10950
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 23308 10266 23336 11222
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23032 9722 23060 10202
rect 23112 9988 23164 9994
rect 23112 9930 23164 9936
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23124 9178 23152 9930
rect 23400 9908 23428 12838
rect 23492 12782 23520 12854
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23584 11778 23612 18566
rect 23676 18222 23704 18686
rect 23940 18702 23992 18708
rect 23754 18663 23810 18672
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23676 17814 23704 18022
rect 23664 17808 23716 17814
rect 23664 17750 23716 17756
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 23846 17368 23902 17377
rect 23846 17303 23902 17312
rect 23754 16960 23810 16969
rect 23754 16895 23810 16904
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23676 13734 23704 14486
rect 23768 14362 23796 16895
rect 23860 15706 23888 17303
rect 24044 17066 24072 17614
rect 24032 17060 24084 17066
rect 24032 17002 24084 17008
rect 24044 15910 24072 17002
rect 24136 16425 24164 19790
rect 24674 19680 24730 19689
rect 24289 19612 24585 19632
rect 24674 19615 24730 19624
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24492 19236 24544 19242
rect 24492 19178 24544 19184
rect 24504 18902 24532 19178
rect 24492 18896 24544 18902
rect 24492 18838 24544 18844
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24228 17542 24256 18226
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24122 16416 24178 16425
rect 24122 16351 24178 16360
rect 24228 15978 24256 17478
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24398 17096 24454 17105
rect 24398 17031 24454 17040
rect 24412 16794 24440 17031
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24216 15972 24268 15978
rect 24216 15914 24268 15920
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 24122 15736 24178 15745
rect 23848 15700 23900 15706
rect 23900 15660 23980 15688
rect 24122 15671 24178 15680
rect 23848 15642 23900 15648
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23860 15162 23888 15506
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23860 14482 23888 15098
rect 23952 14958 23980 15660
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 23938 14512 23994 14521
rect 23848 14476 23900 14482
rect 23938 14447 23994 14456
rect 23848 14418 23900 14424
rect 23768 14334 23888 14362
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 13938 23796 14214
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23676 12458 23704 13670
rect 23754 13560 23810 13569
rect 23754 13495 23756 13504
rect 23808 13495 23810 13504
rect 23756 13466 23808 13472
rect 23768 12646 23796 13466
rect 23860 13326 23888 14334
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23676 12430 23796 12458
rect 23662 12064 23718 12073
rect 23662 11999 23718 12008
rect 23676 11898 23704 11999
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23584 11750 23704 11778
rect 23570 11656 23626 11665
rect 23570 11591 23626 11600
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23492 11121 23520 11494
rect 23478 11112 23534 11121
rect 23478 11047 23534 11056
rect 23584 10810 23612 11591
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23216 9880 23428 9908
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 22928 9104 22980 9110
rect 22928 9046 22980 9052
rect 22834 8936 22890 8945
rect 22834 8871 22890 8880
rect 22940 8634 22968 9046
rect 23124 8634 23152 9114
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 23216 7954 23244 9880
rect 23676 9722 23704 11750
rect 23768 10656 23796 12430
rect 23860 10810 23888 13126
rect 23952 12714 23980 14447
rect 24044 13530 24072 15302
rect 24136 13705 24164 15671
rect 24228 15094 24256 15914
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15162 24716 19615
rect 24780 18442 24808 20839
rect 24872 20058 24900 21558
rect 25056 21350 25084 22034
rect 25044 21344 25096 21350
rect 25042 21312 25044 21321
rect 25096 21312 25098 21321
rect 25042 21247 25098 21256
rect 25148 21162 25176 22086
rect 25320 22034 25372 22040
rect 25410 21992 25466 22001
rect 25410 21927 25466 21936
rect 25228 21888 25280 21894
rect 25228 21830 25280 21836
rect 24964 21134 25176 21162
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 24860 19712 24912 19718
rect 24860 19654 24912 19660
rect 24872 18970 24900 19654
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24780 18426 24900 18442
rect 24780 18420 24912 18426
rect 24780 18414 24860 18420
rect 24860 18362 24912 18368
rect 24766 17504 24822 17513
rect 24766 17439 24822 17448
rect 24780 15688 24808 17439
rect 24780 15660 24900 15688
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24216 15088 24268 15094
rect 24216 15030 24268 15036
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24214 14648 24270 14657
rect 24214 14583 24270 14592
rect 24122 13696 24178 13705
rect 24122 13631 24178 13640
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 24044 12918 24072 13466
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 24136 12986 24164 13262
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 24228 12866 24256 14583
rect 24412 14414 24440 14962
rect 24780 14618 24808 15506
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24308 14408 24360 14414
rect 24306 14376 24308 14385
rect 24400 14408 24452 14414
rect 24360 14376 24362 14385
rect 24400 14350 24452 14356
rect 24306 14311 24362 14320
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24766 13968 24822 13977
rect 24766 13903 24822 13912
rect 24308 13864 24360 13870
rect 24306 13832 24308 13841
rect 24360 13832 24362 13841
rect 24306 13767 24362 13776
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24400 12912 24452 12918
rect 24228 12850 24348 12866
rect 24400 12854 24452 12860
rect 24228 12844 24360 12850
rect 24228 12838 24308 12844
rect 24308 12786 24360 12792
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 24308 12708 24360 12714
rect 24308 12650 24360 12656
rect 24320 12322 24348 12650
rect 24412 12442 24440 12854
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24596 12374 24624 12582
rect 24228 12294 24348 12322
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24228 12186 24256 12294
rect 24136 12158 24256 12186
rect 24306 12200 24362 12209
rect 24030 11928 24086 11937
rect 24030 11863 24086 11872
rect 24044 11694 24072 11863
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 24136 11642 24164 12158
rect 24306 12135 24308 12144
rect 24360 12135 24362 12144
rect 24308 12106 24360 12112
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 24228 11762 24256 12038
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24044 11354 24072 11630
rect 24136 11614 24348 11642
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 24320 11121 24348 11614
rect 24306 11112 24362 11121
rect 24306 11047 24362 11056
rect 24124 11008 24176 11014
rect 24124 10950 24176 10956
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 23768 10628 23980 10656
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 9926 23888 10406
rect 23848 9920 23900 9926
rect 23846 9888 23848 9897
rect 23900 9888 23902 9897
rect 23846 9823 23902 9832
rect 23952 9738 23980 10628
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23860 9710 23980 9738
rect 23308 8974 23336 9658
rect 23754 9616 23810 9625
rect 23754 9551 23810 9560
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23308 8566 23336 8910
rect 23478 8800 23534 8809
rect 23478 8735 23534 8744
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23216 7546 23244 7890
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22282 6624 22338 6633
rect 22282 6559 22338 6568
rect 20442 4720 20498 4729
rect 20442 4655 20498 4664
rect 23492 4185 23520 8735
rect 23570 8528 23626 8537
rect 23570 8463 23626 8472
rect 23584 5273 23612 8463
rect 23676 7954 23704 9454
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23676 7546 23704 7890
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23662 7440 23718 7449
rect 23768 7410 23796 9551
rect 23860 9217 23888 9710
rect 23940 9512 23992 9518
rect 23940 9454 23992 9460
rect 23846 9208 23902 9217
rect 23846 9143 23902 9152
rect 23860 9042 23888 9143
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23846 8392 23902 8401
rect 23846 8327 23902 8336
rect 23662 7375 23718 7384
rect 23756 7404 23808 7410
rect 23676 7342 23704 7375
rect 23756 7346 23808 7352
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 23754 7304 23810 7313
rect 23754 7239 23810 7248
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23676 6769 23704 6802
rect 23662 6760 23718 6769
rect 23662 6695 23718 6704
rect 23676 6458 23704 6695
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23570 5264 23626 5273
rect 23570 5199 23626 5208
rect 23570 4584 23626 4593
rect 23570 4519 23626 4528
rect 23478 4176 23534 4185
rect 23478 4111 23534 4120
rect 20166 3904 20222 3913
rect 19622 3836 19918 3856
rect 20166 3839 20222 3848
rect 23478 3904 23534 3913
rect 23478 3839 23534 3848
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 22190 3768 22246 3777
rect 22190 3703 22246 3712
rect 18510 3632 18566 3641
rect 18510 3567 18566 3576
rect 22006 3632 22062 3641
rect 22204 3618 22232 3703
rect 22062 3590 22232 3618
rect 22006 3567 22062 3576
rect 23202 3496 23258 3505
rect 23202 3431 23258 3440
rect 17038 3088 17094 3097
rect 17038 3023 17094 3032
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14646 1592 14702 1601
rect 14646 1527 14702 1536
rect 23216 480 23244 3431
rect 23492 921 23520 3839
rect 23584 2553 23612 4519
rect 23570 2544 23626 2553
rect 23570 2479 23626 2488
rect 23768 2009 23796 7239
rect 23860 7177 23888 8327
rect 23952 8090 23980 9454
rect 24044 8634 24072 10746
rect 24136 10606 24164 10950
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24136 10266 24164 10542
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24136 9722 24164 10066
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24122 8664 24178 8673
rect 24032 8628 24084 8634
rect 24122 8599 24178 8608
rect 24032 8570 24084 8576
rect 24044 8430 24072 8570
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 24044 7478 24072 8230
rect 24136 7857 24164 8599
rect 24122 7848 24178 7857
rect 24122 7783 24178 7792
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 23846 7168 23902 7177
rect 23846 7103 23902 7112
rect 24122 2136 24178 2145
rect 24228 2122 24256 10406
rect 24582 10296 24638 10305
rect 24582 10231 24584 10240
rect 24636 10231 24638 10240
rect 24584 10202 24636 10208
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9654 24716 12786
rect 24676 9648 24728 9654
rect 24676 9590 24728 9596
rect 24674 9208 24730 9217
rect 24780 9178 24808 13903
rect 24872 11898 24900 15660
rect 24964 15473 24992 21134
rect 25240 20777 25268 21830
rect 25320 21480 25372 21486
rect 25318 21448 25320 21457
rect 25372 21448 25374 21457
rect 25318 21383 25374 21392
rect 25226 20768 25282 20777
rect 25226 20703 25282 20712
rect 25424 20602 25452 21927
rect 25608 21690 25636 22471
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25502 21448 25558 21457
rect 25502 21383 25558 21392
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25226 20088 25282 20097
rect 25226 20023 25282 20032
rect 25412 20052 25464 20058
rect 25044 19168 25096 19174
rect 25044 19110 25096 19116
rect 25056 18358 25084 19110
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 25240 18222 25268 20023
rect 25412 19994 25464 20000
rect 25320 19848 25372 19854
rect 25318 19816 25320 19825
rect 25372 19816 25374 19825
rect 25318 19751 25374 19760
rect 25332 19514 25360 19751
rect 25320 19508 25372 19514
rect 25320 19450 25372 19456
rect 25424 18834 25452 19994
rect 25516 18970 25544 21383
rect 25596 20256 25648 20262
rect 25596 20198 25648 20204
rect 25608 19854 25636 20198
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25608 19446 25636 19790
rect 25596 19440 25648 19446
rect 25596 19382 25648 19388
rect 25504 18964 25556 18970
rect 25504 18906 25556 18912
rect 25608 18902 25636 19382
rect 25596 18896 25648 18902
rect 25596 18838 25648 18844
rect 25412 18828 25464 18834
rect 25412 18770 25464 18776
rect 25596 18760 25648 18766
rect 25596 18702 25648 18708
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25608 17542 25636 18702
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25044 16992 25096 16998
rect 25042 16960 25044 16969
rect 25096 16960 25098 16969
rect 25042 16895 25098 16904
rect 25148 16833 25176 17478
rect 25134 16824 25190 16833
rect 25134 16759 25190 16768
rect 25502 16280 25558 16289
rect 25502 16215 25558 16224
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25240 15502 25268 15846
rect 25228 15496 25280 15502
rect 24950 15464 25006 15473
rect 25228 15438 25280 15444
rect 24950 15399 25006 15408
rect 25240 15094 25268 15438
rect 25228 15088 25280 15094
rect 25228 15030 25280 15036
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 25148 13938 25176 14418
rect 25136 13932 25188 13938
rect 25136 13874 25188 13880
rect 25044 13456 25096 13462
rect 25044 13398 25096 13404
rect 25056 12986 25084 13398
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 24950 12880 25006 12889
rect 24950 12815 25006 12824
rect 24964 12442 24992 12815
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 24952 12436 25004 12442
rect 24952 12378 25004 12384
rect 25056 12322 25084 12718
rect 24964 12294 25084 12322
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24964 11354 24992 12294
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 25056 11830 25084 12174
rect 25044 11824 25096 11830
rect 25044 11766 25096 11772
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24950 11248 25006 11257
rect 24950 11183 24952 11192
rect 25004 11183 25006 11192
rect 24952 11154 25004 11160
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24872 10470 24900 11086
rect 24964 10810 24992 11154
rect 25044 11008 25096 11014
rect 25148 10985 25176 13874
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 25044 10950 25096 10956
rect 25134 10976 25190 10985
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 25056 10266 25084 10950
rect 25134 10911 25190 10920
rect 25240 10826 25268 13806
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25320 13388 25372 13394
rect 25320 13330 25372 13336
rect 25332 12918 25360 13330
rect 25320 12912 25372 12918
rect 25424 12889 25452 13670
rect 25320 12854 25372 12860
rect 25410 12880 25466 12889
rect 25332 12753 25360 12854
rect 25410 12815 25466 12824
rect 25318 12744 25374 12753
rect 25318 12679 25374 12688
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25424 12345 25452 12582
rect 25410 12336 25466 12345
rect 25410 12271 25466 12280
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 25318 10976 25374 10985
rect 25318 10911 25374 10920
rect 25148 10798 25268 10826
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 24872 9654 24900 10134
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24964 9450 24992 9862
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 24858 9344 24914 9353
rect 24858 9279 24914 9288
rect 24674 9143 24730 9152
rect 24768 9172 24820 9178
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24178 2094 24256 2122
rect 24122 2071 24178 2080
rect 23754 2000 23810 2009
rect 23754 1935 23810 1944
rect 23478 912 23534 921
rect 23478 847 23534 856
rect 3238 368 3294 377
rect 3238 303 3294 312
rect 4618 0 4674 480
rect 13910 0 13966 480
rect 23202 0 23258 480
rect 24688 377 24716 9143
rect 24768 9114 24820 9120
rect 24766 9072 24822 9081
rect 24766 9007 24822 9016
rect 24780 8430 24808 9007
rect 24872 8634 24900 9279
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 25056 8634 25084 8978
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 25148 8090 25176 10798
rect 25332 10742 25360 10911
rect 25320 10736 25372 10742
rect 25226 10704 25282 10713
rect 25320 10678 25372 10684
rect 25226 10639 25282 10648
rect 25240 10606 25268 10639
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25424 8566 25452 11290
rect 25516 10810 25544 16215
rect 25608 13410 25636 17478
rect 25700 14618 25728 23598
rect 25688 14612 25740 14618
rect 25688 14554 25740 14560
rect 25792 13530 25820 24686
rect 26528 24426 26556 27520
rect 27080 24857 27108 27520
rect 27066 24848 27122 24857
rect 27066 24783 27122 24792
rect 26160 24398 26556 24426
rect 26160 22778 26188 24398
rect 27632 24041 27660 27520
rect 27618 24032 27674 24041
rect 27618 23967 27674 23976
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 26238 18728 26294 18737
rect 26238 18663 26294 18672
rect 26252 18426 26280 18663
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 25872 17740 25924 17746
rect 25872 17682 25924 17688
rect 25884 16998 25912 17682
rect 25872 16992 25924 16998
rect 25872 16934 25924 16940
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 25608 13382 25820 13410
rect 25594 13288 25650 13297
rect 25594 13223 25650 13232
rect 25608 12442 25636 13223
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25608 11354 25636 12378
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25700 9926 25728 11630
rect 25688 9920 25740 9926
rect 25688 9862 25740 9868
rect 25412 8560 25464 8566
rect 25412 8502 25464 8508
rect 25792 8294 25820 13382
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 24766 7984 24822 7993
rect 24766 7919 24768 7928
rect 24820 7919 24822 7928
rect 24768 7890 24820 7896
rect 24780 7546 24808 7890
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 25884 6730 25912 16934
rect 26148 12164 26200 12170
rect 26148 12106 26200 12112
rect 26160 11898 26188 12106
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 25872 6724 25924 6730
rect 25872 6666 25924 6672
rect 24674 368 24730 377
rect 24674 303 24730 312
<< via2 >>
rect 4434 27648 4490 27704
rect 1214 26560 1270 26616
rect 1306 24792 1362 24848
rect 1674 25336 1730 25392
rect 2502 25200 2558 25256
rect 2318 24792 2374 24848
rect 2042 23704 2098 23760
rect 3054 26016 3110 26072
rect 1766 22380 1768 22400
rect 1768 22380 1820 22400
rect 1820 22380 1822 22400
rect 1766 22344 1822 22380
rect 1582 21120 1638 21176
rect 1398 20032 1454 20088
rect 294 15408 350 15464
rect 1490 17720 1546 17776
rect 1950 22616 2006 22672
rect 1582 17448 1638 17504
rect 1858 19760 1914 19816
rect 2042 18944 2098 19000
rect 1950 17856 2006 17912
rect 2962 24928 3018 24984
rect 2410 23024 2466 23080
rect 2870 23432 2926 23488
rect 2410 21256 2466 21312
rect 2318 20168 2374 20224
rect 1582 15680 1638 15736
rect 1582 14592 1638 14648
rect 1490 13912 1546 13968
rect 1582 13368 1638 13424
rect 1582 12824 1638 12880
rect 2226 16224 2282 16280
rect 2962 23296 3018 23352
rect 2410 16496 2466 16552
rect 3054 23160 3110 23216
rect 2962 21392 3018 21448
rect 2962 19488 3018 19544
rect 2962 18844 2964 18864
rect 2964 18844 3016 18864
rect 3016 18844 3018 18864
rect 2962 18808 3018 18844
rect 2778 18128 2834 18184
rect 3330 24520 3386 24576
rect 3238 23180 3294 23216
rect 3238 23160 3240 23180
rect 3240 23160 3292 23180
rect 3292 23160 3294 23180
rect 3606 24112 3662 24168
rect 3790 24248 3846 24304
rect 3330 21004 3386 21040
rect 3330 20984 3332 21004
rect 3332 20984 3384 21004
rect 3384 20984 3386 21004
rect 3238 20712 3294 20768
rect 3330 20460 3386 20496
rect 3330 20440 3332 20460
rect 3332 20440 3384 20460
rect 3384 20440 3386 20460
rect 3146 19760 3202 19816
rect 2502 15020 2558 15056
rect 2502 15000 2504 15020
rect 2504 15000 2556 15020
rect 2556 15000 2558 15020
rect 2686 15136 2742 15192
rect 2134 12588 2136 12608
rect 2136 12588 2188 12608
rect 2188 12588 2190 12608
rect 2134 12552 2190 12588
rect 2686 12280 2742 12336
rect 3330 20168 3386 20224
rect 3514 19352 3570 19408
rect 3330 15700 3386 15736
rect 3330 15680 3332 15700
rect 3332 15680 3384 15700
rect 3384 15680 3386 15700
rect 3238 14728 3294 14784
rect 3054 13504 3110 13560
rect 3146 12824 3202 12880
rect 3054 12688 3110 12744
rect 3606 19216 3662 19272
rect 4066 23432 4122 23488
rect 3882 21392 3938 21448
rect 3882 20848 3938 20904
rect 4066 20848 4122 20904
rect 23938 27648 23994 27704
rect 4802 27104 4858 27160
rect 4526 21528 4582 21584
rect 4618 21256 4674 21312
rect 4802 20204 4804 20224
rect 4804 20204 4856 20224
rect 4856 20204 4858 20224
rect 4802 20168 4858 20204
rect 4434 20052 4490 20088
rect 4434 20032 4436 20052
rect 4436 20032 4488 20052
rect 4488 20032 4490 20052
rect 4342 19896 4398 19952
rect 4342 19660 4344 19680
rect 4344 19660 4396 19680
rect 4396 19660 4398 19680
rect 4342 19624 4398 19660
rect 4342 19488 4398 19544
rect 4526 19216 4582 19272
rect 4250 17720 4306 17776
rect 4250 16788 4306 16824
rect 4250 16768 4252 16788
rect 4252 16768 4304 16788
rect 4304 16768 4306 16788
rect 3698 15564 3754 15600
rect 3698 15544 3700 15564
rect 3700 15544 3752 15564
rect 3752 15544 3754 15564
rect 3882 15408 3938 15464
rect 4066 14592 4122 14648
rect 3330 13504 3386 13560
rect 3238 11736 3294 11792
rect 2962 9288 3018 9344
rect 1858 9016 1914 9072
rect 2962 7112 3018 7168
rect 3146 3576 3202 3632
rect 3698 13640 3754 13696
rect 4066 11736 4122 11792
rect 3882 10376 3938 10432
rect 3698 9424 3754 9480
rect 3514 9152 3570 9208
rect 4434 11328 4490 11384
rect 5906 25220 5962 25256
rect 5906 25200 5908 25220
rect 5908 25200 5960 25220
rect 5960 25200 5962 25220
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 6090 24928 6146 24984
rect 5998 24656 6054 24712
rect 5354 24112 5410 24168
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5998 23296 6054 23352
rect 5998 23024 6054 23080
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 6090 22752 6146 22808
rect 5538 22380 5540 22400
rect 5540 22380 5592 22400
rect 5592 22380 5594 22400
rect 5538 22344 5594 22380
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5354 20712 5410 20768
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 6642 23704 6698 23760
rect 6458 21800 6514 21856
rect 6366 21140 6422 21176
rect 6366 21120 6368 21140
rect 6368 21120 6420 21140
rect 6420 21120 6422 21140
rect 6366 20032 6422 20088
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5446 18400 5502 18456
rect 4894 17720 4950 17776
rect 5814 18028 5816 18048
rect 5816 18028 5868 18048
rect 5868 18028 5870 18048
rect 5814 17992 5870 18028
rect 5538 17876 5594 17912
rect 5538 17856 5540 17876
rect 5540 17856 5592 17876
rect 5592 17856 5594 17876
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5538 17196 5594 17232
rect 5538 17176 5540 17196
rect 5540 17176 5592 17196
rect 5592 17176 5594 17196
rect 5354 17040 5410 17096
rect 5446 16088 5502 16144
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 4986 15816 5042 15872
rect 5354 15272 5410 15328
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5538 14356 5540 14376
rect 5540 14356 5592 14376
rect 5592 14356 5594 14376
rect 5538 14320 5594 14356
rect 6182 17720 6238 17776
rect 6182 15408 6238 15464
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5354 13912 5410 13968
rect 6274 14612 6330 14648
rect 6274 14592 6276 14612
rect 6276 14592 6328 14612
rect 6328 14592 6330 14612
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5630 12824 5686 12880
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6826 24792 6882 24848
rect 7286 24792 7342 24848
rect 6826 23704 6882 23760
rect 6734 22888 6790 22944
rect 6918 23180 6974 23216
rect 6918 23160 6920 23180
rect 6920 23160 6972 23180
rect 6972 23160 6974 23180
rect 7010 21936 7066 21992
rect 7286 24248 7342 24304
rect 7470 22772 7526 22808
rect 7470 22752 7472 22772
rect 7472 22752 7524 22772
rect 7524 22752 7526 22772
rect 6918 21392 6974 21448
rect 6918 21120 6974 21176
rect 7194 21392 7250 21448
rect 7010 20848 7066 20904
rect 6734 20712 6790 20768
rect 6826 20596 6882 20632
rect 6826 20576 6828 20596
rect 6828 20576 6880 20596
rect 6880 20576 6882 20596
rect 7194 20848 7250 20904
rect 7102 19080 7158 19136
rect 6550 18128 6606 18184
rect 7286 18808 7342 18864
rect 7194 16632 7250 16688
rect 7378 17448 7434 17504
rect 7378 16904 7434 16960
rect 7010 15408 7066 15464
rect 6734 14864 6790 14920
rect 7010 12688 7066 12744
rect 7930 24132 7986 24168
rect 7930 24112 7932 24132
rect 7932 24112 7984 24132
rect 7984 24112 7986 24132
rect 7838 23432 7894 23488
rect 7838 22752 7894 22808
rect 8114 24656 8170 24712
rect 8114 23568 8170 23624
rect 7562 17040 7618 17096
rect 7470 15408 7526 15464
rect 7470 15272 7526 15328
rect 7286 12708 7342 12744
rect 7286 12688 7288 12708
rect 7288 12688 7340 12708
rect 7340 12688 7342 12708
rect 7378 12316 7380 12336
rect 7380 12316 7432 12336
rect 7432 12316 7434 12336
rect 7378 12280 7434 12316
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 4526 10240 4582 10296
rect 4066 9968 4122 10024
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 6550 8200 6606 8256
rect 6550 7656 6606 7712
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 7838 18944 7894 19000
rect 7838 18708 7840 18728
rect 7840 18708 7892 18728
rect 7892 18708 7894 18728
rect 7838 18672 7894 18708
rect 7838 18300 7840 18320
rect 7840 18300 7892 18320
rect 7892 18300 7894 18320
rect 7838 18264 7894 18300
rect 8022 19624 8078 19680
rect 8022 17312 8078 17368
rect 7838 16940 7840 16960
rect 7840 16940 7892 16960
rect 7892 16940 7894 16960
rect 7838 16904 7894 16940
rect 7838 15680 7894 15736
rect 7838 14340 7894 14376
rect 7838 14320 7840 14340
rect 7840 14320 7892 14340
rect 7892 14320 7894 14340
rect 7838 13640 7894 13696
rect 8022 16632 8078 16688
rect 8022 15544 8078 15600
rect 8298 22344 8354 22400
rect 8298 21548 8354 21584
rect 8298 21528 8300 21548
rect 8300 21528 8352 21548
rect 8352 21528 8354 21548
rect 8390 20748 8392 20768
rect 8392 20748 8444 20768
rect 8444 20748 8446 20768
rect 8390 20712 8446 20748
rect 8666 23468 8668 23488
rect 8668 23468 8720 23488
rect 8720 23468 8722 23488
rect 8666 23432 8722 23468
rect 8758 23060 8760 23080
rect 8760 23060 8812 23080
rect 8812 23060 8814 23080
rect 8758 23024 8814 23060
rect 8574 21292 8576 21312
rect 8576 21292 8628 21312
rect 8628 21292 8630 21312
rect 8574 21256 8630 21292
rect 8298 19352 8354 19408
rect 8206 18164 8208 18184
rect 8208 18164 8260 18184
rect 8260 18164 8262 18184
rect 8206 18128 8262 18164
rect 8390 17584 8446 17640
rect 8390 17040 8446 17096
rect 8298 16088 8354 16144
rect 8482 16088 8538 16144
rect 8114 14048 8170 14104
rect 8574 15952 8630 16008
rect 9402 23704 9458 23760
rect 8850 20052 8906 20088
rect 8850 20032 8852 20052
rect 8852 20032 8904 20052
rect 8904 20032 8906 20052
rect 8850 16360 8906 16416
rect 8482 13524 8538 13560
rect 8482 13504 8484 13524
rect 8484 13504 8536 13524
rect 8536 13504 8538 13524
rect 8390 12824 8446 12880
rect 8390 11328 8446 11384
rect 8850 13096 8906 13152
rect 9034 20440 9090 20496
rect 9034 18400 9090 18456
rect 9034 17740 9090 17776
rect 9034 17720 9036 17740
rect 9036 17720 9088 17740
rect 9088 17720 9090 17740
rect 9586 19352 9642 19408
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10414 25220 10470 25256
rect 10414 25200 10416 25220
rect 10416 25200 10468 25220
rect 10468 25200 10470 25220
rect 10690 24656 10746 24712
rect 10138 24520 10194 24576
rect 10046 24384 10102 24440
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10138 23840 10194 23896
rect 11150 24792 11206 24848
rect 10966 24284 10968 24304
rect 10968 24284 11020 24304
rect 11020 24284 11022 24304
rect 10966 24248 11022 24284
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 11058 23468 11060 23488
rect 11060 23468 11112 23488
rect 11112 23468 11114 23488
rect 11058 23432 11114 23468
rect 10138 23160 10194 23216
rect 9954 22888 10010 22944
rect 9862 22072 9918 22128
rect 9310 18536 9366 18592
rect 9402 17856 9458 17912
rect 9494 17720 9550 17776
rect 9402 17212 9404 17232
rect 9404 17212 9456 17232
rect 9456 17212 9458 17232
rect 9402 17176 9458 17212
rect 9126 13368 9182 13424
rect 9034 12588 9036 12608
rect 9036 12588 9088 12608
rect 9088 12588 9090 12608
rect 9034 12552 9090 12588
rect 9310 13776 9366 13832
rect 9678 17604 9734 17640
rect 9678 17584 9680 17604
rect 9680 17584 9732 17604
rect 9732 17584 9734 17604
rect 9678 16904 9734 16960
rect 9678 16088 9734 16144
rect 10138 22888 10194 22944
rect 10966 22888 11022 22944
rect 11334 22616 11390 22672
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10690 22208 10746 22264
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10046 20204 10048 20224
rect 10048 20204 10100 20224
rect 10100 20204 10102 20224
rect 10046 20168 10102 20204
rect 10046 19660 10048 19680
rect 10048 19660 10100 19680
rect 10100 19660 10102 19680
rect 10046 19624 10102 19660
rect 9402 12688 9458 12744
rect 9402 11600 9458 11656
rect 9218 11192 9274 11248
rect 8850 11056 8906 11112
rect 8758 10648 8814 10704
rect 8666 9424 8722 9480
rect 9678 9424 9734 9480
rect 8022 8880 8078 8936
rect 10230 20576 10286 20632
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10230 19488 10286 19544
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10138 18672 10194 18728
rect 10506 18708 10508 18728
rect 10508 18708 10560 18728
rect 10560 18708 10562 18728
rect 10506 18672 10562 18708
rect 10322 18536 10378 18592
rect 10230 18264 10286 18320
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10322 15444 10324 15464
rect 10324 15444 10376 15464
rect 10376 15444 10378 15464
rect 10322 15408 10378 15444
rect 10138 14764 10140 14784
rect 10140 14764 10192 14784
rect 10192 14764 10194 14784
rect 10138 14728 10194 14764
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10046 10512 10102 10568
rect 10966 21664 11022 21720
rect 10966 21528 11022 21584
rect 10874 21004 10930 21040
rect 10874 20984 10876 21004
rect 10876 20984 10928 21004
rect 10928 20984 10930 21004
rect 11794 24792 11850 24848
rect 11794 23704 11850 23760
rect 11518 21800 11574 21856
rect 11150 20440 11206 20496
rect 11058 20304 11114 20360
rect 10874 20032 10930 20088
rect 10966 19760 11022 19816
rect 10874 19488 10930 19544
rect 10782 16940 10784 16960
rect 10784 16940 10836 16960
rect 10836 16940 10838 16960
rect 10782 16904 10838 16940
rect 11150 19624 11206 19680
rect 11058 19216 11114 19272
rect 11058 17312 11114 17368
rect 10874 16224 10930 16280
rect 11978 25780 11980 25800
rect 11980 25780 12032 25800
rect 12032 25780 12034 25800
rect 11978 25744 12034 25780
rect 12162 25336 12218 25392
rect 12070 23860 12126 23896
rect 12070 23840 12072 23860
rect 12072 23840 12124 23860
rect 12124 23840 12126 23860
rect 11518 21256 11574 21312
rect 11518 21140 11574 21176
rect 11518 21120 11520 21140
rect 11520 21120 11572 21140
rect 11572 21120 11574 21140
rect 11334 17312 11390 17368
rect 11426 16788 11482 16824
rect 11426 16768 11428 16788
rect 11428 16768 11480 16788
rect 11480 16768 11482 16788
rect 11150 16224 11206 16280
rect 10782 15156 10838 15192
rect 10782 15136 10784 15156
rect 10784 15136 10836 15156
rect 10836 15136 10838 15156
rect 11150 15272 11206 15328
rect 11150 14184 11206 14240
rect 10782 12280 10838 12336
rect 10874 11076 10930 11112
rect 10874 11056 10876 11076
rect 10876 11056 10928 11076
rect 10928 11056 10930 11076
rect 10138 10376 10194 10432
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10046 10240 10102 10296
rect 11794 21528 11850 21584
rect 12070 21256 12126 21312
rect 11886 20440 11942 20496
rect 11610 17856 11666 17912
rect 11334 15952 11390 16008
rect 9862 9324 9864 9344
rect 9864 9324 9916 9344
rect 9916 9324 9918 9344
rect 9862 9288 9918 9324
rect 9954 9152 10010 9208
rect 9770 7928 9826 7984
rect 7470 7520 7526 7576
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10138 7384 10194 7440
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10782 6840 10838 6896
rect 4066 6704 4122 6760
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 4066 6024 4122 6080
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 4066 5344 4122 5400
rect 3974 5208 4030 5264
rect 3882 4800 3938 4856
rect 10690 4936 10746 4992
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 4066 4664 4122 4720
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 3974 4256 4030 4312
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 11150 11736 11206 11792
rect 11242 11056 11298 11112
rect 11610 15000 11666 15056
rect 11426 12164 11482 12200
rect 11426 12144 11428 12164
rect 11428 12144 11480 12164
rect 11480 12144 11482 12164
rect 12254 23840 12310 23896
rect 12806 25780 12808 25800
rect 12808 25780 12860 25800
rect 12860 25780 12862 25800
rect 12806 25744 12862 25780
rect 12898 24656 12954 24712
rect 12714 24112 12770 24168
rect 12806 23704 12862 23760
rect 12622 22072 12678 22128
rect 12622 21428 12624 21448
rect 12624 21428 12676 21448
rect 12676 21428 12678 21448
rect 12622 21392 12678 21428
rect 12254 18808 12310 18864
rect 12162 18400 12218 18456
rect 12254 17992 12310 18048
rect 12162 13796 12218 13832
rect 12162 13776 12164 13796
rect 12164 13776 12216 13796
rect 12216 13776 12218 13796
rect 11886 12008 11942 12064
rect 11702 11872 11758 11928
rect 12162 11620 12218 11656
rect 12162 11600 12164 11620
rect 12164 11600 12216 11620
rect 12216 11600 12218 11620
rect 12438 17176 12494 17232
rect 12806 20848 12862 20904
rect 12806 18672 12862 18728
rect 12714 18128 12770 18184
rect 12898 18264 12954 18320
rect 12530 16224 12586 16280
rect 13174 17312 13230 17368
rect 13358 24248 13414 24304
rect 13542 23044 13598 23080
rect 13542 23024 13544 23044
rect 13544 23024 13596 23044
rect 13596 23024 13598 23044
rect 13726 23432 13782 23488
rect 13634 22888 13690 22944
rect 13542 22616 13598 22672
rect 13634 22344 13690 22400
rect 13358 19896 13414 19952
rect 13818 19216 13874 19272
rect 13450 18284 13506 18320
rect 13450 18264 13452 18284
rect 13452 18264 13504 18284
rect 13504 18264 13506 18284
rect 13358 17756 13360 17776
rect 13360 17756 13412 17776
rect 13412 17756 13414 17776
rect 13358 17720 13414 17756
rect 13634 16224 13690 16280
rect 12346 14728 12402 14784
rect 13358 15136 13414 15192
rect 13358 14068 13414 14104
rect 13358 14048 13360 14068
rect 13360 14048 13412 14068
rect 13412 14048 13414 14068
rect 12990 13912 13046 13968
rect 13174 13912 13230 13968
rect 13542 13776 13598 13832
rect 12438 12688 12494 12744
rect 13450 13232 13506 13288
rect 13542 12824 13598 12880
rect 12070 11192 12126 11248
rect 10690 3440 10746 3496
rect 11058 3440 11114 3496
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 3146 856 3202 912
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 3514 2624 3570 2680
rect 4618 2352 4674 2408
rect 3514 1536 3570 1592
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 12254 9696 12310 9752
rect 12070 9288 12126 9344
rect 11886 3576 11942 3632
rect 12162 7928 12218 7984
rect 13542 10376 13598 10432
rect 13266 10240 13322 10296
rect 12714 7284 12716 7304
rect 12716 7284 12768 7304
rect 12768 7284 12770 7304
rect 12714 7248 12770 7284
rect 12622 6296 12678 6352
rect 11978 2488 12034 2544
rect 13266 8472 13322 8528
rect 13818 18536 13874 18592
rect 13818 16360 13874 16416
rect 13818 15988 13820 16008
rect 13820 15988 13872 16008
rect 13872 15988 13874 16008
rect 13818 15952 13874 15988
rect 13726 15680 13782 15736
rect 13726 13232 13782 13288
rect 15474 25372 15476 25392
rect 15476 25372 15528 25392
rect 15528 25372 15530 25392
rect 15474 25336 15530 25372
rect 14278 24132 14334 24168
rect 14278 24112 14280 24132
rect 14280 24112 14332 24132
rect 14332 24112 14334 24132
rect 14278 23296 14334 23352
rect 14094 22480 14150 22536
rect 14094 21664 14150 21720
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14738 23860 14794 23896
rect 14738 23840 14740 23860
rect 14740 23840 14792 23860
rect 14792 23840 14794 23860
rect 14554 20984 14610 21040
rect 14186 19352 14242 19408
rect 14094 18672 14150 18728
rect 14462 19216 14518 19272
rect 14186 16360 14242 16416
rect 14094 15428 14150 15464
rect 14094 15408 14096 15428
rect 14096 15408 14148 15428
rect 14148 15408 14150 15428
rect 14002 13368 14058 13424
rect 14186 13368 14242 13424
rect 14002 12824 14058 12880
rect 14186 11328 14242 11384
rect 14370 16652 14426 16688
rect 14370 16632 14372 16652
rect 14372 16632 14424 16652
rect 14424 16632 14426 16652
rect 15290 23024 15346 23080
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15290 22616 15346 22672
rect 14830 22480 14886 22536
rect 14646 16088 14702 16144
rect 14370 15136 14426 15192
rect 13634 10104 13690 10160
rect 13818 8064 13874 8120
rect 14186 9968 14242 10024
rect 14186 7656 14242 7712
rect 14462 14728 14518 14784
rect 14462 14476 14518 14512
rect 14462 14456 14464 14476
rect 14464 14456 14516 14476
rect 14516 14456 14518 14476
rect 14646 14184 14702 14240
rect 14554 11872 14610 11928
rect 14554 9696 14610 9752
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14830 20848 14886 20904
rect 15474 22038 15530 22094
rect 15658 24792 15714 24848
rect 15382 20748 15384 20768
rect 15384 20748 15436 20768
rect 15436 20748 15438 20768
rect 15382 20712 15438 20748
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15842 24384 15898 24440
rect 15750 22616 15806 22672
rect 15750 21936 15806 21992
rect 15750 21392 15806 21448
rect 15474 20032 15530 20088
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 16394 23704 16450 23760
rect 16762 24656 16818 24712
rect 17130 24792 17186 24848
rect 17038 24520 17094 24576
rect 16854 23740 16856 23760
rect 16856 23740 16908 23760
rect 16908 23740 16910 23760
rect 16854 23704 16910 23740
rect 16670 23296 16726 23352
rect 16302 21256 16358 21312
rect 16762 20984 16818 21040
rect 16210 19760 16266 19816
rect 16394 19624 16450 19680
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15382 17604 15438 17640
rect 15382 17584 15384 17604
rect 15384 17584 15436 17604
rect 15436 17584 15438 17604
rect 15290 17040 15346 17096
rect 15106 16652 15162 16688
rect 15106 16632 15108 16652
rect 15108 16632 15160 16652
rect 15160 16632 15162 16652
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14738 10648 14794 10704
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15382 13812 15384 13832
rect 15384 13812 15436 13832
rect 15436 13812 15438 13832
rect 15382 13776 15438 13812
rect 15382 12688 15438 12744
rect 15290 11736 15346 11792
rect 15842 16632 15898 16688
rect 15658 15272 15714 15328
rect 17406 23044 17462 23080
rect 17406 23024 17408 23044
rect 17408 23024 17460 23044
rect 17460 23024 17462 23044
rect 17774 23588 17830 23624
rect 17774 23568 17776 23588
rect 17776 23568 17828 23588
rect 17828 23568 17830 23588
rect 18234 24384 18290 24440
rect 18050 23432 18106 23488
rect 17406 21972 17408 21992
rect 17408 21972 17460 21992
rect 17460 21972 17462 21992
rect 17406 21936 17462 21972
rect 17130 20712 17186 20768
rect 16762 17856 16818 17912
rect 16762 17448 16818 17504
rect 16118 16088 16174 16144
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15290 10532 15346 10568
rect 15290 10512 15292 10532
rect 15292 10512 15344 10532
rect 15344 10512 15346 10532
rect 15382 10412 15384 10432
rect 15384 10412 15436 10432
rect 15436 10412 15438 10432
rect 15382 10376 15438 10412
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15750 11192 15806 11248
rect 16302 13132 16304 13152
rect 16304 13132 16356 13152
rect 16356 13132 16358 13152
rect 16302 13096 16358 13132
rect 15658 9968 15714 10024
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14554 7928 14610 7984
rect 14370 6704 14426 6760
rect 11978 2388 11980 2408
rect 11980 2388 12032 2408
rect 12032 2388 12034 2408
rect 11978 2352 12034 2388
rect 11794 1536 11850 1592
rect 14738 7520 14794 7576
rect 15106 8200 15162 8256
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15382 8472 15438 8528
rect 16210 12144 16266 12200
rect 16854 15272 16910 15328
rect 17314 20440 17370 20496
rect 17682 15852 17684 15872
rect 17684 15852 17736 15872
rect 17736 15852 17738 15872
rect 17682 15816 17738 15852
rect 16670 10376 16726 10432
rect 16118 8916 16120 8936
rect 16120 8916 16172 8936
rect 16172 8916 16174 8936
rect 15934 8064 15990 8120
rect 16118 8880 16174 8916
rect 16210 7792 16266 7848
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 16762 8200 16818 8256
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 16946 4528 17002 4584
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 17498 10512 17554 10568
rect 17958 23196 17960 23216
rect 17960 23196 18012 23216
rect 18012 23196 18014 23216
rect 17958 23160 18014 23196
rect 18510 22888 18566 22944
rect 18878 25200 18934 25256
rect 18694 22480 18750 22536
rect 17866 20596 17922 20632
rect 17866 20576 17868 20596
rect 17868 20576 17920 20596
rect 17920 20576 17922 20596
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19246 24792 19302 24848
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19890 23860 19946 23896
rect 19890 23840 19892 23860
rect 19892 23840 19944 23860
rect 19944 23840 19946 23860
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19338 22344 19394 22400
rect 19706 22752 19762 22808
rect 19890 22480 19946 22536
rect 20350 23740 20352 23760
rect 20352 23740 20404 23760
rect 20404 23740 20406 23760
rect 20350 23704 20406 23740
rect 20626 22888 20682 22944
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19430 22208 19486 22264
rect 19706 21956 19762 21992
rect 19706 21936 19708 21956
rect 19708 21936 19760 21956
rect 19760 21936 19762 21956
rect 19246 21528 19302 21584
rect 19062 20576 19118 20632
rect 18510 17312 18566 17368
rect 18694 17040 18750 17096
rect 18510 16904 18566 16960
rect 18050 16632 18106 16688
rect 18142 15680 18198 15736
rect 18694 16788 18750 16824
rect 18694 16768 18696 16788
rect 18696 16768 18748 16788
rect 18748 16768 18750 16788
rect 18050 14864 18106 14920
rect 18050 13096 18106 13152
rect 18602 13368 18658 13424
rect 18142 11872 18198 11928
rect 18142 11348 18198 11384
rect 18142 11328 18144 11348
rect 18144 11328 18196 11348
rect 18196 11328 18198 11348
rect 18602 12144 18658 12200
rect 18234 11056 18290 11112
rect 18694 10512 18750 10568
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19614 20576 19670 20632
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 20074 20032 20130 20088
rect 19062 18028 19064 18048
rect 19064 18028 19116 18048
rect 19116 18028 19118 18048
rect 19062 17992 19118 18028
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 18878 16632 18934 16688
rect 18786 10240 18842 10296
rect 19062 13268 19064 13288
rect 19064 13268 19116 13288
rect 19116 13268 19118 13288
rect 19062 13232 19118 13268
rect 19982 18264 20038 18320
rect 19338 17720 19394 17776
rect 19246 16904 19302 16960
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19338 15952 19394 16008
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 21270 24792 21326 24848
rect 21546 24248 21602 24304
rect 21270 23568 21326 23624
rect 21914 23296 21970 23352
rect 21546 22752 21602 22808
rect 21822 22652 21824 22672
rect 21824 22652 21876 22672
rect 21876 22652 21878 22672
rect 21822 22616 21878 22652
rect 22742 24792 22798 24848
rect 22466 24248 22522 24304
rect 22374 23840 22430 23896
rect 22098 22480 22154 22536
rect 21362 21256 21418 21312
rect 21270 19896 21326 19952
rect 20810 19624 20866 19680
rect 20902 18808 20958 18864
rect 20810 18400 20866 18456
rect 20810 18128 20866 18184
rect 21086 18128 21142 18184
rect 20902 17448 20958 17504
rect 19246 14356 19248 14376
rect 19248 14356 19300 14376
rect 19300 14356 19302 14376
rect 19246 14320 19302 14356
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19430 14184 19486 14240
rect 19706 14220 19708 14240
rect 19708 14220 19760 14240
rect 19760 14220 19762 14240
rect 19706 14184 19762 14220
rect 19338 13912 19394 13968
rect 18510 8900 18566 8936
rect 18510 8880 18512 8900
rect 18512 8880 18564 8900
rect 18564 8880 18566 8900
rect 18878 8880 18934 8936
rect 18234 7792 18290 7848
rect 17590 6568 17646 6624
rect 18234 5072 18290 5128
rect 17406 4936 17462 4992
rect 17130 3984 17186 4040
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 20350 12824 20406 12880
rect 20074 11872 20130 11928
rect 19982 11600 20038 11656
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19982 10684 19984 10704
rect 19984 10684 20036 10704
rect 20036 10684 20038 10704
rect 19982 10648 20038 10684
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19982 9832 20038 9888
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19890 8508 19892 8528
rect 19892 8508 19944 8528
rect 19944 8508 19946 8528
rect 19890 8472 19946 8508
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19338 7964 19340 7984
rect 19340 7964 19392 7984
rect 19392 7964 19394 7984
rect 19154 6840 19210 6896
rect 19338 7928 19394 7964
rect 20350 10240 20406 10296
rect 20258 9560 20314 9616
rect 20626 12008 20682 12064
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 18786 5208 18842 5264
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 20902 15544 20958 15600
rect 20994 13912 21050 13968
rect 20902 8608 20958 8664
rect 20902 8356 20958 8392
rect 20902 8336 20904 8356
rect 20904 8336 20956 8356
rect 20956 8336 20958 8356
rect 20810 7928 20866 7984
rect 21086 12144 21142 12200
rect 21086 7812 21142 7848
rect 21086 7792 21088 7812
rect 21088 7792 21140 7812
rect 21140 7792 21142 7812
rect 21454 19352 21510 19408
rect 21270 16632 21326 16688
rect 21270 15000 21326 15056
rect 21270 13368 21326 13424
rect 21638 17176 21694 17232
rect 21914 21936 21970 21992
rect 21822 20168 21878 20224
rect 22098 18400 22154 18456
rect 22006 15000 22062 15056
rect 21914 13776 21970 13832
rect 21362 10648 21418 10704
rect 21270 8744 21326 8800
rect 21270 8472 21326 8528
rect 21822 10648 21878 10704
rect 22006 9460 22008 9480
rect 22008 9460 22060 9480
rect 22060 9460 22062 9480
rect 22006 9424 22062 9460
rect 21730 9288 21786 9344
rect 21546 8880 21602 8936
rect 21546 8608 21602 8664
rect 22558 21956 22614 21992
rect 22558 21936 22560 21956
rect 22560 21936 22612 21956
rect 22612 21936 22614 21956
rect 23018 24656 23074 24712
rect 23202 24676 23258 24712
rect 23202 24656 23204 24676
rect 23204 24656 23256 24676
rect 23256 24656 23258 24676
rect 22742 20984 22798 21040
rect 22374 16360 22430 16416
rect 22282 14340 22338 14376
rect 22282 14320 22284 14340
rect 22284 14320 22336 14340
rect 22336 14320 22338 14340
rect 22650 17856 22706 17912
rect 22650 14864 22706 14920
rect 22558 13504 22614 13560
rect 22558 12960 22614 13016
rect 22466 9560 22522 9616
rect 22834 18128 22890 18184
rect 22834 13932 22890 13968
rect 22834 13912 22836 13932
rect 22836 13912 22888 13932
rect 22888 13912 22890 13932
rect 22834 13640 22890 13696
rect 23202 23024 23258 23080
rect 23754 27104 23810 27160
rect 23570 24112 23626 24168
rect 23478 22752 23534 22808
rect 23478 21936 23534 21992
rect 23662 20848 23718 20904
rect 24214 26560 24270 26616
rect 24122 24792 24178 24848
rect 25226 26016 25282 26072
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24582 23704 24638 23760
rect 24398 23296 24454 23352
rect 25502 25336 25558 25392
rect 25410 24792 25466 24848
rect 24950 23568 25006 23624
rect 25410 23976 25466 24032
rect 24674 23160 24730 23216
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 25594 22480 25650 22536
rect 24122 20304 24178 20360
rect 23846 19216 23902 19272
rect 24122 20204 24124 20224
rect 24124 20204 24176 20224
rect 24176 20204 24178 20224
rect 24122 20168 24178 20204
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 20848 24822 20904
rect 24674 20460 24730 20496
rect 24674 20440 24676 20460
rect 24676 20440 24728 20460
rect 24728 20440 24730 20460
rect 23938 18944 23994 19000
rect 23938 18808 23994 18864
rect 23294 16904 23350 16960
rect 23386 15272 23442 15328
rect 23478 12960 23534 13016
rect 22926 11736 22982 11792
rect 22834 10920 22890 10976
rect 22742 9696 22798 9752
rect 22650 9016 22706 9072
rect 23754 18672 23810 18728
rect 23846 17312 23902 17368
rect 23754 16904 23810 16960
rect 24674 19624 24730 19680
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24122 16360 24178 16416
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24398 17040 24454 17096
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24122 15680 24178 15736
rect 23938 14456 23994 14512
rect 23754 13524 23810 13560
rect 23754 13504 23756 13524
rect 23756 13504 23808 13524
rect 23808 13504 23810 13524
rect 23662 12008 23718 12064
rect 23570 11600 23626 11656
rect 23478 11056 23534 11112
rect 22834 8880 22890 8936
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 25042 21292 25044 21312
rect 25044 21292 25096 21312
rect 25096 21292 25098 21312
rect 25042 21256 25098 21292
rect 25410 21936 25466 21992
rect 24766 17448 24822 17504
rect 24214 14592 24270 14648
rect 24122 13640 24178 13696
rect 24306 14356 24308 14376
rect 24308 14356 24360 14376
rect 24360 14356 24362 14376
rect 24306 14320 24362 14356
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 13912 24822 13968
rect 24306 13812 24308 13832
rect 24308 13812 24360 13832
rect 24360 13812 24362 13832
rect 24306 13776 24362 13812
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24306 12164 24362 12200
rect 24030 11872 24086 11928
rect 24306 12144 24308 12164
rect 24308 12144 24360 12164
rect 24360 12144 24362 12164
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24306 11056 24362 11112
rect 23846 9868 23848 9888
rect 23848 9868 23900 9888
rect 23900 9868 23902 9888
rect 23846 9832 23902 9868
rect 23754 9560 23810 9616
rect 23478 8744 23534 8800
rect 22282 6568 22338 6624
rect 20442 4664 20498 4720
rect 23570 8472 23626 8528
rect 23662 7384 23718 7440
rect 23846 9152 23902 9208
rect 23846 8336 23902 8392
rect 23754 7248 23810 7304
rect 23662 6704 23718 6760
rect 23570 5208 23626 5264
rect 23570 4528 23626 4584
rect 23478 4120 23534 4176
rect 20166 3848 20222 3904
rect 23478 3848 23534 3904
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 22190 3712 22246 3768
rect 18510 3576 18566 3632
rect 22006 3576 22062 3632
rect 23202 3440 23258 3496
rect 17038 3032 17094 3088
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14646 1536 14702 1592
rect 23570 2488 23626 2544
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24122 8608 24178 8664
rect 24122 7792 24178 7848
rect 23846 7112 23902 7168
rect 24122 2080 24178 2136
rect 24582 10260 24638 10296
rect 24582 10240 24584 10260
rect 24584 10240 24636 10260
rect 24636 10240 24638 10260
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24674 9152 24730 9208
rect 25318 21428 25320 21448
rect 25320 21428 25372 21448
rect 25372 21428 25374 21448
rect 25318 21392 25374 21428
rect 25226 20712 25282 20768
rect 25502 21392 25558 21448
rect 25226 20032 25282 20088
rect 25318 19796 25320 19816
rect 25320 19796 25372 19816
rect 25372 19796 25374 19816
rect 25318 19760 25374 19796
rect 25042 16940 25044 16960
rect 25044 16940 25096 16960
rect 25096 16940 25098 16960
rect 25042 16904 25098 16940
rect 25134 16768 25190 16824
rect 25502 16224 25558 16280
rect 24950 15408 25006 15464
rect 24950 12824 25006 12880
rect 24950 11212 25006 11248
rect 24950 11192 24952 11212
rect 24952 11192 25004 11212
rect 25004 11192 25006 11212
rect 25134 10920 25190 10976
rect 25410 12824 25466 12880
rect 25318 12688 25374 12744
rect 25410 12280 25466 12336
rect 25318 10920 25374 10976
rect 24858 9288 24914 9344
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23754 1944 23810 2000
rect 23478 856 23534 912
rect 3238 312 3294 368
rect 24766 9016 24822 9072
rect 25226 10648 25282 10704
rect 27066 24792 27122 24848
rect 27618 23976 27674 24032
rect 26238 18672 26294 18728
rect 25594 13232 25650 13288
rect 24766 7948 24822 7984
rect 24766 7928 24768 7948
rect 24768 7928 24820 7948
rect 24820 7928 24822 7948
rect 24674 312 24730 368
<< metal3 >>
rect 0 27706 480 27736
rect 4429 27706 4495 27709
rect 0 27704 4495 27706
rect 0 27648 4434 27704
rect 4490 27648 4495 27704
rect 0 27646 4495 27648
rect 0 27616 480 27646
rect 4429 27643 4495 27646
rect 23933 27706 23999 27709
rect 27520 27706 28000 27736
rect 23933 27704 28000 27706
rect 23933 27648 23938 27704
rect 23994 27648 28000 27704
rect 23933 27646 28000 27648
rect 23933 27643 23999 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 4797 27162 4863 27165
rect 0 27160 4863 27162
rect 0 27104 4802 27160
rect 4858 27104 4863 27160
rect 0 27102 4863 27104
rect 0 27072 480 27102
rect 4797 27099 4863 27102
rect 23749 27162 23815 27165
rect 27520 27162 28000 27192
rect 23749 27160 28000 27162
rect 23749 27104 23754 27160
rect 23810 27104 28000 27160
rect 23749 27102 28000 27104
rect 23749 27099 23815 27102
rect 27520 27072 28000 27102
rect 0 26618 480 26648
rect 1209 26618 1275 26621
rect 0 26616 1275 26618
rect 0 26560 1214 26616
rect 1270 26560 1275 26616
rect 0 26558 1275 26560
rect 0 26528 480 26558
rect 1209 26555 1275 26558
rect 24209 26618 24275 26621
rect 27520 26618 28000 26648
rect 24209 26616 28000 26618
rect 24209 26560 24214 26616
rect 24270 26560 28000 26616
rect 24209 26558 28000 26560
rect 24209 26555 24275 26558
rect 27520 26528 28000 26558
rect 0 26074 480 26104
rect 3049 26074 3115 26077
rect 0 26072 3115 26074
rect 0 26016 3054 26072
rect 3110 26016 3115 26072
rect 0 26014 3115 26016
rect 0 25984 480 26014
rect 3049 26011 3115 26014
rect 25221 26074 25287 26077
rect 27520 26074 28000 26104
rect 25221 26072 28000 26074
rect 25221 26016 25226 26072
rect 25282 26016 28000 26072
rect 25221 26014 28000 26016
rect 25221 26011 25287 26014
rect 27520 25984 28000 26014
rect 11973 25802 12039 25805
rect 12801 25802 12867 25805
rect 11973 25800 12867 25802
rect 11973 25744 11978 25800
rect 12034 25744 12806 25800
rect 12862 25744 12867 25800
rect 11973 25742 12867 25744
rect 11973 25739 12039 25742
rect 12801 25739 12867 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 1669 25394 1735 25397
rect 0 25392 1735 25394
rect 0 25336 1674 25392
rect 1730 25336 1735 25392
rect 0 25334 1735 25336
rect 0 25304 480 25334
rect 1669 25331 1735 25334
rect 12157 25394 12223 25397
rect 15469 25394 15535 25397
rect 12157 25392 15535 25394
rect 12157 25336 12162 25392
rect 12218 25336 15474 25392
rect 15530 25336 15535 25392
rect 12157 25334 15535 25336
rect 12157 25331 12223 25334
rect 15469 25331 15535 25334
rect 25497 25394 25563 25397
rect 27520 25394 28000 25424
rect 25497 25392 28000 25394
rect 25497 25336 25502 25392
rect 25558 25336 28000 25392
rect 25497 25334 28000 25336
rect 25497 25331 25563 25334
rect 27520 25304 28000 25334
rect 2497 25258 2563 25261
rect 5901 25258 5967 25261
rect 2497 25256 5967 25258
rect 2497 25200 2502 25256
rect 2558 25200 5906 25256
rect 5962 25200 5967 25256
rect 2497 25198 5967 25200
rect 2497 25195 2563 25198
rect 5901 25195 5967 25198
rect 10409 25258 10475 25261
rect 18873 25258 18939 25261
rect 10409 25256 18939 25258
rect 10409 25200 10414 25256
rect 10470 25200 18878 25256
rect 18934 25200 18939 25256
rect 10409 25198 18939 25200
rect 10409 25195 10475 25198
rect 18873 25195 18939 25198
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 2957 24986 3023 24989
rect 6085 24986 6151 24989
rect 9438 24986 9444 24988
rect 2957 24984 3066 24986
rect 2957 24928 2962 24984
rect 3018 24928 3066 24984
rect 2957 24923 3066 24928
rect 6085 24984 9444 24986
rect 6085 24928 6090 24984
rect 6146 24928 9444 24984
rect 6085 24926 9444 24928
rect 6085 24923 6151 24926
rect 9438 24924 9444 24926
rect 9508 24924 9514 24988
rect 0 24850 480 24880
rect 1301 24850 1367 24853
rect 0 24848 1367 24850
rect 0 24792 1306 24848
rect 1362 24792 1367 24848
rect 0 24790 1367 24792
rect 0 24760 480 24790
rect 1301 24787 1367 24790
rect 2313 24850 2379 24853
rect 3006 24850 3066 24923
rect 6821 24850 6887 24853
rect 2313 24848 6887 24850
rect 2313 24792 2318 24848
rect 2374 24792 6826 24848
rect 6882 24792 6887 24848
rect 2313 24790 6887 24792
rect 2313 24787 2379 24790
rect 6821 24787 6887 24790
rect 7281 24850 7347 24853
rect 11145 24850 11211 24853
rect 7281 24848 11211 24850
rect 7281 24792 7286 24848
rect 7342 24792 11150 24848
rect 11206 24792 11211 24848
rect 7281 24790 11211 24792
rect 7281 24787 7347 24790
rect 11145 24787 11211 24790
rect 11789 24850 11855 24853
rect 15653 24850 15719 24853
rect 17125 24850 17191 24853
rect 11789 24848 15578 24850
rect 11789 24792 11794 24848
rect 11850 24792 15578 24848
rect 11789 24790 15578 24792
rect 11789 24787 11855 24790
rect 5993 24714 6059 24717
rect 8109 24714 8175 24717
rect 5993 24712 8175 24714
rect 5993 24656 5998 24712
rect 6054 24656 8114 24712
rect 8170 24656 8175 24712
rect 5993 24654 8175 24656
rect 5993 24651 6059 24654
rect 8109 24651 8175 24654
rect 10685 24714 10751 24717
rect 12893 24714 12959 24717
rect 10685 24712 12959 24714
rect 10685 24656 10690 24712
rect 10746 24656 12898 24712
rect 12954 24656 12959 24712
rect 10685 24654 12959 24656
rect 10685 24651 10751 24654
rect 12893 24651 12959 24654
rect 3325 24578 3391 24581
rect 10133 24578 10199 24581
rect 3325 24576 10199 24578
rect 3325 24520 3330 24576
rect 3386 24520 10138 24576
rect 10194 24520 10199 24576
rect 3325 24518 10199 24520
rect 15518 24578 15578 24790
rect 15653 24848 17191 24850
rect 15653 24792 15658 24848
rect 15714 24792 17130 24848
rect 17186 24792 17191 24848
rect 15653 24790 17191 24792
rect 15653 24787 15719 24790
rect 17125 24787 17191 24790
rect 19241 24850 19307 24853
rect 21265 24850 21331 24853
rect 19241 24848 21331 24850
rect 19241 24792 19246 24848
rect 19302 24792 21270 24848
rect 21326 24792 21331 24848
rect 19241 24790 21331 24792
rect 19241 24787 19307 24790
rect 21265 24787 21331 24790
rect 22737 24850 22803 24853
rect 24117 24850 24183 24853
rect 22737 24848 24183 24850
rect 22737 24792 22742 24848
rect 22798 24792 24122 24848
rect 24178 24792 24183 24848
rect 22737 24790 24183 24792
rect 22737 24787 22803 24790
rect 24117 24787 24183 24790
rect 25405 24850 25471 24853
rect 27061 24850 27127 24853
rect 27520 24850 28000 24880
rect 25405 24848 27127 24850
rect 25405 24792 25410 24848
rect 25466 24792 27066 24848
rect 27122 24792 27127 24848
rect 25405 24790 27127 24792
rect 25405 24787 25471 24790
rect 27061 24787 27127 24790
rect 27294 24790 28000 24850
rect 16757 24714 16823 24717
rect 23013 24714 23079 24717
rect 16757 24712 23079 24714
rect 16757 24656 16762 24712
rect 16818 24656 23018 24712
rect 23074 24656 23079 24712
rect 16757 24654 23079 24656
rect 16757 24651 16823 24654
rect 23013 24651 23079 24654
rect 23197 24714 23263 24717
rect 27294 24714 27354 24790
rect 27520 24760 28000 24790
rect 23197 24712 27354 24714
rect 23197 24656 23202 24712
rect 23258 24656 27354 24712
rect 23197 24654 27354 24656
rect 23197 24651 23263 24654
rect 17033 24578 17099 24581
rect 15518 24576 17099 24578
rect 15518 24520 17038 24576
rect 17094 24520 17099 24576
rect 15518 24518 17099 24520
rect 3325 24515 3391 24518
rect 10133 24515 10199 24518
rect 17033 24515 17099 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 10041 24442 10107 24445
rect 6318 24440 10107 24442
rect 6318 24384 10046 24440
rect 10102 24384 10107 24440
rect 6318 24382 10107 24384
rect 0 24306 480 24336
rect 3785 24306 3851 24309
rect 6318 24306 6378 24382
rect 10041 24379 10107 24382
rect 15837 24442 15903 24445
rect 18229 24442 18295 24445
rect 15837 24440 18295 24442
rect 15837 24384 15842 24440
rect 15898 24384 18234 24440
rect 18290 24384 18295 24440
rect 15837 24382 18295 24384
rect 15837 24379 15903 24382
rect 18229 24379 18295 24382
rect 0 24304 3851 24306
rect 0 24248 3790 24304
rect 3846 24248 3851 24304
rect 0 24246 3851 24248
rect 0 24216 480 24246
rect 3785 24243 3851 24246
rect 3926 24246 6378 24306
rect 7281 24306 7347 24309
rect 10961 24306 11027 24309
rect 7281 24304 11027 24306
rect 7281 24248 7286 24304
rect 7342 24248 10966 24304
rect 11022 24248 11027 24304
rect 7281 24246 11027 24248
rect 3601 24170 3667 24173
rect 3926 24170 3986 24246
rect 7281 24243 7347 24246
rect 10961 24243 11027 24246
rect 13353 24306 13419 24309
rect 21541 24306 21607 24309
rect 13353 24304 21607 24306
rect 13353 24248 13358 24304
rect 13414 24248 21546 24304
rect 21602 24248 21607 24304
rect 13353 24246 21607 24248
rect 13353 24243 13419 24246
rect 21541 24243 21607 24246
rect 22461 24306 22527 24309
rect 27520 24306 28000 24336
rect 22461 24304 28000 24306
rect 22461 24248 22466 24304
rect 22522 24248 28000 24304
rect 22461 24246 28000 24248
rect 22461 24243 22527 24246
rect 27520 24216 28000 24246
rect 3601 24168 3986 24170
rect 3601 24112 3606 24168
rect 3662 24112 3986 24168
rect 3601 24110 3986 24112
rect 5349 24170 5415 24173
rect 7925 24170 7991 24173
rect 5349 24168 7991 24170
rect 5349 24112 5354 24168
rect 5410 24112 7930 24168
rect 7986 24112 7991 24168
rect 5349 24110 7991 24112
rect 3601 24107 3667 24110
rect 5349 24107 5415 24110
rect 7925 24107 7991 24110
rect 9622 24108 9628 24172
rect 9692 24170 9698 24172
rect 12709 24170 12775 24173
rect 9692 24168 12775 24170
rect 9692 24112 12714 24168
rect 12770 24112 12775 24168
rect 9692 24110 12775 24112
rect 9692 24108 9698 24110
rect 12709 24107 12775 24110
rect 14273 24170 14339 24173
rect 23565 24170 23631 24173
rect 14273 24168 23631 24170
rect 14273 24112 14278 24168
rect 14334 24112 23570 24168
rect 23626 24112 23631 24168
rect 14273 24110 23631 24112
rect 14273 24107 14339 24110
rect 23565 24107 23631 24110
rect 25405 24034 25471 24037
rect 27613 24034 27679 24037
rect 25405 24032 27679 24034
rect 25405 23976 25410 24032
rect 25466 23976 27618 24032
rect 27674 23976 27679 24032
rect 25405 23974 27679 23976
rect 25405 23971 25471 23974
rect 27613 23971 27679 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10133 23898 10199 23901
rect 12065 23898 12131 23901
rect 10133 23896 12131 23898
rect 10133 23840 10138 23896
rect 10194 23840 12070 23896
rect 12126 23840 12131 23896
rect 10133 23838 12131 23840
rect 10133 23835 10199 23838
rect 12065 23835 12131 23838
rect 12249 23898 12315 23901
rect 14733 23898 14799 23901
rect 12249 23896 14799 23898
rect 12249 23840 12254 23896
rect 12310 23840 14738 23896
rect 14794 23840 14799 23896
rect 12249 23838 14799 23840
rect 12249 23835 12315 23838
rect 14733 23835 14799 23838
rect 19885 23898 19951 23901
rect 22369 23898 22435 23901
rect 19885 23896 22435 23898
rect 19885 23840 19890 23896
rect 19946 23840 22374 23896
rect 22430 23840 22435 23896
rect 19885 23838 22435 23840
rect 19885 23835 19951 23838
rect 22369 23835 22435 23838
rect 0 23762 480 23792
rect 2037 23762 2103 23765
rect 6637 23762 6703 23765
rect 0 23702 1226 23762
rect 0 23672 480 23702
rect 1166 23490 1226 23702
rect 2037 23760 6703 23762
rect 2037 23704 2042 23760
rect 2098 23704 6642 23760
rect 6698 23704 6703 23760
rect 2037 23702 6703 23704
rect 2037 23699 2103 23702
rect 6637 23699 6703 23702
rect 6821 23762 6887 23765
rect 9397 23762 9463 23765
rect 11789 23762 11855 23765
rect 6821 23760 11855 23762
rect 6821 23704 6826 23760
rect 6882 23704 9402 23760
rect 9458 23704 11794 23760
rect 11850 23704 11855 23760
rect 6821 23702 11855 23704
rect 6821 23699 6887 23702
rect 9397 23699 9463 23702
rect 11789 23699 11855 23702
rect 12801 23762 12867 23765
rect 16389 23762 16455 23765
rect 16849 23762 16915 23765
rect 12801 23760 16915 23762
rect 12801 23704 12806 23760
rect 12862 23704 16394 23760
rect 16450 23704 16854 23760
rect 16910 23704 16915 23760
rect 12801 23702 16915 23704
rect 12801 23699 12867 23702
rect 16389 23699 16455 23702
rect 16849 23699 16915 23702
rect 20345 23762 20411 23765
rect 24577 23762 24643 23765
rect 27520 23762 28000 23792
rect 20345 23760 28000 23762
rect 20345 23704 20350 23760
rect 20406 23704 24582 23760
rect 24638 23704 28000 23760
rect 20345 23702 28000 23704
rect 20345 23699 20411 23702
rect 24577 23699 24643 23702
rect 27520 23672 28000 23702
rect 8109 23626 8175 23629
rect 17769 23626 17835 23629
rect 8109 23624 17835 23626
rect 8109 23568 8114 23624
rect 8170 23568 17774 23624
rect 17830 23568 17835 23624
rect 8109 23566 17835 23568
rect 8109 23563 8175 23566
rect 17769 23563 17835 23566
rect 21265 23626 21331 23629
rect 24945 23626 25011 23629
rect 21265 23624 25011 23626
rect 21265 23568 21270 23624
rect 21326 23568 24950 23624
rect 25006 23568 25011 23624
rect 21265 23566 25011 23568
rect 21265 23563 21331 23566
rect 24945 23563 25011 23566
rect 2865 23490 2931 23493
rect 1166 23488 2931 23490
rect 1166 23432 2870 23488
rect 2926 23432 2931 23488
rect 1166 23430 2931 23432
rect 2865 23427 2931 23430
rect 4061 23490 4127 23493
rect 7833 23490 7899 23493
rect 8661 23490 8727 23493
rect 11053 23492 11119 23493
rect 11053 23490 11100 23492
rect 4061 23488 8727 23490
rect 4061 23432 4066 23488
rect 4122 23432 7838 23488
rect 7894 23432 8666 23488
rect 8722 23432 8727 23488
rect 4061 23430 8727 23432
rect 11008 23488 11100 23490
rect 11008 23432 11058 23488
rect 11008 23430 11100 23432
rect 4061 23427 4127 23430
rect 7833 23427 7899 23430
rect 8661 23427 8727 23430
rect 11053 23428 11100 23430
rect 11164 23428 11170 23492
rect 13721 23490 13787 23493
rect 18045 23490 18111 23493
rect 13721 23488 18111 23490
rect 13721 23432 13726 23488
rect 13782 23432 18050 23488
rect 18106 23432 18111 23488
rect 13721 23430 18111 23432
rect 11053 23427 11119 23428
rect 13721 23427 13787 23430
rect 18045 23427 18111 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 2957 23354 3023 23357
rect 5993 23354 6059 23357
rect 2957 23352 6059 23354
rect 2957 23296 2962 23352
rect 3018 23296 5998 23352
rect 6054 23296 6059 23352
rect 2957 23294 6059 23296
rect 2957 23291 3023 23294
rect 5993 23291 6059 23294
rect 14273 23354 14339 23357
rect 16665 23354 16731 23357
rect 14273 23352 16731 23354
rect 14273 23296 14278 23352
rect 14334 23296 16670 23352
rect 16726 23296 16731 23352
rect 14273 23294 16731 23296
rect 14273 23291 14339 23294
rect 16665 23291 16731 23294
rect 21909 23354 21975 23357
rect 24393 23354 24459 23357
rect 21909 23352 24459 23354
rect 21909 23296 21914 23352
rect 21970 23296 24398 23352
rect 24454 23296 24459 23352
rect 21909 23294 24459 23296
rect 21909 23291 21975 23294
rect 24393 23291 24459 23294
rect 0 23218 480 23248
rect 3049 23218 3115 23221
rect 0 23216 3115 23218
rect 0 23160 3054 23216
rect 3110 23160 3115 23216
rect 0 23158 3115 23160
rect 0 23128 480 23158
rect 3049 23155 3115 23158
rect 3233 23218 3299 23221
rect 6913 23218 6979 23221
rect 3233 23216 6979 23218
rect 3233 23160 3238 23216
rect 3294 23160 6918 23216
rect 6974 23160 6979 23216
rect 3233 23158 6979 23160
rect 3233 23155 3299 23158
rect 6913 23155 6979 23158
rect 10133 23218 10199 23221
rect 17953 23218 18019 23221
rect 10133 23216 18019 23218
rect 10133 23160 10138 23216
rect 10194 23160 17958 23216
rect 18014 23160 18019 23216
rect 10133 23158 18019 23160
rect 10133 23155 10199 23158
rect 17953 23155 18019 23158
rect 24669 23218 24735 23221
rect 27520 23218 28000 23248
rect 24669 23216 28000 23218
rect 24669 23160 24674 23216
rect 24730 23160 28000 23216
rect 24669 23158 28000 23160
rect 24669 23155 24735 23158
rect 27520 23128 28000 23158
rect 2405 23082 2471 23085
rect 5993 23082 6059 23085
rect 2405 23080 6059 23082
rect 2405 23024 2410 23080
rect 2466 23024 5998 23080
rect 6054 23024 6059 23080
rect 2405 23022 6059 23024
rect 2405 23019 2471 23022
rect 5993 23019 6059 23022
rect 8753 23082 8819 23085
rect 11094 23082 11100 23084
rect 8753 23080 11100 23082
rect 8753 23024 8758 23080
rect 8814 23024 11100 23080
rect 8753 23022 11100 23024
rect 8753 23019 8819 23022
rect 11094 23020 11100 23022
rect 11164 23020 11170 23084
rect 13537 23082 13603 23085
rect 15285 23082 15351 23085
rect 13537 23080 15351 23082
rect 13537 23024 13542 23080
rect 13598 23024 15290 23080
rect 15346 23024 15351 23080
rect 13537 23022 15351 23024
rect 13537 23019 13603 23022
rect 15285 23019 15351 23022
rect 17401 23082 17467 23085
rect 23197 23082 23263 23085
rect 17401 23080 23263 23082
rect 17401 23024 17406 23080
rect 17462 23024 23202 23080
rect 23258 23024 23263 23080
rect 17401 23022 23263 23024
rect 17401 23019 17467 23022
rect 23197 23019 23263 23022
rect 6729 22946 6795 22949
rect 9949 22946 10015 22949
rect 10133 22946 10199 22949
rect 6729 22944 10199 22946
rect 6729 22888 6734 22944
rect 6790 22888 9954 22944
rect 10010 22888 10138 22944
rect 10194 22888 10199 22944
rect 6729 22886 10199 22888
rect 6729 22883 6795 22886
rect 9949 22883 10015 22886
rect 10133 22883 10199 22886
rect 10961 22946 11027 22949
rect 13629 22946 13695 22949
rect 10961 22944 13695 22946
rect 10961 22888 10966 22944
rect 11022 22888 13634 22944
rect 13690 22888 13695 22944
rect 10961 22886 13695 22888
rect 10961 22883 11027 22886
rect 13629 22883 13695 22886
rect 18505 22946 18571 22949
rect 20621 22946 20687 22949
rect 18505 22944 20687 22946
rect 18505 22888 18510 22944
rect 18566 22888 20626 22944
rect 20682 22888 20687 22944
rect 18505 22886 20687 22888
rect 18505 22883 18571 22886
rect 20621 22883 20687 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 6085 22810 6151 22813
rect 7465 22810 7531 22813
rect 6085 22808 7531 22810
rect 6085 22752 6090 22808
rect 6146 22752 7470 22808
rect 7526 22752 7531 22808
rect 6085 22750 7531 22752
rect 6085 22747 6151 22750
rect 7465 22747 7531 22750
rect 7833 22810 7899 22813
rect 19701 22810 19767 22813
rect 21541 22810 21607 22813
rect 23473 22810 23539 22813
rect 7833 22808 13876 22810
rect 7833 22752 7838 22808
rect 7894 22752 13876 22808
rect 7833 22750 13876 22752
rect 7833 22747 7899 22750
rect 1945 22674 2011 22677
rect 11329 22674 11395 22677
rect 13537 22674 13603 22677
rect 1945 22672 7666 22674
rect 1945 22616 1950 22672
rect 2006 22616 7666 22672
rect 1945 22614 7666 22616
rect 1945 22611 2011 22614
rect 0 22538 480 22568
rect 7606 22538 7666 22614
rect 11329 22672 13603 22674
rect 11329 22616 11334 22672
rect 11390 22616 13542 22672
rect 13598 22616 13603 22672
rect 11329 22614 13603 22616
rect 13816 22674 13876 22750
rect 19701 22808 23539 22810
rect 19701 22752 19706 22808
rect 19762 22752 21546 22808
rect 21602 22752 23478 22808
rect 23534 22752 23539 22808
rect 19701 22750 23539 22752
rect 19701 22747 19767 22750
rect 21541 22747 21607 22750
rect 23473 22747 23539 22750
rect 15285 22674 15351 22677
rect 13816 22672 15351 22674
rect 13816 22616 15290 22672
rect 15346 22616 15351 22672
rect 13816 22614 15351 22616
rect 11329 22611 11395 22614
rect 13537 22611 13603 22614
rect 15285 22611 15351 22614
rect 15745 22674 15811 22677
rect 21817 22674 21883 22677
rect 15745 22672 21883 22674
rect 15745 22616 15750 22672
rect 15806 22616 21822 22672
rect 21878 22616 21883 22672
rect 15745 22614 21883 22616
rect 15745 22611 15811 22614
rect 21817 22611 21883 22614
rect 14089 22538 14155 22541
rect 0 22478 5826 22538
rect 7606 22536 14155 22538
rect 7606 22480 14094 22536
rect 14150 22480 14155 22536
rect 7606 22478 14155 22480
rect 0 22448 480 22478
rect 1761 22402 1827 22405
rect 5533 22402 5599 22405
rect 1761 22400 5599 22402
rect 1761 22344 1766 22400
rect 1822 22344 5538 22400
rect 5594 22344 5599 22400
rect 1761 22342 5599 22344
rect 5766 22402 5826 22478
rect 14089 22475 14155 22478
rect 14825 22538 14891 22541
rect 18689 22538 18755 22541
rect 14825 22536 18755 22538
rect 14825 22480 14830 22536
rect 14886 22480 18694 22536
rect 18750 22480 18755 22536
rect 14825 22478 18755 22480
rect 14825 22475 14891 22478
rect 18689 22475 18755 22478
rect 19885 22538 19951 22541
rect 22093 22538 22159 22541
rect 19885 22536 22159 22538
rect 19885 22480 19890 22536
rect 19946 22480 22098 22536
rect 22154 22480 22159 22536
rect 19885 22478 22159 22480
rect 19885 22475 19951 22478
rect 22093 22475 22159 22478
rect 25589 22538 25655 22541
rect 27520 22538 28000 22568
rect 25589 22536 28000 22538
rect 25589 22480 25594 22536
rect 25650 22480 28000 22536
rect 25589 22478 28000 22480
rect 25589 22475 25655 22478
rect 27520 22448 28000 22478
rect 8293 22402 8359 22405
rect 5766 22400 8359 22402
rect 5766 22344 8298 22400
rect 8354 22344 8359 22400
rect 5766 22342 8359 22344
rect 1761 22339 1827 22342
rect 5533 22339 5599 22342
rect 8293 22339 8359 22342
rect 13629 22402 13695 22405
rect 19333 22402 19399 22405
rect 13629 22400 19399 22402
rect 13629 22344 13634 22400
rect 13690 22344 19338 22400
rect 19394 22344 19399 22400
rect 13629 22342 19399 22344
rect 13629 22339 13695 22342
rect 19333 22339 19399 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 10685 22266 10751 22269
rect 19425 22266 19491 22269
rect 10685 22264 19491 22266
rect 10685 22208 10690 22264
rect 10746 22208 19430 22264
rect 19486 22208 19491 22264
rect 10685 22206 19491 22208
rect 10685 22203 10751 22206
rect 19425 22203 19491 22206
rect 9857 22130 9923 22133
rect 12617 22130 12683 22133
rect 9857 22128 12683 22130
rect 9857 22072 9862 22128
rect 9918 22072 12622 22128
rect 12678 22072 12683 22128
rect 9857 22070 12683 22072
rect 9857 22067 9923 22070
rect 12617 22067 12683 22070
rect 15469 22096 15535 22099
rect 15469 22094 15578 22096
rect 15469 22038 15474 22094
rect 15530 22038 15578 22094
rect 15469 22033 15578 22038
rect 0 21994 480 22024
rect 7005 21994 7071 21997
rect 0 21992 7071 21994
rect 0 21936 7010 21992
rect 7066 21936 7071 21992
rect 0 21934 7071 21936
rect 15518 21994 15578 22033
rect 15745 21994 15811 21997
rect 15518 21992 15811 21994
rect 15518 21936 15750 21992
rect 15806 21936 15811 21992
rect 15518 21934 15811 21936
rect 0 21904 480 21934
rect 7005 21931 7071 21934
rect 15745 21931 15811 21934
rect 17401 21994 17467 21997
rect 19701 21994 19767 21997
rect 17401 21992 19767 21994
rect 17401 21936 17406 21992
rect 17462 21936 19706 21992
rect 19762 21936 19767 21992
rect 17401 21934 19767 21936
rect 17401 21931 17467 21934
rect 19701 21931 19767 21934
rect 21909 21994 21975 21997
rect 22553 21994 22619 21997
rect 23473 21994 23539 21997
rect 21909 21992 23539 21994
rect 21909 21936 21914 21992
rect 21970 21936 22558 21992
rect 22614 21936 23478 21992
rect 23534 21936 23539 21992
rect 21909 21934 23539 21936
rect 21909 21931 21975 21934
rect 22553 21931 22619 21934
rect 23473 21931 23539 21934
rect 25405 21994 25471 21997
rect 27520 21994 28000 22024
rect 25405 21992 28000 21994
rect 25405 21936 25410 21992
rect 25466 21936 28000 21992
rect 25405 21934 28000 21936
rect 25405 21931 25471 21934
rect 27520 21904 28000 21934
rect 6453 21858 6519 21861
rect 11513 21858 11579 21861
rect 6453 21856 11579 21858
rect 6453 21800 6458 21856
rect 6514 21800 11518 21856
rect 11574 21800 11579 21856
rect 6453 21798 11579 21800
rect 6453 21795 6519 21798
rect 11513 21795 11579 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 10961 21722 11027 21725
rect 14089 21722 14155 21725
rect 10961 21720 14155 21722
rect 10961 21664 10966 21720
rect 11022 21664 14094 21720
rect 14150 21664 14155 21720
rect 10961 21662 14155 21664
rect 10961 21659 11027 21662
rect 14089 21659 14155 21662
rect 4521 21586 4587 21589
rect 8293 21586 8359 21589
rect 4521 21584 8359 21586
rect 4521 21528 4526 21584
rect 4582 21528 8298 21584
rect 8354 21528 8359 21584
rect 4521 21526 8359 21528
rect 4521 21523 4587 21526
rect 8293 21523 8359 21526
rect 10961 21586 11027 21589
rect 11789 21586 11855 21589
rect 19241 21586 19307 21589
rect 10961 21584 19307 21586
rect 10961 21528 10966 21584
rect 11022 21528 11794 21584
rect 11850 21528 19246 21584
rect 19302 21528 19307 21584
rect 10961 21526 19307 21528
rect 10961 21523 11027 21526
rect 11789 21523 11855 21526
rect 19241 21523 19307 21526
rect 0 21450 480 21480
rect 2957 21450 3023 21453
rect 0 21448 3023 21450
rect 0 21392 2962 21448
rect 3018 21392 3023 21448
rect 0 21390 3023 21392
rect 0 21360 480 21390
rect 2957 21387 3023 21390
rect 3877 21450 3943 21453
rect 6913 21450 6979 21453
rect 3877 21448 6979 21450
rect 3877 21392 3882 21448
rect 3938 21392 6918 21448
rect 6974 21392 6979 21448
rect 3877 21390 6979 21392
rect 3877 21387 3943 21390
rect 6913 21387 6979 21390
rect 7189 21450 7255 21453
rect 12617 21450 12683 21453
rect 7189 21448 12683 21450
rect 7189 21392 7194 21448
rect 7250 21392 12622 21448
rect 12678 21392 12683 21448
rect 7189 21390 12683 21392
rect 7189 21387 7255 21390
rect 12617 21387 12683 21390
rect 15745 21450 15811 21453
rect 25313 21450 25379 21453
rect 15745 21448 25379 21450
rect 15745 21392 15750 21448
rect 15806 21392 25318 21448
rect 25374 21392 25379 21448
rect 15745 21390 25379 21392
rect 15745 21387 15811 21390
rect 25313 21387 25379 21390
rect 25497 21450 25563 21453
rect 27520 21450 28000 21480
rect 25497 21448 28000 21450
rect 25497 21392 25502 21448
rect 25558 21392 28000 21448
rect 25497 21390 28000 21392
rect 25497 21387 25563 21390
rect 27520 21360 28000 21390
rect 2405 21314 2471 21317
rect 4613 21314 4679 21317
rect 8569 21314 8635 21317
rect 2405 21312 8635 21314
rect 2405 21256 2410 21312
rect 2466 21256 4618 21312
rect 4674 21256 8574 21312
rect 8630 21256 8635 21312
rect 2405 21254 8635 21256
rect 2405 21251 2471 21254
rect 4613 21251 4679 21254
rect 8569 21251 8635 21254
rect 11513 21314 11579 21317
rect 12065 21314 12131 21317
rect 16297 21314 16363 21317
rect 11513 21312 16363 21314
rect 11513 21256 11518 21312
rect 11574 21256 12070 21312
rect 12126 21256 16302 21312
rect 16358 21256 16363 21312
rect 11513 21254 16363 21256
rect 11513 21251 11579 21254
rect 12065 21251 12131 21254
rect 16297 21251 16363 21254
rect 21357 21314 21423 21317
rect 25037 21314 25103 21317
rect 21357 21312 25103 21314
rect 21357 21256 21362 21312
rect 21418 21256 25042 21312
rect 25098 21256 25103 21312
rect 21357 21254 25103 21256
rect 21357 21251 21423 21254
rect 25037 21251 25103 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1577 21178 1643 21181
rect 6361 21178 6427 21181
rect 1577 21176 6427 21178
rect 1577 21120 1582 21176
rect 1638 21120 6366 21176
rect 6422 21120 6427 21176
rect 1577 21118 6427 21120
rect 1577 21115 1643 21118
rect 6361 21115 6427 21118
rect 6913 21178 6979 21181
rect 9622 21178 9628 21180
rect 6913 21176 9628 21178
rect 6913 21120 6918 21176
rect 6974 21120 9628 21176
rect 6913 21118 9628 21120
rect 6913 21115 6979 21118
rect 9622 21116 9628 21118
rect 9692 21116 9698 21180
rect 11513 21178 11579 21181
rect 10688 21176 11579 21178
rect 10688 21120 11518 21176
rect 11574 21120 11579 21176
rect 10688 21118 11579 21120
rect 3325 21042 3391 21045
rect 10688 21042 10748 21118
rect 11513 21115 11579 21118
rect 3325 21040 10748 21042
rect 3325 20984 3330 21040
rect 3386 20984 10748 21040
rect 3325 20982 10748 20984
rect 10869 21042 10935 21045
rect 14549 21042 14615 21045
rect 10869 21040 14615 21042
rect 10869 20984 10874 21040
rect 10930 20984 14554 21040
rect 14610 20984 14615 21040
rect 10869 20982 14615 20984
rect 3325 20979 3391 20982
rect 10869 20979 10935 20982
rect 14549 20979 14615 20982
rect 16757 21042 16823 21045
rect 22737 21042 22803 21045
rect 16757 21040 22803 21042
rect 16757 20984 16762 21040
rect 16818 20984 22742 21040
rect 22798 20984 22803 21040
rect 16757 20982 22803 20984
rect 16757 20979 16823 20982
rect 22737 20979 22803 20982
rect 0 20906 480 20936
rect 3877 20906 3943 20909
rect 0 20904 3943 20906
rect 0 20848 3882 20904
rect 3938 20848 3943 20904
rect 0 20846 3943 20848
rect 0 20816 480 20846
rect 3877 20843 3943 20846
rect 4061 20906 4127 20909
rect 7005 20906 7071 20909
rect 4061 20904 7071 20906
rect 4061 20848 4066 20904
rect 4122 20848 7010 20904
rect 7066 20848 7071 20904
rect 4061 20846 7071 20848
rect 4061 20843 4127 20846
rect 7005 20843 7071 20846
rect 7189 20906 7255 20909
rect 12801 20906 12867 20909
rect 7189 20904 12867 20906
rect 7189 20848 7194 20904
rect 7250 20848 12806 20904
rect 12862 20848 12867 20904
rect 7189 20846 12867 20848
rect 7189 20843 7255 20846
rect 12801 20843 12867 20846
rect 14825 20906 14891 20909
rect 23657 20906 23723 20909
rect 14825 20904 23723 20906
rect 14825 20848 14830 20904
rect 14886 20848 23662 20904
rect 23718 20848 23723 20904
rect 14825 20846 23723 20848
rect 14825 20843 14891 20846
rect 23657 20843 23723 20846
rect 24761 20906 24827 20909
rect 27520 20906 28000 20936
rect 24761 20904 28000 20906
rect 24761 20848 24766 20904
rect 24822 20848 28000 20904
rect 24761 20846 28000 20848
rect 24761 20843 24827 20846
rect 27520 20816 28000 20846
rect 3233 20770 3299 20773
rect 5349 20770 5415 20773
rect 3233 20768 5415 20770
rect 3233 20712 3238 20768
rect 3294 20712 5354 20768
rect 5410 20712 5415 20768
rect 3233 20710 5415 20712
rect 3233 20707 3299 20710
rect 5349 20707 5415 20710
rect 6729 20770 6795 20773
rect 8385 20770 8451 20773
rect 6729 20768 8451 20770
rect 6729 20712 6734 20768
rect 6790 20712 8390 20768
rect 8446 20712 8451 20768
rect 6729 20710 8451 20712
rect 6729 20707 6795 20710
rect 8385 20707 8451 20710
rect 15377 20770 15443 20773
rect 17125 20770 17191 20773
rect 15377 20768 17191 20770
rect 15377 20712 15382 20768
rect 15438 20712 17130 20768
rect 17186 20712 17191 20768
rect 15377 20710 17191 20712
rect 15377 20707 15443 20710
rect 17125 20707 17191 20710
rect 25221 20770 25287 20773
rect 25221 20768 25330 20770
rect 25221 20712 25226 20768
rect 25282 20712 25330 20768
rect 25221 20707 25330 20712
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 6821 20634 6887 20637
rect 10225 20634 10291 20637
rect 6821 20632 10291 20634
rect 6821 20576 6826 20632
rect 6882 20576 10230 20632
rect 10286 20576 10291 20632
rect 6821 20574 10291 20576
rect 6821 20571 6887 20574
rect 10225 20571 10291 20574
rect 17861 20634 17927 20637
rect 19057 20634 19123 20637
rect 19609 20634 19675 20637
rect 17861 20632 19675 20634
rect 17861 20576 17866 20632
rect 17922 20576 19062 20632
rect 19118 20576 19614 20632
rect 19670 20576 19675 20632
rect 17861 20574 19675 20576
rect 17861 20571 17927 20574
rect 19057 20571 19123 20574
rect 19609 20571 19675 20574
rect 3325 20498 3391 20501
rect 9029 20498 9095 20501
rect 3325 20496 9095 20498
rect 3325 20440 3330 20496
rect 3386 20440 9034 20496
rect 9090 20440 9095 20496
rect 3325 20438 9095 20440
rect 3325 20435 3391 20438
rect 9029 20435 9095 20438
rect 9622 20436 9628 20500
rect 9692 20498 9698 20500
rect 11145 20498 11211 20501
rect 9692 20496 11211 20498
rect 9692 20440 11150 20496
rect 11206 20440 11211 20496
rect 9692 20438 11211 20440
rect 9692 20436 9698 20438
rect 11145 20435 11211 20438
rect 11881 20498 11947 20501
rect 17309 20498 17375 20501
rect 24669 20498 24735 20501
rect 11881 20496 24735 20498
rect 11881 20440 11886 20496
rect 11942 20440 17314 20496
rect 17370 20440 24674 20496
rect 24730 20440 24735 20496
rect 11881 20438 24735 20440
rect 11881 20435 11947 20438
rect 17309 20435 17375 20438
rect 24669 20435 24735 20438
rect 0 20362 480 20392
rect 11053 20362 11119 20365
rect 0 20360 11119 20362
rect 0 20304 11058 20360
rect 11114 20304 11119 20360
rect 0 20302 11119 20304
rect 0 20272 480 20302
rect 11053 20299 11119 20302
rect 24117 20362 24183 20365
rect 25270 20362 25330 20707
rect 27520 20362 28000 20392
rect 24117 20360 24410 20362
rect 24117 20304 24122 20360
rect 24178 20304 24410 20360
rect 24117 20302 24410 20304
rect 25270 20302 28000 20362
rect 24117 20299 24183 20302
rect 2313 20226 2379 20229
rect 3325 20226 3391 20229
rect 2313 20224 3391 20226
rect 2313 20168 2318 20224
rect 2374 20168 3330 20224
rect 3386 20168 3391 20224
rect 2313 20166 3391 20168
rect 2313 20163 2379 20166
rect 3325 20163 3391 20166
rect 4797 20226 4863 20229
rect 10041 20226 10107 20229
rect 4797 20224 10107 20226
rect 4797 20168 4802 20224
rect 4858 20168 10046 20224
rect 10102 20168 10107 20224
rect 4797 20166 10107 20168
rect 4797 20163 4863 20166
rect 10041 20163 10107 20166
rect 21817 20226 21883 20229
rect 24117 20226 24183 20229
rect 21817 20224 24183 20226
rect 21817 20168 21822 20224
rect 21878 20168 24122 20224
rect 24178 20168 24183 20224
rect 21817 20166 24183 20168
rect 21817 20163 21883 20166
rect 24117 20163 24183 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1393 20090 1459 20093
rect 4429 20090 4495 20093
rect 1393 20088 4495 20090
rect 1393 20032 1398 20088
rect 1454 20032 4434 20088
rect 4490 20032 4495 20088
rect 1393 20030 4495 20032
rect 1393 20027 1459 20030
rect 4429 20027 4495 20030
rect 6361 20090 6427 20093
rect 8845 20090 8911 20093
rect 6361 20088 8911 20090
rect 6361 20032 6366 20088
rect 6422 20032 8850 20088
rect 8906 20032 8911 20088
rect 6361 20030 8911 20032
rect 6361 20027 6427 20030
rect 8845 20027 8911 20030
rect 10869 20090 10935 20093
rect 15469 20090 15535 20093
rect 10869 20088 15535 20090
rect 10869 20032 10874 20088
rect 10930 20032 15474 20088
rect 15530 20032 15535 20088
rect 10869 20030 15535 20032
rect 10869 20027 10935 20030
rect 15469 20027 15535 20030
rect 20069 20090 20135 20093
rect 24350 20090 24410 20302
rect 27520 20272 28000 20302
rect 25221 20090 25287 20093
rect 20069 20088 25287 20090
rect 20069 20032 20074 20088
rect 20130 20032 25226 20088
rect 25282 20032 25287 20088
rect 20069 20030 25287 20032
rect 20069 20027 20135 20030
rect 25221 20027 25287 20030
rect 4337 19954 4403 19957
rect 13353 19954 13419 19957
rect 21265 19954 21331 19957
rect 4337 19952 13419 19954
rect 4337 19896 4342 19952
rect 4398 19896 13358 19952
rect 13414 19896 13419 19952
rect 4337 19894 13419 19896
rect 4337 19891 4403 19894
rect 13353 19891 13419 19894
rect 16070 19952 21331 19954
rect 16070 19896 21270 19952
rect 21326 19896 21331 19952
rect 16070 19894 21331 19896
rect 1853 19818 1919 19821
rect 3141 19818 3207 19821
rect 1853 19816 3207 19818
rect 1853 19760 1858 19816
rect 1914 19760 3146 19816
rect 3202 19760 3207 19816
rect 1853 19758 3207 19760
rect 1853 19755 1919 19758
rect 3141 19755 3207 19758
rect 10961 19818 11027 19821
rect 16070 19818 16130 19894
rect 21265 19891 21331 19894
rect 10961 19816 16130 19818
rect 10961 19760 10966 19816
rect 11022 19760 16130 19816
rect 10961 19758 16130 19760
rect 16205 19818 16271 19821
rect 25313 19818 25379 19821
rect 16205 19816 25379 19818
rect 16205 19760 16210 19816
rect 16266 19760 25318 19816
rect 25374 19760 25379 19816
rect 16205 19758 25379 19760
rect 10961 19755 11027 19758
rect 16205 19755 16271 19758
rect 25313 19755 25379 19758
rect 0 19682 480 19712
rect 4337 19682 4403 19685
rect 0 19680 4403 19682
rect 0 19624 4342 19680
rect 4398 19624 4403 19680
rect 0 19622 4403 19624
rect 0 19592 480 19622
rect 4337 19619 4403 19622
rect 8017 19682 8083 19685
rect 10041 19682 10107 19685
rect 11145 19684 11211 19685
rect 11094 19682 11100 19684
rect 8017 19680 10107 19682
rect 8017 19624 8022 19680
rect 8078 19624 10046 19680
rect 10102 19624 10107 19680
rect 8017 19622 10107 19624
rect 11054 19622 11100 19682
rect 11164 19680 11211 19684
rect 11206 19624 11211 19680
rect 8017 19619 8083 19622
rect 10041 19619 10107 19622
rect 11094 19620 11100 19622
rect 11164 19620 11211 19624
rect 11145 19619 11211 19620
rect 16389 19682 16455 19685
rect 20805 19682 20871 19685
rect 16389 19680 20871 19682
rect 16389 19624 16394 19680
rect 16450 19624 20810 19680
rect 20866 19624 20871 19680
rect 16389 19622 20871 19624
rect 16389 19619 16455 19622
rect 20805 19619 20871 19622
rect 24669 19682 24735 19685
rect 27520 19682 28000 19712
rect 24669 19680 28000 19682
rect 24669 19624 24674 19680
rect 24730 19624 28000 19680
rect 24669 19622 28000 19624
rect 24669 19619 24735 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 27520 19592 28000 19622
rect 24277 19551 24597 19552
rect 2957 19546 3023 19549
rect 4337 19546 4403 19549
rect 2957 19544 4403 19546
rect 2957 19488 2962 19544
rect 3018 19488 4342 19544
rect 4398 19488 4403 19544
rect 2957 19486 4403 19488
rect 2957 19483 3023 19486
rect 4337 19483 4403 19486
rect 10225 19546 10291 19549
rect 10869 19546 10935 19549
rect 10225 19544 10935 19546
rect 10225 19488 10230 19544
rect 10286 19488 10874 19544
rect 10930 19488 10935 19544
rect 10225 19486 10935 19488
rect 10225 19483 10291 19486
rect 10869 19483 10935 19486
rect 3509 19410 3575 19413
rect 8293 19410 8359 19413
rect 3509 19408 8359 19410
rect 3509 19352 3514 19408
rect 3570 19352 8298 19408
rect 8354 19352 8359 19408
rect 3509 19350 8359 19352
rect 3509 19347 3575 19350
rect 8293 19347 8359 19350
rect 9581 19410 9647 19413
rect 14181 19410 14247 19413
rect 9581 19408 11346 19410
rect 9581 19352 9586 19408
rect 9642 19352 11346 19408
rect 9581 19350 11346 19352
rect 9581 19347 9647 19350
rect 3601 19274 3667 19277
rect 4521 19274 4587 19277
rect 11053 19274 11119 19277
rect 3601 19272 11119 19274
rect 3601 19216 3606 19272
rect 3662 19216 4526 19272
rect 4582 19216 11058 19272
rect 11114 19216 11119 19272
rect 3601 19214 11119 19216
rect 11286 19274 11346 19350
rect 14046 19408 14247 19410
rect 14046 19352 14186 19408
rect 14242 19352 14247 19408
rect 14046 19350 14247 19352
rect 13813 19274 13879 19277
rect 11286 19272 13879 19274
rect 11286 19216 13818 19272
rect 13874 19216 13879 19272
rect 11286 19214 13879 19216
rect 3601 19211 3667 19214
rect 4521 19211 4587 19214
rect 11053 19211 11119 19214
rect 13813 19211 13879 19214
rect 0 19138 480 19168
rect 7097 19138 7163 19141
rect 0 19136 7163 19138
rect 0 19080 7102 19136
rect 7158 19080 7163 19136
rect 0 19078 7163 19080
rect 0 19048 480 19078
rect 7097 19075 7163 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 2037 19002 2103 19005
rect 7833 19002 7899 19005
rect 2037 19000 7899 19002
rect 2037 18944 2042 19000
rect 2098 18944 7838 19000
rect 7894 18944 7899 19000
rect 2037 18942 7899 18944
rect 2037 18939 2103 18942
rect 7833 18939 7899 18942
rect 2957 18866 3023 18869
rect 7281 18866 7347 18869
rect 12249 18866 12315 18869
rect 2957 18864 6056 18866
rect 2957 18808 2962 18864
rect 3018 18808 6056 18864
rect 2957 18806 6056 18808
rect 2957 18803 3023 18806
rect 0 18594 480 18624
rect 5996 18594 6056 18806
rect 7281 18864 12315 18866
rect 7281 18808 7286 18864
rect 7342 18808 12254 18864
rect 12310 18808 12315 18864
rect 7281 18806 12315 18808
rect 7281 18803 7347 18806
rect 12249 18803 12315 18806
rect 14046 18733 14106 19350
rect 14181 19347 14247 19350
rect 21449 19410 21515 19413
rect 21449 19408 24778 19410
rect 21449 19352 21454 19408
rect 21510 19352 24778 19408
rect 21449 19350 24778 19352
rect 21449 19347 21515 19350
rect 14457 19274 14523 19277
rect 23841 19274 23907 19277
rect 14457 19272 23907 19274
rect 14457 19216 14462 19272
rect 14518 19216 23846 19272
rect 23902 19216 23907 19272
rect 14457 19214 23907 19216
rect 14457 19211 14523 19214
rect 23841 19211 23907 19214
rect 24718 19138 24778 19350
rect 27520 19138 28000 19168
rect 24718 19078 28000 19138
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 23606 18940 23612 19004
rect 23676 19002 23682 19004
rect 23933 19002 23999 19005
rect 23676 19000 23999 19002
rect 23676 18944 23938 19000
rect 23994 18944 23999 19000
rect 23676 18942 23999 18944
rect 23676 18940 23682 18942
rect 23933 18939 23999 18942
rect 20897 18866 20963 18869
rect 23933 18866 23999 18869
rect 20897 18864 23999 18866
rect 20897 18808 20902 18864
rect 20958 18808 23938 18864
rect 23994 18808 23999 18864
rect 20897 18806 23999 18808
rect 20897 18803 20963 18806
rect 23933 18803 23999 18806
rect 7833 18730 7899 18733
rect 10133 18730 10199 18733
rect 7833 18728 10199 18730
rect 7833 18672 7838 18728
rect 7894 18672 10138 18728
rect 10194 18672 10199 18728
rect 7833 18670 10199 18672
rect 7833 18667 7899 18670
rect 10133 18667 10199 18670
rect 10501 18730 10567 18733
rect 12801 18730 12867 18733
rect 10501 18728 12867 18730
rect 10501 18672 10506 18728
rect 10562 18672 12806 18728
rect 12862 18672 12867 18728
rect 10501 18670 12867 18672
rect 14046 18728 14155 18733
rect 14046 18672 14094 18728
rect 14150 18672 14155 18728
rect 14046 18670 14155 18672
rect 10501 18667 10567 18670
rect 12801 18667 12867 18670
rect 14089 18667 14155 18670
rect 23749 18730 23815 18733
rect 26233 18730 26299 18733
rect 23749 18728 26299 18730
rect 23749 18672 23754 18728
rect 23810 18672 26238 18728
rect 26294 18672 26299 18728
rect 23749 18670 26299 18672
rect 23749 18667 23815 18670
rect 26233 18667 26299 18670
rect 9305 18594 9371 18597
rect 0 18534 2744 18594
rect 5996 18592 9371 18594
rect 5996 18536 9310 18592
rect 9366 18536 9371 18592
rect 5996 18534 9371 18536
rect 0 18504 480 18534
rect 2684 18458 2744 18534
rect 9305 18531 9371 18534
rect 10317 18594 10383 18597
rect 13813 18594 13879 18597
rect 27520 18594 28000 18624
rect 10317 18592 13879 18594
rect 10317 18536 10322 18592
rect 10378 18536 13818 18592
rect 13874 18536 13879 18592
rect 10317 18534 13879 18536
rect 10317 18531 10383 18534
rect 13813 18531 13879 18534
rect 24902 18534 28000 18594
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 5441 18458 5507 18461
rect 2684 18456 5507 18458
rect 2684 18400 5446 18456
rect 5502 18400 5507 18456
rect 2684 18398 5507 18400
rect 5441 18395 5507 18398
rect 9029 18458 9095 18461
rect 12157 18458 12223 18461
rect 20805 18458 20871 18461
rect 22093 18460 22159 18461
rect 22093 18458 22140 18460
rect 9029 18456 12223 18458
rect 9029 18400 9034 18456
rect 9090 18400 12162 18456
rect 12218 18400 12223 18456
rect 9029 18398 12223 18400
rect 9029 18395 9095 18398
rect 12157 18395 12223 18398
rect 19750 18456 20871 18458
rect 19750 18400 20810 18456
rect 20866 18400 20871 18456
rect 19750 18398 20871 18400
rect 22048 18456 22140 18458
rect 22048 18400 22098 18456
rect 22048 18398 22140 18400
rect 7833 18322 7899 18325
rect 10225 18322 10291 18325
rect 12893 18322 12959 18325
rect 7833 18320 12959 18322
rect 7833 18264 7838 18320
rect 7894 18264 10230 18320
rect 10286 18264 12898 18320
rect 12954 18264 12959 18320
rect 7833 18262 12959 18264
rect 7833 18259 7899 18262
rect 10225 18259 10291 18262
rect 12893 18259 12959 18262
rect 13445 18322 13511 18325
rect 19750 18322 19810 18398
rect 20805 18395 20871 18398
rect 22093 18396 22140 18398
rect 22204 18396 22210 18460
rect 22093 18395 22159 18396
rect 13445 18320 19810 18322
rect 13445 18264 13450 18320
rect 13506 18264 19810 18320
rect 13445 18262 19810 18264
rect 19977 18322 20043 18325
rect 24902 18322 24962 18534
rect 27520 18504 28000 18534
rect 19977 18320 24962 18322
rect 19977 18264 19982 18320
rect 20038 18264 24962 18320
rect 19977 18262 24962 18264
rect 13445 18259 13511 18262
rect 19977 18259 20043 18262
rect 2773 18186 2839 18189
rect 6545 18186 6611 18189
rect 2773 18184 6611 18186
rect 2773 18128 2778 18184
rect 2834 18128 6550 18184
rect 6606 18128 6611 18184
rect 2773 18126 6611 18128
rect 2773 18123 2839 18126
rect 6545 18123 6611 18126
rect 8201 18186 8267 18189
rect 12709 18186 12775 18189
rect 8201 18184 12775 18186
rect 8201 18128 8206 18184
rect 8262 18128 12714 18184
rect 12770 18128 12775 18184
rect 8201 18126 12775 18128
rect 8201 18123 8267 18126
rect 12709 18123 12775 18126
rect 20805 18186 20871 18189
rect 21081 18186 21147 18189
rect 22829 18186 22895 18189
rect 20805 18184 22895 18186
rect 20805 18128 20810 18184
rect 20866 18128 21086 18184
rect 21142 18128 22834 18184
rect 22890 18128 22895 18184
rect 20805 18126 22895 18128
rect 20805 18123 20871 18126
rect 21081 18123 21147 18126
rect 22829 18123 22895 18126
rect 0 18050 480 18080
rect 5809 18050 5875 18053
rect 0 18048 5875 18050
rect 0 17992 5814 18048
rect 5870 17992 5875 18048
rect 0 17990 5875 17992
rect 0 17960 480 17990
rect 5809 17987 5875 17990
rect 12249 18050 12315 18053
rect 19057 18050 19123 18053
rect 19374 18050 19380 18052
rect 12249 18048 19380 18050
rect 12249 17992 12254 18048
rect 12310 17992 19062 18048
rect 19118 17992 19380 18048
rect 12249 17990 19380 17992
rect 12249 17987 12315 17990
rect 19057 17987 19123 17990
rect 19374 17988 19380 17990
rect 19444 17988 19450 18052
rect 27520 18050 28000 18080
rect 23430 17990 28000 18050
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 1945 17914 2011 17917
rect 5533 17914 5599 17917
rect 9397 17914 9463 17917
rect 1945 17912 5599 17914
rect 1945 17856 1950 17912
rect 2006 17856 5538 17912
rect 5594 17856 5599 17912
rect 1945 17854 5599 17856
rect 1945 17851 2011 17854
rect 5533 17851 5599 17854
rect 5766 17912 9463 17914
rect 5766 17856 9402 17912
rect 9458 17856 9463 17912
rect 5766 17854 9463 17856
rect 1485 17778 1551 17781
rect 4245 17778 4311 17781
rect 4889 17778 4955 17781
rect 5766 17778 5826 17854
rect 9397 17851 9463 17854
rect 11605 17914 11671 17917
rect 16757 17914 16823 17917
rect 11605 17912 16823 17914
rect 11605 17856 11610 17912
rect 11666 17856 16762 17912
rect 16818 17856 16823 17912
rect 11605 17854 16823 17856
rect 11605 17851 11671 17854
rect 16757 17851 16823 17854
rect 22645 17914 22711 17917
rect 23430 17914 23490 17990
rect 27520 17960 28000 17990
rect 22645 17912 23490 17914
rect 22645 17856 22650 17912
rect 22706 17856 23490 17912
rect 22645 17854 23490 17856
rect 22645 17851 22711 17854
rect 1485 17776 1778 17778
rect 1485 17720 1490 17776
rect 1546 17720 1778 17776
rect 1485 17718 1778 17720
rect 1485 17715 1551 17718
rect 0 17506 480 17536
rect 1577 17506 1643 17509
rect 0 17504 1643 17506
rect 0 17448 1582 17504
rect 1638 17448 1643 17504
rect 0 17446 1643 17448
rect 0 17416 480 17446
rect 1577 17443 1643 17446
rect 1718 16962 1778 17718
rect 4245 17776 5826 17778
rect 4245 17720 4250 17776
rect 4306 17720 4894 17776
rect 4950 17720 5826 17776
rect 4245 17718 5826 17720
rect 6177 17778 6243 17781
rect 9029 17778 9095 17781
rect 6177 17776 9095 17778
rect 6177 17720 6182 17776
rect 6238 17720 9034 17776
rect 9090 17720 9095 17776
rect 6177 17718 9095 17720
rect 4245 17715 4311 17718
rect 4889 17715 4955 17718
rect 6177 17715 6243 17718
rect 9029 17715 9095 17718
rect 9489 17778 9555 17781
rect 13353 17778 13419 17781
rect 19333 17778 19399 17781
rect 9489 17776 13419 17778
rect 9489 17720 9494 17776
rect 9550 17720 13358 17776
rect 13414 17720 13419 17776
rect 9489 17718 13419 17720
rect 9489 17715 9555 17718
rect 13353 17715 13419 17718
rect 13678 17776 19399 17778
rect 13678 17720 19338 17776
rect 19394 17720 19399 17776
rect 13678 17718 19399 17720
rect 8385 17644 8451 17645
rect 8334 17580 8340 17644
rect 8404 17642 8451 17644
rect 9673 17642 9739 17645
rect 13678 17642 13738 17718
rect 19333 17715 19399 17718
rect 15377 17642 15443 17645
rect 8404 17640 8496 17642
rect 8446 17584 8496 17640
rect 8404 17582 8496 17584
rect 9673 17640 13738 17642
rect 9673 17584 9678 17640
rect 9734 17584 13738 17640
rect 9673 17582 13738 17584
rect 13862 17640 15443 17642
rect 13862 17584 15382 17640
rect 15438 17584 15443 17640
rect 13862 17582 15443 17584
rect 8404 17580 8451 17582
rect 8385 17579 8451 17580
rect 9673 17579 9739 17582
rect 7373 17506 7439 17509
rect 13862 17506 13922 17582
rect 15377 17579 15443 17582
rect 7373 17504 13922 17506
rect 7373 17448 7378 17504
rect 7434 17448 13922 17504
rect 7373 17446 13922 17448
rect 16757 17506 16823 17509
rect 20897 17506 20963 17509
rect 16757 17504 20963 17506
rect 16757 17448 16762 17504
rect 16818 17448 20902 17504
rect 20958 17448 20963 17504
rect 16757 17446 20963 17448
rect 7373 17443 7439 17446
rect 16757 17443 16823 17446
rect 20897 17443 20963 17446
rect 24761 17506 24827 17509
rect 27520 17506 28000 17536
rect 24761 17504 28000 17506
rect 24761 17448 24766 17504
rect 24822 17448 28000 17504
rect 24761 17446 28000 17448
rect 24761 17443 24827 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17446
rect 24277 17375 24597 17376
rect 8017 17370 8083 17373
rect 11053 17370 11119 17373
rect 8017 17368 11119 17370
rect 8017 17312 8022 17368
rect 8078 17312 11058 17368
rect 11114 17312 11119 17368
rect 8017 17310 11119 17312
rect 8017 17307 8083 17310
rect 11053 17307 11119 17310
rect 11329 17370 11395 17373
rect 13169 17370 13235 17373
rect 11329 17368 13235 17370
rect 11329 17312 11334 17368
rect 11390 17312 13174 17368
rect 13230 17312 13235 17368
rect 11329 17310 13235 17312
rect 11329 17307 11395 17310
rect 13169 17307 13235 17310
rect 18505 17370 18571 17373
rect 23841 17370 23907 17373
rect 18505 17368 23907 17370
rect 18505 17312 18510 17368
rect 18566 17312 23846 17368
rect 23902 17312 23907 17368
rect 18505 17310 23907 17312
rect 18505 17307 18571 17310
rect 23841 17307 23907 17310
rect 5533 17234 5599 17237
rect 9397 17234 9463 17237
rect 5533 17232 9463 17234
rect 5533 17176 5538 17232
rect 5594 17176 9402 17232
rect 9458 17176 9463 17232
rect 5533 17174 9463 17176
rect 5533 17171 5599 17174
rect 9397 17171 9463 17174
rect 12433 17234 12499 17237
rect 21633 17234 21699 17237
rect 12433 17232 21699 17234
rect 12433 17176 12438 17232
rect 12494 17176 21638 17232
rect 21694 17176 21699 17232
rect 12433 17174 21699 17176
rect 12433 17171 12499 17174
rect 21633 17171 21699 17174
rect 5349 17098 5415 17101
rect 7557 17098 7623 17101
rect 5349 17096 7623 17098
rect 5349 17040 5354 17096
rect 5410 17040 7562 17096
rect 7618 17040 7623 17096
rect 5349 17038 7623 17040
rect 5349 17035 5415 17038
rect 7557 17035 7623 17038
rect 8385 17098 8451 17101
rect 15285 17098 15351 17101
rect 8385 17096 15351 17098
rect 8385 17040 8390 17096
rect 8446 17040 15290 17096
rect 15346 17040 15351 17096
rect 8385 17038 15351 17040
rect 8385 17035 8451 17038
rect 15285 17035 15351 17038
rect 18689 17098 18755 17101
rect 24393 17098 24459 17101
rect 18689 17096 24459 17098
rect 18689 17040 18694 17096
rect 18750 17040 24398 17096
rect 24454 17040 24459 17096
rect 18689 17038 24459 17040
rect 18689 17035 18755 17038
rect 24393 17035 24459 17038
rect 7373 16962 7439 16965
rect 1718 16960 7439 16962
rect 1718 16904 7378 16960
rect 7434 16904 7439 16960
rect 1718 16902 7439 16904
rect 7373 16899 7439 16902
rect 7833 16962 7899 16965
rect 9673 16962 9739 16965
rect 7833 16960 9739 16962
rect 7833 16904 7838 16960
rect 7894 16904 9678 16960
rect 9734 16904 9739 16960
rect 7833 16902 9739 16904
rect 7833 16899 7899 16902
rect 9673 16899 9739 16902
rect 10777 16962 10843 16965
rect 18505 16962 18571 16965
rect 19241 16962 19307 16965
rect 10777 16960 19307 16962
rect 10777 16904 10782 16960
rect 10838 16904 18510 16960
rect 18566 16904 19246 16960
rect 19302 16904 19307 16960
rect 10777 16902 19307 16904
rect 10777 16899 10843 16902
rect 18505 16899 18571 16902
rect 19241 16899 19307 16902
rect 23289 16962 23355 16965
rect 23749 16962 23815 16965
rect 25037 16962 25103 16965
rect 23289 16960 25103 16962
rect 23289 16904 23294 16960
rect 23350 16904 23754 16960
rect 23810 16904 25042 16960
rect 25098 16904 25103 16960
rect 23289 16902 25103 16904
rect 23289 16899 23355 16902
rect 23749 16899 23815 16902
rect 25037 16899 25103 16902
rect 10277 16896 10597 16897
rect 0 16826 480 16856
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 4245 16826 4311 16829
rect 0 16824 4311 16826
rect 0 16768 4250 16824
rect 4306 16768 4311 16824
rect 0 16766 4311 16768
rect 0 16736 480 16766
rect 4245 16763 4311 16766
rect 11421 16826 11487 16829
rect 18689 16826 18755 16829
rect 11421 16824 18755 16826
rect 11421 16768 11426 16824
rect 11482 16768 18694 16824
rect 18750 16768 18755 16824
rect 11421 16766 18755 16768
rect 11421 16763 11487 16766
rect 18689 16763 18755 16766
rect 25129 16826 25195 16829
rect 27520 16826 28000 16856
rect 25129 16824 28000 16826
rect 25129 16768 25134 16824
rect 25190 16768 28000 16824
rect 25129 16766 28000 16768
rect 25129 16763 25195 16766
rect 27520 16736 28000 16766
rect 7189 16688 7255 16693
rect 7189 16632 7194 16688
rect 7250 16632 7255 16688
rect 7189 16627 7255 16632
rect 8017 16690 8083 16693
rect 14365 16690 14431 16693
rect 8017 16688 14431 16690
rect 8017 16632 8022 16688
rect 8078 16632 14370 16688
rect 14426 16632 14431 16688
rect 8017 16630 14431 16632
rect 8017 16627 8083 16630
rect 14365 16627 14431 16630
rect 15101 16690 15167 16693
rect 15837 16690 15903 16693
rect 18045 16690 18111 16693
rect 15101 16688 18111 16690
rect 15101 16632 15106 16688
rect 15162 16632 15842 16688
rect 15898 16632 18050 16688
rect 18106 16632 18111 16688
rect 15101 16630 18111 16632
rect 15101 16627 15167 16630
rect 15837 16627 15903 16630
rect 18045 16627 18111 16630
rect 18873 16690 18939 16693
rect 21265 16690 21331 16693
rect 18873 16688 21331 16690
rect 18873 16632 18878 16688
rect 18934 16632 21270 16688
rect 21326 16632 21331 16688
rect 18873 16630 21331 16632
rect 18873 16627 18939 16630
rect 21265 16627 21331 16630
rect 2405 16554 2471 16557
rect 7192 16554 7252 16627
rect 23422 16554 23428 16556
rect 2405 16552 7114 16554
rect 2405 16496 2410 16552
rect 2466 16496 7114 16552
rect 2405 16494 7114 16496
rect 7192 16494 23428 16554
rect 2405 16491 2471 16494
rect 5610 16352 5930 16353
rect 0 16282 480 16312
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 2221 16282 2287 16285
rect 0 16280 2287 16282
rect 0 16224 2226 16280
rect 2282 16224 2287 16280
rect 0 16222 2287 16224
rect 7054 16282 7114 16494
rect 23422 16492 23428 16494
rect 23492 16492 23498 16556
rect 8845 16418 8911 16421
rect 13813 16418 13879 16421
rect 14181 16418 14247 16421
rect 8845 16416 14247 16418
rect 8845 16360 8850 16416
rect 8906 16360 13818 16416
rect 13874 16360 14186 16416
rect 14242 16360 14247 16416
rect 8845 16358 14247 16360
rect 8845 16355 8911 16358
rect 13813 16355 13879 16358
rect 14181 16355 14247 16358
rect 22369 16418 22435 16421
rect 24117 16418 24183 16421
rect 22369 16416 24183 16418
rect 22369 16360 22374 16416
rect 22430 16360 24122 16416
rect 24178 16360 24183 16416
rect 22369 16358 24183 16360
rect 22369 16355 22435 16358
rect 24117 16355 24183 16358
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 10869 16282 10935 16285
rect 7054 16280 10935 16282
rect 7054 16224 10874 16280
rect 10930 16224 10935 16280
rect 7054 16222 10935 16224
rect 0 16192 480 16222
rect 2221 16219 2287 16222
rect 10869 16219 10935 16222
rect 11145 16282 11211 16285
rect 12525 16282 12591 16285
rect 13629 16282 13695 16285
rect 11145 16280 13695 16282
rect 11145 16224 11150 16280
rect 11206 16224 12530 16280
rect 12586 16224 13634 16280
rect 13690 16224 13695 16280
rect 11145 16222 13695 16224
rect 11145 16219 11211 16222
rect 12525 16219 12591 16222
rect 13629 16219 13695 16222
rect 25497 16282 25563 16285
rect 27520 16282 28000 16312
rect 25497 16280 28000 16282
rect 25497 16224 25502 16280
rect 25558 16224 28000 16280
rect 25497 16222 28000 16224
rect 25497 16219 25563 16222
rect 27520 16192 28000 16222
rect 5441 16146 5507 16149
rect 8293 16146 8359 16149
rect 8477 16146 8543 16149
rect 5441 16144 8543 16146
rect 5441 16088 5446 16144
rect 5502 16088 8298 16144
rect 8354 16088 8482 16144
rect 8538 16088 8543 16144
rect 5441 16086 8543 16088
rect 5441 16083 5507 16086
rect 8293 16083 8359 16086
rect 8477 16083 8543 16086
rect 9673 16146 9739 16149
rect 14641 16146 14707 16149
rect 16113 16146 16179 16149
rect 9673 16144 14060 16146
rect 9673 16088 9678 16144
rect 9734 16088 14060 16144
rect 9673 16086 14060 16088
rect 9673 16083 9739 16086
rect 8569 16010 8635 16013
rect 11329 16010 11395 16013
rect 13813 16010 13879 16013
rect 7468 16008 10748 16010
rect 7468 15952 8574 16008
rect 8630 15952 10748 16008
rect 7468 15950 10748 15952
rect 4981 15874 5047 15877
rect 7468 15874 7528 15950
rect 8569 15947 8635 15950
rect 4981 15872 7528 15874
rect 4981 15816 4986 15872
rect 5042 15816 7528 15872
rect 4981 15814 7528 15816
rect 10688 15874 10748 15950
rect 11329 16008 13879 16010
rect 11329 15952 11334 16008
rect 11390 15952 13818 16008
rect 13874 15952 13879 16008
rect 11329 15950 13879 15952
rect 14000 16010 14060 16086
rect 14641 16144 16179 16146
rect 14641 16088 14646 16144
rect 14702 16088 16118 16144
rect 16174 16088 16179 16144
rect 14641 16086 16179 16088
rect 14641 16083 14707 16086
rect 16113 16083 16179 16086
rect 19333 16010 19399 16013
rect 14000 16008 19399 16010
rect 14000 15952 19338 16008
rect 19394 15952 19399 16008
rect 14000 15950 19399 15952
rect 11329 15947 11395 15950
rect 13813 15947 13879 15950
rect 19333 15947 19399 15950
rect 17677 15874 17743 15877
rect 10688 15872 17743 15874
rect 10688 15816 17682 15872
rect 17738 15816 17743 15872
rect 10688 15814 17743 15816
rect 4981 15811 5047 15814
rect 17677 15811 17743 15814
rect 10277 15808 10597 15809
rect 0 15738 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 1577 15738 1643 15741
rect 0 15736 1643 15738
rect 0 15680 1582 15736
rect 1638 15680 1643 15736
rect 0 15678 1643 15680
rect 0 15648 480 15678
rect 1577 15675 1643 15678
rect 3325 15738 3391 15741
rect 7833 15738 7899 15741
rect 3325 15736 7899 15738
rect 3325 15680 3330 15736
rect 3386 15680 7838 15736
rect 7894 15680 7899 15736
rect 3325 15678 7899 15680
rect 3325 15675 3391 15678
rect 7833 15675 7899 15678
rect 13721 15738 13787 15741
rect 18137 15738 18203 15741
rect 13721 15736 18203 15738
rect 13721 15680 13726 15736
rect 13782 15680 18142 15736
rect 18198 15680 18203 15736
rect 13721 15678 18203 15680
rect 13721 15675 13787 15678
rect 18137 15675 18203 15678
rect 24117 15738 24183 15741
rect 27520 15738 28000 15768
rect 24117 15736 28000 15738
rect 24117 15680 24122 15736
rect 24178 15680 28000 15736
rect 24117 15678 28000 15680
rect 24117 15675 24183 15678
rect 27520 15648 28000 15678
rect 3693 15602 3759 15605
rect 8017 15602 8083 15605
rect 3693 15600 8083 15602
rect 3693 15544 3698 15600
rect 3754 15544 8022 15600
rect 8078 15544 8083 15600
rect 3693 15542 8083 15544
rect 3693 15539 3759 15542
rect 8017 15539 8083 15542
rect 20897 15602 20963 15605
rect 23974 15602 23980 15604
rect 20897 15600 23980 15602
rect 20897 15544 20902 15600
rect 20958 15544 23980 15600
rect 20897 15542 23980 15544
rect 20897 15539 20963 15542
rect 23974 15540 23980 15542
rect 24044 15540 24050 15604
rect 289 15466 355 15469
rect 3877 15466 3943 15469
rect 6177 15466 6243 15469
rect 7005 15466 7071 15469
rect 289 15464 674 15466
rect 289 15408 294 15464
rect 350 15408 674 15464
rect 289 15406 674 15408
rect 289 15403 355 15406
rect 614 15330 674 15406
rect 3877 15464 7071 15466
rect 3877 15408 3882 15464
rect 3938 15408 6182 15464
rect 6238 15408 7010 15464
rect 7066 15408 7071 15464
rect 3877 15406 7071 15408
rect 3877 15403 3943 15406
rect 6177 15403 6243 15406
rect 7005 15403 7071 15406
rect 7465 15466 7531 15469
rect 10317 15466 10383 15469
rect 7465 15464 10383 15466
rect 7465 15408 7470 15464
rect 7526 15408 10322 15464
rect 10378 15408 10383 15464
rect 7465 15406 10383 15408
rect 7465 15403 7531 15406
rect 10317 15403 10383 15406
rect 14089 15466 14155 15469
rect 24945 15466 25011 15469
rect 14089 15464 25011 15466
rect 14089 15408 14094 15464
rect 14150 15408 24950 15464
rect 25006 15408 25011 15464
rect 14089 15406 25011 15408
rect 14089 15403 14155 15406
rect 24945 15403 25011 15406
rect 5349 15330 5415 15333
rect 614 15328 5415 15330
rect 614 15272 5354 15328
rect 5410 15272 5415 15328
rect 614 15270 5415 15272
rect 5349 15267 5415 15270
rect 7465 15330 7531 15333
rect 11145 15330 11211 15333
rect 7465 15328 11211 15330
rect 7465 15272 7470 15328
rect 7526 15272 11150 15328
rect 11206 15272 11211 15328
rect 7465 15270 11211 15272
rect 7465 15267 7531 15270
rect 11145 15267 11211 15270
rect 15653 15330 15719 15333
rect 16849 15330 16915 15333
rect 23381 15330 23447 15333
rect 15653 15328 23447 15330
rect 15653 15272 15658 15328
rect 15714 15272 16854 15328
rect 16910 15272 23386 15328
rect 23442 15272 23447 15328
rect 15653 15270 23447 15272
rect 15653 15267 15719 15270
rect 16849 15267 16915 15270
rect 23381 15267 23447 15270
rect 5610 15264 5930 15265
rect 0 15194 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 2681 15194 2747 15197
rect 0 15192 2747 15194
rect 0 15136 2686 15192
rect 2742 15136 2747 15192
rect 0 15134 2747 15136
rect 0 15104 480 15134
rect 2681 15131 2747 15134
rect 10777 15194 10843 15197
rect 13353 15194 13419 15197
rect 10777 15192 13419 15194
rect 10777 15136 10782 15192
rect 10838 15136 13358 15192
rect 13414 15136 13419 15192
rect 10777 15134 13419 15136
rect 10777 15131 10843 15134
rect 13353 15131 13419 15134
rect 14365 15194 14431 15197
rect 27520 15194 28000 15224
rect 14365 15192 14842 15194
rect 14365 15136 14370 15192
rect 14426 15136 14842 15192
rect 14365 15134 14842 15136
rect 14365 15131 14431 15134
rect 2497 15058 2563 15061
rect 11605 15058 11671 15061
rect 2497 15056 11671 15058
rect 2497 15000 2502 15056
rect 2558 15000 11610 15056
rect 11666 15000 11671 15056
rect 2497 14998 11671 15000
rect 14782 15058 14842 15134
rect 24672 15134 28000 15194
rect 21265 15058 21331 15061
rect 14782 15056 21331 15058
rect 14782 15000 21270 15056
rect 21326 15000 21331 15056
rect 14782 14998 21331 15000
rect 2497 14995 2563 14998
rect 11605 14995 11671 14998
rect 21265 14995 21331 14998
rect 22001 15058 22067 15061
rect 24672 15058 24732 15134
rect 27520 15104 28000 15134
rect 22001 15056 24732 15058
rect 22001 15000 22006 15056
rect 22062 15000 24732 15056
rect 22001 14998 24732 15000
rect 22001 14995 22067 14998
rect 6729 14922 6795 14925
rect 18045 14922 18111 14925
rect 6729 14920 18111 14922
rect 6729 14864 6734 14920
rect 6790 14864 18050 14920
rect 18106 14864 18111 14920
rect 6729 14862 18111 14864
rect 6729 14859 6795 14862
rect 18045 14859 18111 14862
rect 22134 14860 22140 14924
rect 22204 14922 22210 14924
rect 22645 14922 22711 14925
rect 22204 14920 22711 14922
rect 22204 14864 22650 14920
rect 22706 14864 22711 14920
rect 22204 14862 22711 14864
rect 22204 14860 22210 14862
rect 22645 14859 22711 14862
rect 3233 14786 3299 14789
rect 10133 14786 10199 14789
rect 3233 14784 10199 14786
rect 3233 14728 3238 14784
rect 3294 14728 10138 14784
rect 10194 14728 10199 14784
rect 3233 14726 10199 14728
rect 3233 14723 3299 14726
rect 10133 14723 10199 14726
rect 12341 14786 12407 14789
rect 14457 14786 14523 14789
rect 12341 14784 14523 14786
rect 12341 14728 12346 14784
rect 12402 14728 14462 14784
rect 14518 14728 14523 14784
rect 12341 14726 14523 14728
rect 12341 14723 12407 14726
rect 14457 14723 14523 14726
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1577 14650 1643 14653
rect 0 14648 1643 14650
rect 0 14592 1582 14648
rect 1638 14592 1643 14648
rect 0 14590 1643 14592
rect 0 14560 480 14590
rect 1577 14587 1643 14590
rect 4061 14650 4127 14653
rect 6269 14650 6335 14653
rect 4061 14648 6335 14650
rect 4061 14592 4066 14648
rect 4122 14592 6274 14648
rect 6330 14592 6335 14648
rect 4061 14590 6335 14592
rect 4061 14587 4127 14590
rect 6269 14587 6335 14590
rect 24209 14650 24275 14653
rect 27520 14650 28000 14680
rect 24209 14648 28000 14650
rect 24209 14592 24214 14648
rect 24270 14592 28000 14648
rect 24209 14590 28000 14592
rect 24209 14587 24275 14590
rect 27520 14560 28000 14590
rect 14457 14514 14523 14517
rect 23933 14514 23999 14517
rect 14457 14512 23999 14514
rect 14457 14456 14462 14512
rect 14518 14456 23938 14512
rect 23994 14456 23999 14512
rect 14457 14454 23999 14456
rect 14457 14451 14523 14454
rect 23933 14451 23999 14454
rect 5533 14378 5599 14381
rect 7833 14378 7899 14381
rect 19241 14378 19307 14381
rect 22277 14378 22343 14381
rect 5533 14376 7899 14378
rect 5533 14320 5538 14376
rect 5594 14320 7838 14376
rect 7894 14320 7899 14376
rect 5533 14318 7899 14320
rect 5533 14315 5599 14318
rect 7833 14315 7899 14318
rect 14782 14318 19074 14378
rect 11145 14242 11211 14245
rect 14641 14242 14707 14245
rect 14782 14242 14842 14318
rect 11145 14240 14842 14242
rect 11145 14184 11150 14240
rect 11206 14184 14646 14240
rect 14702 14184 14842 14240
rect 11145 14182 14842 14184
rect 19014 14242 19074 14318
rect 19241 14376 22343 14378
rect 19241 14320 19246 14376
rect 19302 14320 22282 14376
rect 22338 14320 22343 14376
rect 19241 14318 22343 14320
rect 19241 14315 19307 14318
rect 22277 14315 22343 14318
rect 24301 14378 24367 14381
rect 24710 14378 24716 14380
rect 24301 14376 24716 14378
rect 24301 14320 24306 14376
rect 24362 14320 24716 14376
rect 24301 14318 24716 14320
rect 24301 14315 24367 14318
rect 24710 14316 24716 14318
rect 24780 14316 24786 14380
rect 19425 14242 19491 14245
rect 19701 14242 19767 14245
rect 19014 14240 19767 14242
rect 19014 14184 19430 14240
rect 19486 14184 19706 14240
rect 19762 14184 19767 14240
rect 19014 14182 19767 14184
rect 11145 14179 11211 14182
rect 14641 14179 14707 14182
rect 19425 14179 19491 14182
rect 19701 14179 19767 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 8109 14106 8175 14109
rect 13353 14106 13419 14109
rect 8109 14104 13419 14106
rect 8109 14048 8114 14104
rect 8170 14048 13358 14104
rect 13414 14048 13419 14104
rect 8109 14046 13419 14048
rect 8109 14043 8175 14046
rect 13353 14043 13419 14046
rect 0 13970 480 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 0 13880 480 13910
rect 1485 13907 1551 13910
rect 5349 13970 5415 13973
rect 12985 13970 13051 13973
rect 5349 13968 13051 13970
rect 5349 13912 5354 13968
rect 5410 13912 12990 13968
rect 13046 13912 13051 13968
rect 5349 13910 13051 13912
rect 5349 13907 5415 13910
rect 12985 13907 13051 13910
rect 13169 13970 13235 13973
rect 19333 13970 19399 13973
rect 13169 13968 19399 13970
rect 13169 13912 13174 13968
rect 13230 13912 19338 13968
rect 19394 13912 19399 13968
rect 13169 13910 19399 13912
rect 13169 13907 13235 13910
rect 19333 13907 19399 13910
rect 20989 13970 21055 13973
rect 22829 13970 22895 13973
rect 20989 13968 22895 13970
rect 20989 13912 20994 13968
rect 21050 13912 22834 13968
rect 22890 13912 22895 13968
rect 20989 13910 22895 13912
rect 20989 13907 21055 13910
rect 22829 13907 22895 13910
rect 24761 13970 24827 13973
rect 27520 13970 28000 14000
rect 24761 13968 28000 13970
rect 24761 13912 24766 13968
rect 24822 13912 28000 13968
rect 24761 13910 28000 13912
rect 24761 13907 24827 13910
rect 27520 13880 28000 13910
rect 9305 13834 9371 13837
rect 12157 13834 12223 13837
rect 9305 13832 12223 13834
rect 9305 13776 9310 13832
rect 9366 13776 12162 13832
rect 12218 13776 12223 13832
rect 9305 13774 12223 13776
rect 9305 13771 9371 13774
rect 12157 13771 12223 13774
rect 13537 13834 13603 13837
rect 15377 13834 15443 13837
rect 13537 13832 15443 13834
rect 13537 13776 13542 13832
rect 13598 13776 15382 13832
rect 15438 13776 15443 13832
rect 13537 13774 15443 13776
rect 13537 13771 13603 13774
rect 15377 13771 15443 13774
rect 21909 13834 21975 13837
rect 24301 13834 24367 13837
rect 21909 13832 24367 13834
rect 21909 13776 21914 13832
rect 21970 13776 24306 13832
rect 24362 13776 24367 13832
rect 21909 13774 24367 13776
rect 21909 13771 21975 13774
rect 24301 13771 24367 13774
rect 3693 13698 3759 13701
rect 7833 13698 7899 13701
rect 3693 13696 7899 13698
rect 3693 13640 3698 13696
rect 3754 13640 7838 13696
rect 7894 13640 7899 13696
rect 3693 13638 7899 13640
rect 3693 13635 3759 13638
rect 7833 13635 7899 13638
rect 22829 13698 22895 13701
rect 24117 13698 24183 13701
rect 22829 13696 24183 13698
rect 22829 13640 22834 13696
rect 22890 13640 24122 13696
rect 24178 13640 24183 13696
rect 22829 13638 24183 13640
rect 22829 13635 22895 13638
rect 24117 13635 24183 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3049 13562 3115 13565
rect 3325 13562 3391 13565
rect 8477 13562 8543 13565
rect 3049 13560 3250 13562
rect 3049 13504 3054 13560
rect 3110 13504 3250 13560
rect 3049 13502 3250 13504
rect 3049 13499 3115 13502
rect 0 13426 480 13456
rect 1577 13426 1643 13429
rect 0 13424 1643 13426
rect 0 13368 1582 13424
rect 1638 13368 1643 13424
rect 0 13366 1643 13368
rect 0 13336 480 13366
rect 1577 13363 1643 13366
rect 3190 13290 3250 13502
rect 3325 13560 8543 13562
rect 3325 13504 3330 13560
rect 3386 13504 8482 13560
rect 8538 13504 8543 13560
rect 3325 13502 8543 13504
rect 3325 13499 3391 13502
rect 8477 13499 8543 13502
rect 22553 13562 22619 13565
rect 23749 13562 23815 13565
rect 22553 13560 23815 13562
rect 22553 13504 22558 13560
rect 22614 13504 23754 13560
rect 23810 13504 23815 13560
rect 22553 13502 23815 13504
rect 22553 13499 22619 13502
rect 23749 13499 23815 13502
rect 9121 13426 9187 13429
rect 13997 13426 14063 13429
rect 9121 13424 14063 13426
rect 9121 13368 9126 13424
rect 9182 13368 14002 13424
rect 14058 13368 14063 13424
rect 9121 13366 14063 13368
rect 9121 13363 9187 13366
rect 13997 13363 14063 13366
rect 14181 13426 14247 13429
rect 18597 13426 18663 13429
rect 21265 13426 21331 13429
rect 27520 13426 28000 13456
rect 14181 13424 19258 13426
rect 14181 13368 14186 13424
rect 14242 13368 18602 13424
rect 18658 13368 19258 13424
rect 14181 13366 19258 13368
rect 14181 13363 14247 13366
rect 18597 13363 18663 13366
rect 13445 13290 13511 13293
rect 3190 13288 13511 13290
rect 3190 13232 13450 13288
rect 13506 13232 13511 13288
rect 3190 13230 13511 13232
rect 13445 13227 13511 13230
rect 13721 13290 13787 13293
rect 19057 13290 19123 13293
rect 13721 13288 19123 13290
rect 13721 13232 13726 13288
rect 13782 13232 19062 13288
rect 19118 13232 19123 13288
rect 13721 13230 19123 13232
rect 19198 13290 19258 13366
rect 21265 13424 28000 13426
rect 21265 13368 21270 13424
rect 21326 13368 28000 13424
rect 21265 13366 28000 13368
rect 21265 13363 21331 13366
rect 27520 13336 28000 13366
rect 25589 13290 25655 13293
rect 19198 13288 25655 13290
rect 19198 13232 25594 13288
rect 25650 13232 25655 13288
rect 19198 13230 25655 13232
rect 13721 13227 13787 13230
rect 19057 13227 19123 13230
rect 25589 13227 25655 13230
rect 8845 13154 8911 13157
rect 16297 13154 16363 13157
rect 18045 13154 18111 13157
rect 8845 13152 13922 13154
rect 8845 13096 8850 13152
rect 8906 13096 13922 13152
rect 8845 13094 13922 13096
rect 8845 13091 8911 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 0 12882 480 12912
rect 1577 12882 1643 12885
rect 0 12880 1643 12882
rect 0 12824 1582 12880
rect 1638 12824 1643 12880
rect 0 12822 1643 12824
rect 0 12792 480 12822
rect 1577 12819 1643 12822
rect 3141 12882 3207 12885
rect 5625 12882 5691 12885
rect 3141 12880 5691 12882
rect 3141 12824 3146 12880
rect 3202 12824 5630 12880
rect 5686 12824 5691 12880
rect 3141 12822 5691 12824
rect 3141 12819 3207 12822
rect 5625 12819 5691 12822
rect 8385 12882 8451 12885
rect 13537 12882 13603 12885
rect 8385 12880 13603 12882
rect 8385 12824 8390 12880
rect 8446 12824 13542 12880
rect 13598 12824 13603 12880
rect 8385 12822 13603 12824
rect 8385 12819 8451 12822
rect 13537 12819 13603 12822
rect 3049 12746 3115 12749
rect 7005 12746 7071 12749
rect 7281 12746 7347 12749
rect 3049 12744 7347 12746
rect 3049 12688 3054 12744
rect 3110 12688 7010 12744
rect 7066 12688 7286 12744
rect 7342 12688 7347 12744
rect 3049 12686 7347 12688
rect 3049 12683 3115 12686
rect 7005 12683 7071 12686
rect 7281 12683 7347 12686
rect 9397 12746 9463 12749
rect 12433 12746 12499 12749
rect 9397 12744 12499 12746
rect 9397 12688 9402 12744
rect 9458 12688 12438 12744
rect 12494 12688 12499 12744
rect 9397 12686 12499 12688
rect 13862 12746 13922 13094
rect 16297 13152 18111 13154
rect 16297 13096 16302 13152
rect 16358 13096 18050 13152
rect 18106 13096 18111 13152
rect 16297 13094 18111 13096
rect 16297 13091 16363 13094
rect 18045 13091 18111 13094
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 22553 13018 22619 13021
rect 23473 13020 23539 13021
rect 15334 13016 22619 13018
rect 15334 12960 22558 13016
rect 22614 12960 22619 13016
rect 15334 12958 22619 12960
rect 13997 12882 14063 12885
rect 15334 12882 15394 12958
rect 22553 12955 22619 12958
rect 23422 12956 23428 13020
rect 23492 13018 23539 13020
rect 23492 13016 23584 13018
rect 23534 12960 23584 13016
rect 23492 12958 23584 12960
rect 23492 12956 23539 12958
rect 23473 12955 23539 12956
rect 13997 12880 15394 12882
rect 13997 12824 14002 12880
rect 14058 12824 15394 12880
rect 13997 12822 15394 12824
rect 20345 12882 20411 12885
rect 24945 12882 25011 12885
rect 20345 12880 25011 12882
rect 20345 12824 20350 12880
rect 20406 12824 24950 12880
rect 25006 12824 25011 12880
rect 20345 12822 25011 12824
rect 13997 12819 14063 12822
rect 20345 12819 20411 12822
rect 24945 12819 25011 12822
rect 25405 12882 25471 12885
rect 27520 12882 28000 12912
rect 25405 12880 28000 12882
rect 25405 12824 25410 12880
rect 25466 12824 28000 12880
rect 25405 12822 28000 12824
rect 25405 12819 25471 12822
rect 27520 12792 28000 12822
rect 15377 12746 15443 12749
rect 25313 12746 25379 12749
rect 13862 12744 15443 12746
rect 13862 12688 15382 12744
rect 15438 12688 15443 12744
rect 13862 12686 15443 12688
rect 9397 12683 9463 12686
rect 12433 12683 12499 12686
rect 15377 12683 15443 12686
rect 19198 12744 25379 12746
rect 19198 12688 25318 12744
rect 25374 12688 25379 12744
rect 19198 12686 25379 12688
rect 2129 12610 2195 12613
rect 9029 12610 9095 12613
rect 2129 12608 9095 12610
rect 2129 12552 2134 12608
rect 2190 12552 9034 12608
rect 9090 12552 9095 12608
rect 2129 12550 9095 12552
rect 2129 12547 2195 12550
rect 9029 12547 9095 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 0 12338 480 12368
rect 2681 12338 2747 12341
rect 0 12336 2747 12338
rect 0 12280 2686 12336
rect 2742 12280 2747 12336
rect 0 12278 2747 12280
rect 0 12248 480 12278
rect 2681 12275 2747 12278
rect 7373 12338 7439 12341
rect 8334 12338 8340 12340
rect 7373 12336 8340 12338
rect 7373 12280 7378 12336
rect 7434 12280 8340 12336
rect 7373 12278 8340 12280
rect 7373 12275 7439 12278
rect 8334 12276 8340 12278
rect 8404 12276 8410 12340
rect 10777 12338 10843 12341
rect 19198 12338 19258 12686
rect 25313 12683 25379 12686
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 10777 12336 19258 12338
rect 10777 12280 10782 12336
rect 10838 12280 19258 12336
rect 10777 12278 19258 12280
rect 25405 12338 25471 12341
rect 27520 12338 28000 12368
rect 25405 12336 28000 12338
rect 25405 12280 25410 12336
rect 25466 12280 28000 12336
rect 25405 12278 28000 12280
rect 10777 12275 10843 12278
rect 25405 12275 25471 12278
rect 27520 12248 28000 12278
rect 11421 12202 11487 12205
rect 16205 12202 16271 12205
rect 11421 12200 16271 12202
rect 11421 12144 11426 12200
rect 11482 12144 16210 12200
rect 16266 12144 16271 12200
rect 11421 12142 16271 12144
rect 11421 12139 11487 12142
rect 16205 12139 16271 12142
rect 18597 12202 18663 12205
rect 21081 12202 21147 12205
rect 24301 12202 24367 12205
rect 18597 12200 24367 12202
rect 18597 12144 18602 12200
rect 18658 12144 21086 12200
rect 21142 12144 24306 12200
rect 24362 12144 24367 12200
rect 18597 12142 24367 12144
rect 18597 12139 18663 12142
rect 21081 12139 21147 12142
rect 24301 12139 24367 12142
rect 11881 12066 11947 12069
rect 7284 12064 11947 12066
rect 7284 12008 11886 12064
rect 11942 12008 11947 12064
rect 7284 12006 11947 12008
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 0 11794 480 11824
rect 3233 11794 3299 11797
rect 0 11792 3299 11794
rect 0 11736 3238 11792
rect 3294 11736 3299 11792
rect 0 11734 3299 11736
rect 0 11704 480 11734
rect 3233 11731 3299 11734
rect 4061 11794 4127 11797
rect 7284 11794 7344 12006
rect 11881 12003 11947 12006
rect 20621 12066 20687 12069
rect 23657 12066 23723 12069
rect 20621 12064 23723 12066
rect 20621 12008 20626 12064
rect 20682 12008 23662 12064
rect 23718 12008 23723 12064
rect 20621 12006 23723 12008
rect 20621 12003 20687 12006
rect 23657 12003 23723 12006
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 11697 11930 11763 11933
rect 14549 11930 14615 11933
rect 11697 11928 14615 11930
rect 11697 11872 11702 11928
rect 11758 11872 14554 11928
rect 14610 11872 14615 11928
rect 11697 11870 14615 11872
rect 11697 11867 11763 11870
rect 14549 11867 14615 11870
rect 18137 11930 18203 11933
rect 20069 11930 20135 11933
rect 24025 11930 24091 11933
rect 18137 11928 24091 11930
rect 18137 11872 18142 11928
rect 18198 11872 20074 11928
rect 20130 11872 24030 11928
rect 24086 11872 24091 11928
rect 18137 11870 24091 11872
rect 18137 11867 18203 11870
rect 20069 11867 20135 11870
rect 24025 11867 24091 11870
rect 4061 11792 7344 11794
rect 4061 11736 4066 11792
rect 4122 11736 7344 11792
rect 4061 11734 7344 11736
rect 11145 11794 11211 11797
rect 15285 11794 15351 11797
rect 11145 11792 15351 11794
rect 11145 11736 11150 11792
rect 11206 11736 15290 11792
rect 15346 11736 15351 11792
rect 11145 11734 15351 11736
rect 4061 11731 4127 11734
rect 11145 11731 11211 11734
rect 15285 11731 15351 11734
rect 22921 11794 22987 11797
rect 27520 11794 28000 11824
rect 22921 11792 28000 11794
rect 22921 11736 22926 11792
rect 22982 11736 28000 11792
rect 22921 11734 28000 11736
rect 22921 11731 22987 11734
rect 27520 11704 28000 11734
rect 9397 11658 9463 11661
rect 12157 11658 12223 11661
rect 9397 11656 12223 11658
rect 9397 11600 9402 11656
rect 9458 11600 12162 11656
rect 12218 11600 12223 11656
rect 9397 11598 12223 11600
rect 9397 11595 9463 11598
rect 12157 11595 12223 11598
rect 19977 11658 20043 11661
rect 23565 11658 23631 11661
rect 19977 11656 23631 11658
rect 19977 11600 19982 11656
rect 20038 11600 23570 11656
rect 23626 11600 23631 11656
rect 19977 11598 23631 11600
rect 19977 11595 20043 11598
rect 23565 11595 23631 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 4429 11386 4495 11389
rect 8385 11386 8451 11389
rect 4429 11384 8451 11386
rect 4429 11328 4434 11384
rect 4490 11328 8390 11384
rect 8446 11328 8451 11384
rect 4429 11326 8451 11328
rect 4429 11323 4495 11326
rect 8385 11323 8451 11326
rect 14181 11386 14247 11389
rect 18137 11386 18203 11389
rect 14181 11384 18203 11386
rect 14181 11328 14186 11384
rect 14242 11328 18142 11384
rect 18198 11328 18203 11384
rect 14181 11326 18203 11328
rect 14181 11323 14247 11326
rect 18137 11323 18203 11326
rect 9213 11250 9279 11253
rect 12065 11250 12131 11253
rect 9213 11248 12131 11250
rect 9213 11192 9218 11248
rect 9274 11192 12070 11248
rect 12126 11192 12131 11248
rect 9213 11190 12131 11192
rect 9213 11187 9279 11190
rect 12065 11187 12131 11190
rect 15745 11250 15811 11253
rect 24945 11250 25011 11253
rect 15745 11248 25011 11250
rect 15745 11192 15750 11248
rect 15806 11192 24950 11248
rect 25006 11192 25011 11248
rect 15745 11190 25011 11192
rect 15745 11187 15811 11190
rect 24945 11187 25011 11190
rect 0 11114 480 11144
rect 8845 11114 8911 11117
rect 0 11112 8911 11114
rect 0 11056 8850 11112
rect 8906 11056 8911 11112
rect 0 11054 8911 11056
rect 0 11024 480 11054
rect 8845 11051 8911 11054
rect 10869 11114 10935 11117
rect 11237 11114 11303 11117
rect 18229 11114 18295 11117
rect 23473 11114 23539 11117
rect 10869 11112 23539 11114
rect 10869 11056 10874 11112
rect 10930 11056 11242 11112
rect 11298 11056 18234 11112
rect 18290 11056 23478 11112
rect 23534 11056 23539 11112
rect 10869 11054 23539 11056
rect 10869 11051 10935 11054
rect 11237 11051 11303 11054
rect 18229 11051 18295 11054
rect 23473 11051 23539 11054
rect 24301 11114 24367 11117
rect 27520 11114 28000 11144
rect 24301 11112 28000 11114
rect 24301 11056 24306 11112
rect 24362 11056 28000 11112
rect 24301 11054 28000 11056
rect 24301 11051 24367 11054
rect 27520 11024 28000 11054
rect 19374 10916 19380 10980
rect 19444 10978 19450 10980
rect 22829 10978 22895 10981
rect 19444 10976 22895 10978
rect 19444 10920 22834 10976
rect 22890 10920 22895 10976
rect 19444 10918 22895 10920
rect 19444 10916 19450 10918
rect 22829 10915 22895 10918
rect 25129 10978 25195 10981
rect 25313 10978 25379 10981
rect 25129 10976 25379 10978
rect 25129 10920 25134 10976
rect 25190 10920 25318 10976
rect 25374 10920 25379 10976
rect 25129 10918 25379 10920
rect 25129 10915 25195 10918
rect 25313 10915 25379 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 8753 10706 8819 10709
rect 2454 10704 8819 10706
rect 2454 10648 8758 10704
rect 8814 10648 8819 10704
rect 2454 10646 8819 10648
rect 0 10570 480 10600
rect 2454 10570 2514 10646
rect 8753 10643 8819 10646
rect 14733 10706 14799 10709
rect 19977 10706 20043 10709
rect 14733 10704 20043 10706
rect 14733 10648 14738 10704
rect 14794 10648 19982 10704
rect 20038 10648 20043 10704
rect 14733 10646 20043 10648
rect 14733 10643 14799 10646
rect 19977 10643 20043 10646
rect 21357 10706 21423 10709
rect 21817 10706 21883 10709
rect 25221 10706 25287 10709
rect 21357 10704 25287 10706
rect 21357 10648 21362 10704
rect 21418 10648 21822 10704
rect 21878 10648 25226 10704
rect 25282 10648 25287 10704
rect 21357 10646 25287 10648
rect 21357 10643 21423 10646
rect 21817 10643 21883 10646
rect 25221 10643 25287 10646
rect 0 10510 2514 10570
rect 10041 10570 10107 10573
rect 15285 10570 15351 10573
rect 17493 10570 17559 10573
rect 10041 10568 17559 10570
rect 10041 10512 10046 10568
rect 10102 10512 15290 10568
rect 15346 10512 17498 10568
rect 17554 10512 17559 10568
rect 10041 10510 17559 10512
rect 0 10480 480 10510
rect 10041 10507 10107 10510
rect 15285 10507 15351 10510
rect 16622 10437 16682 10510
rect 17493 10507 17559 10510
rect 18689 10570 18755 10573
rect 27520 10570 28000 10600
rect 18689 10568 20362 10570
rect 18689 10512 18694 10568
rect 18750 10512 20362 10568
rect 18689 10510 20362 10512
rect 18689 10507 18755 10510
rect 3877 10434 3943 10437
rect 10133 10434 10199 10437
rect 3877 10432 10199 10434
rect 3877 10376 3882 10432
rect 3938 10376 10138 10432
rect 10194 10376 10199 10432
rect 3877 10374 10199 10376
rect 3877 10371 3943 10374
rect 10133 10371 10199 10374
rect 13537 10434 13603 10437
rect 15377 10434 15443 10437
rect 13537 10432 15443 10434
rect 13537 10376 13542 10432
rect 13598 10376 15382 10432
rect 15438 10376 15443 10432
rect 13537 10374 15443 10376
rect 16622 10432 16731 10437
rect 16622 10376 16670 10432
rect 16726 10376 16731 10432
rect 16622 10374 16731 10376
rect 13537 10371 13603 10374
rect 15377 10371 15443 10374
rect 16665 10371 16731 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 20302 10301 20362 10510
rect 24902 10510 28000 10570
rect 4521 10298 4587 10301
rect 10041 10298 10107 10301
rect 4521 10296 10107 10298
rect 4521 10240 4526 10296
rect 4582 10240 10046 10296
rect 10102 10240 10107 10296
rect 4521 10238 10107 10240
rect 4521 10235 4587 10238
rect 10041 10235 10107 10238
rect 13261 10298 13327 10301
rect 18781 10298 18847 10301
rect 20302 10298 20411 10301
rect 24577 10298 24643 10301
rect 13261 10296 18847 10298
rect 13261 10240 13266 10296
rect 13322 10240 18786 10296
rect 18842 10240 18847 10296
rect 13261 10238 18847 10240
rect 20218 10296 24643 10298
rect 20218 10240 20350 10296
rect 20406 10240 24582 10296
rect 24638 10240 24643 10296
rect 20218 10238 24643 10240
rect 13261 10235 13327 10238
rect 18781 10235 18847 10238
rect 20345 10235 20411 10238
rect 24577 10235 24643 10238
rect 13629 10162 13695 10165
rect 24902 10162 24962 10510
rect 27520 10480 28000 10510
rect 13629 10160 24962 10162
rect 13629 10104 13634 10160
rect 13690 10104 24962 10160
rect 13629 10102 24962 10104
rect 13629 10099 13695 10102
rect 0 10026 480 10056
rect 4061 10026 4127 10029
rect 0 10024 4127 10026
rect 0 9968 4066 10024
rect 4122 9968 4127 10024
rect 0 9966 4127 9968
rect 0 9936 480 9966
rect 4061 9963 4127 9966
rect 14181 10026 14247 10029
rect 15653 10026 15719 10029
rect 27520 10026 28000 10056
rect 14181 10024 15719 10026
rect 14181 9968 14186 10024
rect 14242 9968 15658 10024
rect 15714 9968 15719 10024
rect 14181 9966 15719 9968
rect 14181 9963 14247 9966
rect 15653 9963 15719 9966
rect 25822 9966 28000 10026
rect 19977 9890 20043 9893
rect 23841 9890 23907 9893
rect 19977 9888 23907 9890
rect 19977 9832 19982 9888
rect 20038 9832 23846 9888
rect 23902 9832 23907 9888
rect 19977 9830 23907 9832
rect 19977 9827 20043 9830
rect 23841 9827 23907 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 12249 9754 12315 9757
rect 14549 9754 14615 9757
rect 12249 9752 14615 9754
rect 12249 9696 12254 9752
rect 12310 9696 14554 9752
rect 14610 9696 14615 9752
rect 12249 9694 14615 9696
rect 12249 9691 12315 9694
rect 14549 9691 14615 9694
rect 22737 9754 22803 9757
rect 25822 9754 25882 9966
rect 27520 9936 28000 9966
rect 22737 9752 24042 9754
rect 22737 9696 22742 9752
rect 22798 9696 24042 9752
rect 22737 9694 24042 9696
rect 22737 9691 22803 9694
rect 20253 9618 20319 9621
rect 22461 9618 22527 9621
rect 20253 9616 22527 9618
rect 20253 9560 20258 9616
rect 20314 9560 22466 9616
rect 22522 9560 22527 9616
rect 20253 9558 22527 9560
rect 20253 9555 20319 9558
rect 22461 9555 22527 9558
rect 23606 9556 23612 9620
rect 23676 9618 23682 9620
rect 23749 9618 23815 9621
rect 23676 9616 23815 9618
rect 23676 9560 23754 9616
rect 23810 9560 23815 9616
rect 23676 9558 23815 9560
rect 23982 9618 24042 9694
rect 24718 9694 25882 9754
rect 24718 9618 24778 9694
rect 23982 9558 24778 9618
rect 23676 9556 23682 9558
rect 23749 9555 23815 9558
rect 0 9482 480 9512
rect 3693 9482 3759 9485
rect 0 9480 3759 9482
rect 0 9424 3698 9480
rect 3754 9424 3759 9480
rect 0 9422 3759 9424
rect 0 9392 480 9422
rect 3693 9419 3759 9422
rect 8661 9482 8727 9485
rect 9673 9482 9739 9485
rect 8661 9480 9739 9482
rect 8661 9424 8666 9480
rect 8722 9424 9678 9480
rect 9734 9424 9739 9480
rect 8661 9422 9739 9424
rect 8661 9419 8727 9422
rect 9673 9419 9739 9422
rect 22001 9482 22067 9485
rect 27520 9482 28000 9512
rect 22001 9480 28000 9482
rect 22001 9424 22006 9480
rect 22062 9424 28000 9480
rect 22001 9422 28000 9424
rect 22001 9419 22067 9422
rect 27520 9392 28000 9422
rect 2957 9346 3023 9349
rect 9857 9346 9923 9349
rect 2957 9344 9923 9346
rect 2957 9288 2962 9344
rect 3018 9288 9862 9344
rect 9918 9288 9923 9344
rect 2957 9286 9923 9288
rect 2957 9283 3023 9286
rect 9857 9283 9923 9286
rect 12065 9346 12131 9349
rect 21725 9346 21791 9349
rect 24853 9346 24919 9349
rect 12065 9344 17234 9346
rect 12065 9288 12070 9344
rect 12126 9288 17234 9344
rect 12065 9286 17234 9288
rect 12065 9283 12131 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 3509 9210 3575 9213
rect 9949 9210 10015 9213
rect 3509 9208 10015 9210
rect 3509 9152 3514 9208
rect 3570 9152 9954 9208
rect 10010 9152 10015 9208
rect 3509 9150 10015 9152
rect 3509 9147 3575 9150
rect 9949 9147 10015 9150
rect 1853 9074 1919 9077
rect 17174 9074 17234 9286
rect 21725 9344 24919 9346
rect 21725 9288 21730 9344
rect 21786 9288 24858 9344
rect 24914 9288 24919 9344
rect 21725 9286 24919 9288
rect 21725 9283 21791 9286
rect 24853 9283 24919 9286
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 23841 9210 23907 9213
rect 22510 9208 23907 9210
rect 22510 9152 23846 9208
rect 23902 9152 23907 9208
rect 22510 9150 23907 9152
rect 22510 9074 22570 9150
rect 23841 9147 23907 9150
rect 24669 9212 24735 9213
rect 24669 9208 24716 9212
rect 24780 9210 24786 9212
rect 24669 9152 24674 9208
rect 24669 9148 24716 9152
rect 24780 9150 24826 9210
rect 24780 9148 24786 9150
rect 24669 9147 24735 9148
rect 1853 9072 15946 9074
rect 1853 9016 1858 9072
rect 1914 9016 15946 9072
rect 1853 9014 15946 9016
rect 17174 9014 22570 9074
rect 22645 9074 22711 9077
rect 24761 9074 24827 9077
rect 22645 9072 24827 9074
rect 22645 9016 22650 9072
rect 22706 9016 24766 9072
rect 24822 9016 24827 9072
rect 22645 9014 24827 9016
rect 1853 9011 1919 9014
rect 0 8938 480 8968
rect 8017 8938 8083 8941
rect 0 8878 2698 8938
rect 0 8848 480 8878
rect 2638 8802 2698 8878
rect 8017 8936 15762 8938
rect 8017 8880 8022 8936
rect 8078 8880 15762 8936
rect 8017 8878 15762 8880
rect 8017 8875 8083 8878
rect 2638 8742 2882 8802
rect 2822 8530 2882 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 15702 8666 15762 8878
rect 15886 8802 15946 9014
rect 22645 9011 22711 9014
rect 24761 9011 24827 9014
rect 16113 8938 16179 8941
rect 18505 8938 18571 8941
rect 16113 8936 18571 8938
rect 16113 8880 16118 8936
rect 16174 8880 18510 8936
rect 18566 8880 18571 8936
rect 16113 8878 18571 8880
rect 16113 8875 16179 8878
rect 18505 8875 18571 8878
rect 18873 8938 18939 8941
rect 21541 8938 21607 8941
rect 18873 8936 21607 8938
rect 18873 8880 18878 8936
rect 18934 8880 21546 8936
rect 21602 8880 21607 8936
rect 18873 8878 21607 8880
rect 18873 8875 18939 8878
rect 21541 8875 21607 8878
rect 22829 8938 22895 8941
rect 27520 8938 28000 8968
rect 22829 8936 28000 8938
rect 22829 8880 22834 8936
rect 22890 8880 28000 8936
rect 22829 8878 28000 8880
rect 22829 8875 22895 8878
rect 27520 8848 28000 8878
rect 21265 8802 21331 8805
rect 23473 8802 23539 8805
rect 15886 8800 21331 8802
rect 15886 8744 21270 8800
rect 21326 8744 21331 8800
rect 15886 8742 21331 8744
rect 21265 8739 21331 8742
rect 21406 8800 23539 8802
rect 21406 8744 23478 8800
rect 23534 8744 23539 8800
rect 21406 8742 23539 8744
rect 20897 8666 20963 8669
rect 21406 8666 21466 8742
rect 23473 8739 23539 8742
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 15702 8664 21466 8666
rect 15702 8608 20902 8664
rect 20958 8608 21466 8664
rect 15702 8606 21466 8608
rect 21541 8666 21607 8669
rect 24117 8666 24183 8669
rect 21541 8664 24183 8666
rect 21541 8608 21546 8664
rect 21602 8608 24122 8664
rect 24178 8608 24183 8664
rect 21541 8606 24183 8608
rect 20897 8603 20963 8606
rect 21541 8603 21607 8606
rect 24117 8603 24183 8606
rect 13261 8530 13327 8533
rect 2822 8528 13327 8530
rect 2822 8472 13266 8528
rect 13322 8472 13327 8528
rect 2822 8470 13327 8472
rect 13261 8467 13327 8470
rect 15377 8530 15443 8533
rect 19885 8530 19951 8533
rect 15377 8528 19951 8530
rect 15377 8472 15382 8528
rect 15438 8472 19890 8528
rect 19946 8472 19951 8528
rect 15377 8470 19951 8472
rect 15377 8467 15443 8470
rect 19885 8467 19951 8470
rect 21265 8530 21331 8533
rect 23565 8530 23631 8533
rect 21265 8528 23631 8530
rect 21265 8472 21270 8528
rect 21326 8472 23570 8528
rect 23626 8472 23631 8528
rect 21265 8470 23631 8472
rect 21265 8467 21331 8470
rect 23565 8467 23631 8470
rect 20897 8394 20963 8397
rect 23841 8394 23907 8397
rect 20897 8392 23907 8394
rect 20897 8336 20902 8392
rect 20958 8336 23846 8392
rect 23902 8336 23907 8392
rect 20897 8334 23907 8336
rect 20897 8331 20963 8334
rect 23841 8331 23907 8334
rect 0 8258 480 8288
rect 6545 8258 6611 8261
rect 0 8256 6611 8258
rect 0 8200 6550 8256
rect 6606 8200 6611 8256
rect 0 8198 6611 8200
rect 0 8168 480 8198
rect 6545 8195 6611 8198
rect 15101 8258 15167 8261
rect 16757 8258 16823 8261
rect 15101 8256 16823 8258
rect 15101 8200 15106 8256
rect 15162 8200 16762 8256
rect 16818 8200 16823 8256
rect 15101 8198 16823 8200
rect 15101 8195 15167 8198
rect 16757 8195 16823 8198
rect 23974 8196 23980 8260
rect 24044 8258 24050 8260
rect 27520 8258 28000 8288
rect 24044 8198 28000 8258
rect 24044 8196 24050 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 13813 8122 13879 8125
rect 15929 8122 15995 8125
rect 13813 8120 15995 8122
rect 13813 8064 13818 8120
rect 13874 8064 15934 8120
rect 15990 8064 15995 8120
rect 13813 8062 15995 8064
rect 13813 8059 13879 8062
rect 15929 8059 15995 8062
rect 9765 7986 9831 7989
rect 12157 7986 12223 7989
rect 9765 7984 12223 7986
rect 9765 7928 9770 7984
rect 9826 7928 12162 7984
rect 12218 7928 12223 7984
rect 9765 7926 12223 7928
rect 9765 7923 9831 7926
rect 12157 7923 12223 7926
rect 14549 7986 14615 7989
rect 19333 7986 19399 7989
rect 14549 7984 19399 7986
rect 14549 7928 14554 7984
rect 14610 7928 19338 7984
rect 19394 7928 19399 7984
rect 14549 7926 19399 7928
rect 14549 7923 14615 7926
rect 19333 7923 19399 7926
rect 20805 7986 20871 7989
rect 24761 7986 24827 7989
rect 20805 7984 24827 7986
rect 20805 7928 20810 7984
rect 20866 7928 24766 7984
rect 24822 7928 24827 7984
rect 20805 7926 24827 7928
rect 20805 7923 20871 7926
rect 24761 7923 24827 7926
rect 16205 7850 16271 7853
rect 4846 7848 16271 7850
rect 4846 7792 16210 7848
rect 16266 7792 16271 7848
rect 4846 7790 16271 7792
rect 0 7714 480 7744
rect 0 7654 2698 7714
rect 0 7624 480 7654
rect 2638 7578 2698 7654
rect 4846 7578 4906 7790
rect 16205 7787 16271 7790
rect 18229 7850 18295 7853
rect 21081 7850 21147 7853
rect 18229 7848 21147 7850
rect 18229 7792 18234 7848
rect 18290 7792 21086 7848
rect 21142 7792 21147 7848
rect 18229 7790 21147 7792
rect 18229 7787 18295 7790
rect 21081 7787 21147 7790
rect 24117 7850 24183 7853
rect 24117 7848 24778 7850
rect 24117 7792 24122 7848
rect 24178 7792 24778 7848
rect 24117 7790 24778 7792
rect 24117 7787 24183 7790
rect 6545 7714 6611 7717
rect 14181 7714 14247 7717
rect 6545 7712 14247 7714
rect 6545 7656 6550 7712
rect 6606 7656 14186 7712
rect 14242 7656 14247 7712
rect 6545 7654 14247 7656
rect 24718 7714 24778 7790
rect 27520 7714 28000 7744
rect 24718 7654 28000 7714
rect 6545 7651 6611 7654
rect 14181 7651 14247 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7654
rect 24277 7583 24597 7584
rect 2638 7518 4906 7578
rect 7465 7578 7531 7581
rect 14733 7578 14799 7581
rect 7465 7576 14799 7578
rect 7465 7520 7470 7576
rect 7526 7520 14738 7576
rect 14794 7520 14799 7576
rect 7465 7518 14799 7520
rect 7465 7515 7531 7518
rect 14733 7515 14799 7518
rect 10133 7442 10199 7445
rect 23657 7442 23723 7445
rect 10133 7440 23723 7442
rect 10133 7384 10138 7440
rect 10194 7384 23662 7440
rect 23718 7384 23723 7440
rect 10133 7382 23723 7384
rect 10133 7379 10199 7382
rect 23657 7379 23723 7382
rect 12709 7306 12775 7309
rect 23749 7306 23815 7309
rect 12709 7304 23815 7306
rect 12709 7248 12714 7304
rect 12770 7248 23754 7304
rect 23810 7248 23815 7304
rect 12709 7246 23815 7248
rect 12709 7243 12775 7246
rect 23749 7243 23815 7246
rect 0 7170 480 7200
rect 2957 7170 3023 7173
rect 0 7168 3023 7170
rect 0 7112 2962 7168
rect 3018 7112 3023 7168
rect 0 7110 3023 7112
rect 0 7080 480 7110
rect 2957 7107 3023 7110
rect 23841 7170 23907 7173
rect 27520 7170 28000 7200
rect 23841 7168 28000 7170
rect 23841 7112 23846 7168
rect 23902 7112 28000 7168
rect 23841 7110 28000 7112
rect 23841 7107 23907 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 27520 7080 28000 7110
rect 19610 7039 19930 7040
rect 10777 6898 10843 6901
rect 19149 6898 19215 6901
rect 10777 6896 17234 6898
rect 10777 6840 10782 6896
rect 10838 6840 17234 6896
rect 10777 6838 17234 6840
rect 10777 6835 10843 6838
rect 4061 6762 4127 6765
rect 14365 6762 14431 6765
rect 4061 6760 14431 6762
rect 4061 6704 4066 6760
rect 4122 6704 14370 6760
rect 14426 6704 14431 6760
rect 4061 6702 14431 6704
rect 17174 6762 17234 6838
rect 19149 6896 24962 6898
rect 19149 6840 19154 6896
rect 19210 6840 24962 6896
rect 19149 6838 24962 6840
rect 19149 6835 19215 6838
rect 23657 6762 23723 6765
rect 17174 6760 23723 6762
rect 17174 6704 23662 6760
rect 23718 6704 23723 6760
rect 17174 6702 23723 6704
rect 4061 6699 4127 6702
rect 14365 6699 14431 6702
rect 23657 6699 23723 6702
rect 0 6626 480 6656
rect 17585 6626 17651 6629
rect 22277 6626 22343 6629
rect 0 6566 2698 6626
rect 0 6536 480 6566
rect 2638 6490 2698 6566
rect 17585 6624 22343 6626
rect 17585 6568 17590 6624
rect 17646 6568 22282 6624
rect 22338 6568 22343 6624
rect 17585 6566 22343 6568
rect 24902 6626 24962 6838
rect 27520 6626 28000 6656
rect 24902 6566 28000 6626
rect 17585 6563 17651 6566
rect 22277 6563 22343 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6566
rect 24277 6495 24597 6496
rect 2638 6430 2882 6490
rect 2822 6354 2882 6430
rect 12617 6354 12683 6357
rect 2822 6352 12683 6354
rect 2822 6296 12622 6352
rect 12678 6296 12683 6352
rect 2822 6294 12683 6296
rect 12617 6291 12683 6294
rect 0 6082 480 6112
rect 4061 6082 4127 6085
rect 0 6080 4127 6082
rect 0 6024 4066 6080
rect 4122 6024 4127 6080
rect 0 6022 4127 6024
rect 0 5992 480 6022
rect 4061 6019 4127 6022
rect 23422 6020 23428 6084
rect 23492 6082 23498 6084
rect 27520 6082 28000 6112
rect 23492 6022 28000 6082
rect 23492 6020 23498 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 4061 5402 4127 5405
rect 27520 5402 28000 5432
rect 0 5400 4127 5402
rect 0 5344 4066 5400
rect 4122 5344 4127 5400
rect 0 5342 4127 5344
rect 0 5312 480 5342
rect 4061 5339 4127 5342
rect 24718 5342 28000 5402
rect 3969 5266 4035 5269
rect 18781 5266 18847 5269
rect 3969 5264 18847 5266
rect 3969 5208 3974 5264
rect 4030 5208 18786 5264
rect 18842 5208 18847 5264
rect 3969 5206 18847 5208
rect 3969 5203 4035 5206
rect 18781 5203 18847 5206
rect 23565 5266 23631 5269
rect 24718 5266 24778 5342
rect 27520 5312 28000 5342
rect 23565 5264 24778 5266
rect 23565 5208 23570 5264
rect 23626 5208 24778 5264
rect 23565 5206 24778 5208
rect 23565 5203 23631 5206
rect 18229 5130 18295 5133
rect 18229 5128 22064 5130
rect 18229 5072 18234 5128
rect 18290 5072 22064 5128
rect 18229 5070 22064 5072
rect 18229 5067 18295 5070
rect 10685 4994 10751 4997
rect 17401 4994 17467 4997
rect 10685 4992 17467 4994
rect 10685 4936 10690 4992
rect 10746 4936 17406 4992
rect 17462 4936 17467 4992
rect 10685 4934 17467 4936
rect 22004 4994 22064 5070
rect 22004 4934 22202 4994
rect 10685 4931 10751 4934
rect 17401 4931 17467 4934
rect 10277 4928 10597 4929
rect 0 4858 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 3877 4858 3943 4861
rect 0 4856 3943 4858
rect 0 4800 3882 4856
rect 3938 4800 3943 4856
rect 0 4798 3943 4800
rect 22142 4858 22202 4934
rect 27520 4858 28000 4888
rect 22142 4798 28000 4858
rect 0 4768 480 4798
rect 3877 4795 3943 4798
rect 27520 4768 28000 4798
rect 4061 4722 4127 4725
rect 20437 4722 20503 4725
rect 4061 4720 20503 4722
rect 4061 4664 4066 4720
rect 4122 4664 20442 4720
rect 20498 4664 20503 4720
rect 4061 4662 20503 4664
rect 4061 4659 4127 4662
rect 20437 4659 20503 4662
rect 16941 4586 17007 4589
rect 23565 4586 23631 4589
rect 16941 4584 23631 4586
rect 16941 4528 16946 4584
rect 17002 4528 23570 4584
rect 23626 4528 23631 4584
rect 16941 4526 23631 4528
rect 16941 4523 17007 4526
rect 23565 4523 23631 4526
rect 5610 4384 5930 4385
rect 0 4314 480 4344
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 3969 4314 4035 4317
rect 27520 4314 28000 4344
rect 0 4312 4035 4314
rect 0 4256 3974 4312
rect 4030 4256 4035 4312
rect 0 4254 4035 4256
rect 0 4224 480 4254
rect 3969 4251 4035 4254
rect 24718 4254 28000 4314
rect 23473 4178 23539 4181
rect 24718 4178 24778 4254
rect 27520 4224 28000 4254
rect 23473 4176 24778 4178
rect 23473 4120 23478 4176
rect 23534 4120 24778 4176
rect 23473 4118 24778 4120
rect 23473 4115 23539 4118
rect 17125 4042 17191 4045
rect 2454 4040 17191 4042
rect 2454 3984 17130 4040
rect 17186 3984 17191 4040
rect 2454 3982 17191 3984
rect 0 3770 480 3800
rect 2454 3770 2514 3982
rect 17125 3979 17191 3982
rect 20161 3906 20227 3909
rect 23473 3906 23539 3909
rect 20161 3904 23539 3906
rect 20161 3848 20166 3904
rect 20222 3848 23478 3904
rect 23534 3848 23539 3904
rect 20161 3846 23539 3848
rect 20161 3843 20227 3846
rect 23473 3843 23539 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 0 3710 2514 3770
rect 22185 3770 22251 3773
rect 27520 3770 28000 3800
rect 22185 3768 28000 3770
rect 22185 3712 22190 3768
rect 22246 3712 28000 3768
rect 22185 3710 28000 3712
rect 0 3680 480 3710
rect 22185 3707 22251 3710
rect 27520 3680 28000 3710
rect 3141 3634 3207 3637
rect 11881 3634 11947 3637
rect 3141 3632 11947 3634
rect 3141 3576 3146 3632
rect 3202 3576 11886 3632
rect 11942 3576 11947 3632
rect 3141 3574 11947 3576
rect 3141 3571 3207 3574
rect 11881 3571 11947 3574
rect 18505 3634 18571 3637
rect 22001 3634 22067 3637
rect 18505 3632 22067 3634
rect 18505 3576 18510 3632
rect 18566 3576 22006 3632
rect 22062 3576 22067 3632
rect 18505 3574 22067 3576
rect 18505 3571 18571 3574
rect 22001 3571 22067 3574
rect 10685 3498 10751 3501
rect 2822 3496 10751 3498
rect 2822 3440 10690 3496
rect 10746 3440 10751 3496
rect 2822 3438 10751 3440
rect 2822 3362 2882 3438
rect 10685 3435 10751 3438
rect 11053 3498 11119 3501
rect 23197 3498 23263 3501
rect 11053 3496 23263 3498
rect 11053 3440 11058 3496
rect 11114 3440 23202 3496
rect 23258 3440 23263 3496
rect 11053 3438 23263 3440
rect 11053 3435 11119 3438
rect 23197 3435 23263 3438
rect 2638 3302 2882 3362
rect 0 3226 480 3256
rect 2638 3226 2698 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 27520 3226 28000 3256
rect 0 3166 2698 3226
rect 24902 3166 28000 3226
rect 0 3136 480 3166
rect 17033 3090 17099 3093
rect 24902 3090 24962 3166
rect 27520 3136 28000 3166
rect 17033 3088 24962 3090
rect 17033 3032 17038 3088
rect 17094 3032 24962 3088
rect 17033 3030 24962 3032
rect 17033 3027 17099 3030
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 3509 2682 3575 2685
rect 3190 2680 3575 2682
rect 3190 2624 3514 2680
rect 3570 2624 3575 2680
rect 3190 2622 3575 2624
rect 0 2546 480 2576
rect 3190 2546 3250 2622
rect 3509 2619 3575 2622
rect 11973 2546 12039 2549
rect 0 2486 3250 2546
rect 3374 2544 12039 2546
rect 3374 2488 11978 2544
rect 12034 2488 12039 2544
rect 3374 2486 12039 2488
rect 0 2456 480 2486
rect 0 2002 480 2032
rect 3374 2002 3434 2486
rect 11973 2483 12039 2486
rect 23565 2546 23631 2549
rect 27520 2546 28000 2576
rect 23565 2544 28000 2546
rect 23565 2488 23570 2544
rect 23626 2488 28000 2544
rect 23565 2486 28000 2488
rect 23565 2483 23631 2486
rect 27520 2456 28000 2486
rect 4613 2410 4679 2413
rect 11973 2410 12039 2413
rect 4613 2408 12039 2410
rect 4613 2352 4618 2408
rect 4674 2352 11978 2408
rect 12034 2352 12039 2408
rect 4613 2350 12039 2352
rect 4613 2347 4679 2350
rect 11973 2347 12039 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 24117 2138 24183 2141
rect 17174 2136 24183 2138
rect 17174 2080 24122 2136
rect 24178 2080 24183 2136
rect 17174 2078 24183 2080
rect 17174 2002 17234 2078
rect 24117 2075 24183 2078
rect 0 1942 3434 2002
rect 3558 1942 17234 2002
rect 23749 2002 23815 2005
rect 27520 2002 28000 2032
rect 23749 2000 28000 2002
rect 23749 1944 23754 2000
rect 23810 1944 28000 2000
rect 23749 1942 28000 1944
rect 0 1912 480 1942
rect 3558 1730 3618 1942
rect 23749 1939 23815 1942
rect 27520 1912 28000 1942
rect 3374 1670 3618 1730
rect 0 1458 480 1488
rect 3374 1458 3434 1670
rect 3509 1594 3575 1597
rect 11789 1594 11855 1597
rect 3509 1592 11855 1594
rect 3509 1536 3514 1592
rect 3570 1536 11794 1592
rect 11850 1536 11855 1592
rect 3509 1534 11855 1536
rect 3509 1531 3575 1534
rect 11789 1531 11855 1534
rect 14641 1594 14707 1597
rect 14641 1592 27538 1594
rect 14641 1536 14646 1592
rect 14702 1536 27538 1592
rect 14641 1534 27538 1536
rect 14641 1531 14707 1534
rect 0 1398 3434 1458
rect 27478 1488 27538 1534
rect 27478 1398 28000 1488
rect 0 1368 480 1398
rect 27520 1368 28000 1398
rect 0 914 480 944
rect 3141 914 3207 917
rect 0 912 3207 914
rect 0 856 3146 912
rect 3202 856 3207 912
rect 0 854 3207 856
rect 0 824 480 854
rect 3141 851 3207 854
rect 23473 914 23539 917
rect 27520 914 28000 944
rect 23473 912 28000 914
rect 23473 856 23478 912
rect 23534 856 28000 912
rect 23473 854 28000 856
rect 23473 851 23539 854
rect 27520 824 28000 854
rect 0 370 480 400
rect 3233 370 3299 373
rect 0 368 3299 370
rect 0 312 3238 368
rect 3294 312 3299 368
rect 0 310 3299 312
rect 0 280 480 310
rect 3233 307 3299 310
rect 24669 370 24735 373
rect 27520 370 28000 400
rect 24669 368 28000 370
rect 24669 312 24674 368
rect 24730 312 28000 368
rect 24669 310 28000 312
rect 24669 307 24735 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 9444 24924 9508 24988
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 9628 24108 9692 24172
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 11100 23488 11164 23492
rect 11100 23432 11114 23488
rect 11114 23432 11164 23488
rect 11100 23428 11164 23432
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 11100 23020 11164 23084
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 9628 21116 9692 21180
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 9628 20436 9692 20500
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 11100 19680 11164 19684
rect 11100 19624 11150 19680
rect 11150 19624 11164 19680
rect 11100 19620 11164 19624
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 23612 18940 23676 19004
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 22140 18456 22204 18460
rect 22140 18400 22154 18456
rect 22154 18400 22204 18456
rect 22140 18396 22204 18400
rect 19380 17988 19444 18052
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 8340 17640 8404 17644
rect 8340 17584 8390 17640
rect 8390 17584 8404 17640
rect 8340 17580 8404 17584
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 23428 16492 23492 16556
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 23980 15540 24044 15604
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 22140 14860 22204 14924
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 24716 14316 24780 14380
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 23428 13016 23492 13020
rect 23428 12960 23478 13016
rect 23478 12960 23492 13016
rect 23428 12956 23492 12960
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 8340 12276 8404 12340
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 19380 10916 19444 10980
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 23612 9556 23676 9620
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 24716 9208 24780 9212
rect 24716 9152 24730 9208
rect 24730 9152 24780 9208
rect 24716 9148 24780 9152
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 23980 8196 24044 8260
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 23428 6020 23492 6084
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 9443 24988 9509 24989
rect 9443 24924 9444 24988
rect 9508 24924 9509 24988
rect 9443 24923 9509 24924
rect 9446 24170 9506 24923
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 9627 24172 9693 24173
rect 9627 24170 9628 24172
rect 9446 24110 9628 24170
rect 9627 24108 9628 24110
rect 9692 24108 9693 24172
rect 9627 24107 9693 24108
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 10277 23424 10597 24448
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 11099 23492 11165 23493
rect 11099 23428 11100 23492
rect 11164 23428 11165 23492
rect 11099 23427 11165 23428
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 11102 23085 11162 23427
rect 11099 23084 11165 23085
rect 11099 23020 11100 23084
rect 11164 23020 11165 23084
rect 11099 23019 11165 23020
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 9627 21180 9693 21181
rect 9627 21116 9628 21180
rect 9692 21116 9693 21180
rect 9627 21115 9693 21116
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 9630 20501 9690 21115
rect 9627 20500 9693 20501
rect 9627 20436 9628 20500
rect 9692 20436 9693 20500
rect 9627 20435 9693 20436
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 11102 19685 11162 23019
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 11099 19684 11165 19685
rect 11099 19620 11100 19684
rect 11164 19620 11165 19684
rect 11099 19619 11165 19620
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 8339 17644 8405 17645
rect 8339 17580 8340 17644
rect 8404 17580 8405 17644
rect 8339 17579 8405 17580
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 8342 12341 8402 17579
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 8339 12340 8405 12341
rect 8339 12276 8340 12340
rect 8404 12276 8405 12340
rect 8339 12275 8405 12276
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19379 18052 19445 18053
rect 19379 17988 19380 18052
rect 19444 17988 19445 18052
rect 19379 17987 19445 17988
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 19382 10981 19442 17987
rect 19610 17984 19930 19008
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 23611 19004 23677 19005
rect 23611 18940 23612 19004
rect 23676 18940 23677 19004
rect 23611 18939 23677 18940
rect 22139 18460 22205 18461
rect 22139 18396 22140 18460
rect 22204 18396 22205 18460
rect 22139 18395 22205 18396
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 22142 14925 22202 18395
rect 23427 16556 23493 16557
rect 23427 16492 23428 16556
rect 23492 16492 23493 16556
rect 23427 16491 23493 16492
rect 22139 14924 22205 14925
rect 22139 14860 22140 14924
rect 22204 14860 22205 14924
rect 22139 14859 22205 14860
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 23430 13021 23490 16491
rect 23427 13020 23493 13021
rect 23427 12956 23428 13020
rect 23492 12956 23493 13020
rect 23427 12955 23493 12956
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19379 10980 19445 10981
rect 19379 10916 19380 10980
rect 19444 10916 19445 10980
rect 19379 10915 19445 10916
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 23430 6085 23490 12955
rect 23614 9621 23674 18939
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 23979 15604 24045 15605
rect 23979 15540 23980 15604
rect 24044 15540 24045 15604
rect 23979 15539 24045 15540
rect 23611 9620 23677 9621
rect 23611 9556 23612 9620
rect 23676 9556 23677 9620
rect 23611 9555 23677 9556
rect 23982 8261 24042 15539
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24715 14380 24781 14381
rect 24715 14316 24716 14380
rect 24780 14316 24781 14380
rect 24715 14315 24781 14316
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24718 9213 24778 14315
rect 24715 9212 24781 9213
rect 24715 9148 24716 9212
rect 24780 9148 24781 9212
rect 24715 9147 24781 9148
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 23979 8260 24045 8261
rect 23979 8196 23980 8260
rect 24044 8196 24045 8260
rect 23979 8195 24045 8196
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 23427 6084 23493 6085
rect 23427 6020 23428 6084
rect 23492 6020 23493 6084
rect 23427 6019 23493 6020
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_167
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_176
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_180
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_249
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_261
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_273
timestamp 1586364061
transform 1 0 26220 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_170
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_183
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_187
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_200
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_203
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_207
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_1  mux_right_track_16.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_248
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_260
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_8_272
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_139
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_151
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_158
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _062_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _065_
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_221
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_238
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 590 592
use scs8hd_conb_1  _033_
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24104 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_248
timestamp 1586364061
transform 1 0 23920 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_252
timestamp 1586364061
transform 1 0 24288 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_259
timestamp 1586364061
transform 1 0 24932 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_263
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_275
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_126
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_130
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _061_
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_159
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_1  mux_top_track_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_222
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_234
timestamp 1586364061
transform 1 0 22632 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_238
timestamp 1586364061
transform 1 0 23000 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_1  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24748 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_249
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_260
timestamp 1586364061
transform 1 0 25024 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 774 592
use scs8hd_conb_1  _063_
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_137
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_141
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_163
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_190
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_207
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_224
timestamp 1586364061
transform 1 0 21712 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24104 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_239
timestamp 1586364061
transform 1 0 23092 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_248
timestamp 1586364061
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_252
timestamp 1586364061
transform 1 0 24288 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_259
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_263
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_267
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_275
timestamp 1586364061
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_12_99
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 406 592
use scs8hd_conb_1  _064_
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 774 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_170
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_193
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_197
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_204
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_2  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_241
timestamp 1586364061
transform 1 0 23276 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_259
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_271
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_86
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_99
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_112
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 12512 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_133
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_14_139
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_158
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_160
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_177
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_185
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_189
timestamp 1586364061
transform 1 0 18492 0 -1 10336
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_6  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_206
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_218
timestamp 1586364061
transform 1 0 21160 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_216
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_225
timestamp 1586364061
transform 1 0 21804 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_222
timestamp 1586364061
transform 1 0 21528 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_219
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21620 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_245
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_249
timestamp 1586364061
transform 1 0 24012 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_251
timestamp 1586364061
transform 1 0 24196 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24380 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_266
timestamp 1586364061
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_262
timestamp 1586364061
transform 1 0 25208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_263
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 25392 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_275
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_267
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_70
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_85
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_34.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_146
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_195
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 1786 592
use scs8hd_buf_1  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_210
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_213
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_266
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_270
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_51
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 774 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_73
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_36.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_100
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_121
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_134
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1786 592
use scs8hd_buf_1  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_173
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_177
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_182
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 20976 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 21528 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_220
timestamp 1586364061
transform 1 0 21344 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_38.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_264
timestamp 1586364061
transform 1 0 25392 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_268
timestamp 1586364061
transform 1 0 25760 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_6
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_10
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_30
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_36
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_43
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_55
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_67
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_34.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_84
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_36.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_128
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_151
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_168
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_223
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_227
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 406 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 26128 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_260
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_270
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_274
timestamp 1586364061
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_1  mux_left_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_18
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_38
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_42
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_75
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_30.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_87
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_34.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_107
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_177
timestamp 1586364061
transform 1 0 17388 0 -1 12512
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_183
timestamp 1586364061
transform 1 0 17940 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_186
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22172 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21804 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_223
timestamp 1586364061
transform 1 0 21620 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_250
timestamp 1586364061
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_254
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_267
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _083_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_30
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_70
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 1786 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_119
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 12512 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_131
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_34.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_20_146
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_142
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_162
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_165
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_161
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_38.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_193
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_189
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_216
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21344 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_222
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_235
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_219
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_243
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23276 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_256
timestamp 1586364061
transform 1 0 24656 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_266
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_36.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25392 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_267
timestamp 1586364061
transform 1 0 25668 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_274
timestamp 1586364061
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_270
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26128 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 406 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_19
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use scs8hd_conb_1  _059_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_30.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_60
timestamp 1586364061
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_65
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_84
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_88
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_111
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_115
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 130 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_36.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_126
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_170
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_38.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_180
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_209
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_213
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_217
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_234
timestamp 1586364061
transform 1 0 22632 0 1 13600
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_266
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_270
timestamp 1586364061
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_274
timestamp 1586364061
transform 1 0 26312 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_buf_1  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_12
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4324 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_29
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_37
timestamp 1586364061
transform 1 0 4508 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_54
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_77
timestamp 1586364061
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_30.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_81
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_85
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_116
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_buf_1  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12144 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_6  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16192 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_160
timestamp 1586364061
transform 1 0 15824 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_200
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_204
timestamp 1586364061
transform 1 0 19872 0 -1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22908 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_234
timestamp 1586364061
transform 1 0 22632 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_243
timestamp 1586364061
transform 1 0 23460 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_256
timestamp 1586364061
transform 1 0 24656 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_38.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25392 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_260
timestamp 1586364061
transform 1 0 25024 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_267
timestamp 1586364061
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_28.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_36.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_141
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_166
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_224
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_228
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23828 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_256
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 25392 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_260
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_268
timestamp 1586364061
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_272
timestamp 1586364061
transform 1 0 26128 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_17
timestamp 1586364061
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_21
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_25
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_77
timestamp 1586364061
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 866 592
use scs8hd_buf_1  mux_top_track_30.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_28.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_34.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13892 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_146
timestamp 1586364061
transform 1 0 14536 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_157
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16468 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18952 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_203
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_207
timestamp 1586364061
transform 1 0 20148 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21528 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21344 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_219
timestamp 1586364061
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23460 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_241
timestamp 1586364061
transform 1 0 23276 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_245
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_258
timestamp 1586364061
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_270
timestamp 1586364061
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 1786 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_40
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_30.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_81
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_91
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_28.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_155
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_201
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_218
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_231
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_264
timestamp 1586364061
transform 1 0 25392 0 1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_29
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_33
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_37
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_40
timestamp 1586364061
transform 1 0 4784 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_58
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_54
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_50
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_66
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_70
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_94
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_102
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_28.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_buf_1  mux_top_track_28.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_134
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_130
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_135
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_146
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16192 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15824 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_162
timestamp 1586364061
transform 1 0 16008 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_188
timestamp 1586364061
transform 1 0 18400 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_185
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_189
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18676 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18860 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 19872 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_214
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_221
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_228
timestamp 1586364061
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_235
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_232
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22264 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23000 0 -1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_257
timestamp 1586364061
transform 1 0 24748 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_269
timestamp 1586364061
transform 1 0 25852 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_264
timestamp 1586364061
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_268
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1472 0 -1 17952
box -38 -48 1786 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_63
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_76
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15364 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16928 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_164
timestamp 1586364061
transform 1 0 16192 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_191
timestamp 1586364061
transform 1 0 18676 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  FILLER_28_197
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19504 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_234
timestamp 1586364061
transform 1 0 22632 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_238
timestamp 1586364061
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23368 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24380 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23184 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24748 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_255
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 25484 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1472 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_13
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_17
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_29_21
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_41
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_45
timestamp 1586364061
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_65
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_82
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_109
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 130 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_162
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_166
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 314 592
use scs8hd_conb_1  _060_
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_192
timestamp 1586364061
transform 1 0 18768 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_219
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_223
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_254
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 26128 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_270
timestamp 1586364061
transform 1 0 25944 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_274
timestamp 1586364061
transform 1 0 26312 0 1 17952
box -38 -48 314 592
use scs8hd_conb_1  _056_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_10
timestamp 1586364061
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_29
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_45
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_60
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9844 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_81
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_86
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11408 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_104
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_108
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_131
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_135
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_139
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 314 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_158
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15916 0 -1 19040
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17296 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_170
timestamp 1586364061
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_174
timestamp 1586364061
transform 1 0 17112 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_187
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_191
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_204
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_208
timestamp 1586364061
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_4  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 21804 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 22816 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 21620 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 21252 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_221
timestamp 1586364061
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_234
timestamp 1586364061
transform 1 0 22632 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_238
timestamp 1586364061
transform 1 0 23000 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23368 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23184 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 24380 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 24748 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_255
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25484 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_267
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_12
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_16
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_20
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_24
timestamp 1586364061
transform 1 0 3312 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_81
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_138
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_22.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_142
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_165
timestamp 1586364061
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_169
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20976 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_203
timestamp 1586364061
transform 1 0 19780 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_212
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 22908 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_235
timestamp 1586364061
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_239
timestamp 1586364061
transform 1 0 23092 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_264
timestamp 1586364061
transform 1 0 25392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_268
timestamp 1586364061
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_272
timestamp 1586364061
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_10
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_29
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5888 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_41
timestamp 1586364061
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_45
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_49
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_71
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_75
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_87
timestamp 1586364061
transform 1 0 9108 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 11960 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 11592 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_112
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_116
timestamp 1586364061
transform 1 0 11776 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 12144 0 -1 20128
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_124
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_128
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_132
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_167
timestamp 1586364061
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_171
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_18.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18308 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17664 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_182
timestamp 1586364061
transform 1 0 17848 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21068 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_206
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 21252 0 -1 20128
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 22356 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 21896 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_223
timestamp 1586364061
transform 1 0 21620 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_228
timestamp 1586364061
transform 1 0 22080 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_250
timestamp 1586364061
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_254
timestamp 1586364061
transform 1 0 24472 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_267
timestamp 1586364061
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_conb_1  _058_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_10
timestamp 1586364061
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_28
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_33_45
timestamp 1586364061
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_51
timestamp 1586364061
transform 1 0 5796 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_49
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_55
timestamp 1586364061
transform 1 0 6164 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5980 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6348 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_59
timestamp 1586364061
transform 1 0 6532 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_77
timestamp 1586364061
transform 1 0 8188 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_73
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_75
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_97
timestamp 1586364061
transform 1 0 10028 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_34_101
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_104
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 866 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_115
timestamp 1586364061
transform 1 0 11684 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_111
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_116
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_128
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_134
timestamp 1586364061
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_146
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_150
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _124_
timestamp 1586364061
transform 1 0 15456 0 -1 21216
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_22.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_20.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16652 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16008 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_174
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_178
timestamp 1586364061
transform 1 0 17480 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_160
timestamp 1586364061
transform 1 0 15824 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_164
timestamp 1586364061
transform 1 0 16192 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_168
timestamp 1586364061
transform 1 0 16560 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_188
timestamp 1586364061
transform 1 0 18400 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_187
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_buf_1  mux_top_track_20.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_192
timestamp 1586364061
transform 1 0 18768 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_192
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18952 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19136 0 -1 21216
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_205
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_205
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20148 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_209
timestamp 1586364061
transform 1 0 20332 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_211
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_34_224
timestamp 1586364061
transform 1 0 21712 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 21896 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_232
timestamp 1586364061
transform 1 0 22448 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_228
timestamp 1586364061
transform 1 0 22080 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 22264 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_237
timestamp 1586364061
transform 1 0 22908 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_234
timestamp 1586364061
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 22540 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_238
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  FILLER_34_245
timestamp 1586364061
transform 1 0 23644 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_241
timestamp 1586364061
transform 1 0 23276 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 23460 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_257
timestamp 1586364061
transform 1 0 24748 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_254
timestamp 1586364061
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23920 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_266
timestamp 1586364061
transform 1 0 25576 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_258
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 24932 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 25208 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_273
timestamp 1586364061
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_276
timestamp 1586364061
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_33_270
timestamp 1586364061
transform 1 0 25944 0 1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_261
timestamp 1586364061
transform 1 0 25116 0 -1 21216
box -38 -48 1142 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_14
timestamp 1586364061
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_18
timestamp 1586364061
transform 1 0 2760 0 1 21216
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 3312 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_43
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_79
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_83
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_97
timestamp 1586364061
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_101
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_127
timestamp 1586364061
transform 1 0 12788 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_151
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_155
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_158
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_18.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18952 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18768 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_189
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_213
timestamp 1586364061
transform 1 0 20700 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_217
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 21436 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 22632 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23828 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_240
timestamp 1586364061
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_256
timestamp 1586364061
transform 1 0 24656 0 1 21216
box -38 -48 406 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 25392 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 25944 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_262
timestamp 1586364061
transform 1 0 25208 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_268
timestamp 1586364061
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_272
timestamp 1586364061
transform 1 0 26128 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_276
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1564 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2576 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_14
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_18
timestamp 1586364061
transform 1 0 2760 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2944 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3312 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3680 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_22
timestamp 1586364061
transform 1 0 3128 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_26
timestamp 1586364061
transform 1 0 3496 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_30
timestamp 1586364061
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_41
timestamp 1586364061
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_46
timestamp 1586364061
transform 1 0 5336 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_50
timestamp 1586364061
transform 1 0 5704 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_54
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_75
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_79
timestamp 1586364061
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9844 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_83
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11408 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_104
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13340 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_131
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_135
timestamp 1586364061
transform 1 0 13524 0 -1 22304
box -38 -48 406 592
use scs8hd_buf_2  _122_
timestamp 1586364061
transform 1 0 15640 0 -1 22304
box -38 -48 406 592
use scs8hd_buf_2  _125_
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13892 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15456 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1586364061
transform 1 0 16744 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16192 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_162
timestamp 1586364061
transform 1 0 16008 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_20.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18124 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_179
timestamp 1586364061
transform 1 0 17572 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_183
timestamp 1586364061
transform 1 0 17940 0 -1 22304
box -38 -48 222 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_206
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_210
timestamp 1586364061
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_218
timestamp 1586364061
transform 1 0 21160 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21896 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 21436 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 22908 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_223
timestamp 1586364061
transform 1 0 21620 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_235
timestamp 1586364061
transform 1 0 22724 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23460 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24472 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23276 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_252
timestamp 1586364061
transform 1 0 24288 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_256
timestamp 1586364061
transform 1 0 24656 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 25024 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 24840 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 25576 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_264
timestamp 1586364061
transform 1 0 25392 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_268
timestamp 1586364061
transform 1 0 25760 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_16
timestamp 1586364061
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 3312 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_20
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_33
timestamp 1586364061
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_37
timestamp 1586364061
transform 1 0 4508 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4876 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_43
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7452 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_66
timestamp 1586364061
transform 1 0 7176 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_94
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_111
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_115
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_119
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12604 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_127
timestamp 1586364061
transform 1 0 12788 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_131
timestamp 1586364061
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_37_158
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_164
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _118_
timestamp 1586364061
transform 1 0 18308 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_191
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_195
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_37_199
timestamp 1586364061
transform 1 0 19412 0 1 22304
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_219
timestamp 1586364061
transform 1 0 21252 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_223
timestamp 1586364061
transform 1 0 21620 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 23276 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_243
timestamp 1586364061
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_254
timestamp 1586364061
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 25760 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_266
timestamp 1586364061
transform 1 0 25576 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_270
timestamp 1586364061
transform 1 0 25944 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_276
timestamp 1586364061
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 1840 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_10
timestamp 1586364061
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4232 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_36
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4876 0 -1 23392
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_38_40
timestamp 1586364061
transform 1 0 4784 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_60
timestamp 1586364061
transform 1 0 6624 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_71
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_88
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11500 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_106
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_110
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_132
timestamp 1586364061
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_136
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_2  _121_
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15456 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_149
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_158
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16008 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15824 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1586364061
transform 1 0 19228 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17940 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19044 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18676 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18308 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_181
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_185
timestamp 1586364061
transform 1 0 18124 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_189
timestamp 1586364061
transform 1 0 18492 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21068 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 20240 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_206
timestamp 1586364061
transform 1 0 20056 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_210
timestamp 1586364061
transform 1 0 20424 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 21436 0 -1 23392
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_38_219
timestamp 1586364061
transform 1 0 21252 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23920 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 23644 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_240
timestamp 1586364061
transform 1 0 23184 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_244
timestamp 1586364061
transform 1 0 23552 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_247
timestamp 1586364061
transform 1 0 23828 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_257
timestamp 1586364061
transform 1 0 24748 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_261
timestamp 1586364061
transform 1 0 25116 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_265
timestamp 1586364061
transform 1 0 25484 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_273
timestamp 1586364061
transform 1 0 26220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 1840 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_10
timestamp 1586364061
transform 1 0 2024 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3772 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3956 0 1 23392
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_40_45
timestamp 1586364061
transform 1 0 5244 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_41
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5428 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 5060 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_54
timestamp 1586364061
transform 1 0 6072 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_50
timestamp 1586364061
transform 1 0 5704 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6256 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5888 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5612 0 -1 24480
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_72
timestamp 1586364061
transform 1 0 7728 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_70
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7912 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _067_
timestamp 1586364061
transform 1 0 8096 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_88
timestamp 1586364061
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8648 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_96
timestamp 1586364061
transform 1 0 9936 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_90
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 10120 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_conb_1  _057_
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_113
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_117
timestamp 1586364061
transform 1 0 11868 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_100
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_113
timestamp 1586364061
transform 1 0 11500 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12604 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12236 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_6  FILLER_40_134
timestamp 1586364061
transform 1 0 13432 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_130
timestamp 1586364061
transform 1 0 13064 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13248 0 -1 24480
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12972 0 1 23392
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_148
timestamp 1586364061
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_149
timestamp 1586364061
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_152
timestamp 1586364061
transform 1 0 15088 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14904 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15456 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17204 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17020 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_167
timestamp 1586364061
transform 1 0 16468 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_6  FILLER_40_188
timestamp 1586364061
transform 1 0 18400 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_184
timestamp 1586364061
transform 1 0 18032 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18124 0 1 23392
box -38 -48 866 592
use scs8hd_fill_1  FILLER_40_194
timestamp 1586364061
transform 1 0 18952 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_194
timestamp 1586364061
transform 1 0 18952 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19044 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_206
timestamp 1586364061
transform 1 0 20056 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_206
timestamp 1586364061
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_199
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_210
timestamp 1586364061
transform 1 0 20424 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_210
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21528 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21344 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22540 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_234
timestamp 1586364061
transform 1 0 22632 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_219
timestamp 1586364061
transform 1 0 21252 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_231
timestamp 1586364061
transform 1 0 22356 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_235
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1586364061
transform 1 0 23276 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_254
timestamp 1586364061
transform 1 0 24472 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_250
timestamp 1586364061
transform 1 0 24104 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_254
timestamp 1586364061
transform 1 0 24472 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 24288 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_267
timestamp 1586364061
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_266
timestamp 1586364061
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_260
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1586364061
transform 1 0 24840 0 -1 24480
box -38 -48 866 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_270
timestamp 1586364061
transform 1 0 25944 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 26128 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1564 0 1 24480
box -38 -48 866 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2576 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_14
timestamp 1586364061
transform 1 0 2392 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_18
timestamp 1586364061
transform 1 0 2760 0 1 24480
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 3128 0 1 24480
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 2944 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 5612 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 5060 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 5428 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_41
timestamp 1586364061
transform 1 0 4876 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_45
timestamp 1586364061
transform 1 0 5244 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6900 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_41_72
timestamp 1586364061
transform 1 0 7728 0 1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_41_78
timestamp 1586364061
transform 1 0 8280 0 1 24480
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8556 0 1 24480
box -38 -48 1786 592
use scs8hd_buf_1  mux_top_track_18.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11316 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10948 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_100
timestamp 1586364061
transform 1 0 10304 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_105
timestamp 1586364061
transform 1 0 10764 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_109
timestamp 1586364061
transform 1 0 11132 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12972 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12788 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_138
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_142
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_146
timestamp 1586364061
transform 1 0 14536 0 1 24480
box -38 -48 314 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 16560 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16008 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 16376 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17112 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 17480 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_160
timestamp 1586364061
transform 1 0 15824 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_164
timestamp 1586364061
transform 1 0 16192 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_172
timestamp 1586364061
transform 1 0 16928 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_176
timestamp 1586364061
transform 1 0 17296 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _117_
timestamp 1586364061
transform 1 0 19044 0 1 24480
box -38 -48 406 592
use scs8hd_buf_1  mux_top_track_22.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 18492 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_180
timestamp 1586364061
transform 1 0 17664 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_187
timestamp 1586364061
transform 1 0 18308 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_191
timestamp 1586364061
transform 1 0 18676 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20148 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19964 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_199
timestamp 1586364061
transform 1 0 19412 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_203
timestamp 1586364061
transform 1 0 19780 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_216
timestamp 1586364061
transform 1 0 20976 0 1 24480
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21988 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21804 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 21436 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_223
timestamp 1586364061
transform 1 0 21620 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_236
timestamp 1586364061
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 24656 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_240
timestamp 1586364061
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_254
timestamp 1586364061
transform 1 0 24472 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 25208 0 1 24480
box -38 -48 406 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 25760 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 25024 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_258
timestamp 1586364061
transform 1 0 24840 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_266
timestamp 1586364061
transform 1 0 25576 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_270
timestamp 1586364061
transform 1 0 25944 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_276
timestamp 1586364061
transform 1 0 26496 0 1 24480
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 25568
box -38 -48 866 592
use scs8hd_buf_1  mux_left_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2208 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_6
timestamp 1586364061
transform 1 0 1656 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_10
timestamp 1586364061
transform 1 0 2024 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1586364061
transform 1 0 4324 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 5612 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5980 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6348 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_48
timestamp 1586364061
transform 1 0 5520 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_51
timestamp 1586364061
transform 1 0 5796 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_55
timestamp 1586364061
transform 1 0 6164 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_59
timestamp 1586364061
transform 1 0 6532 0 -1 25568
box -38 -48 314 592
use scs8hd_buf_2  _066_
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8096 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7452 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 7820 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_67
timestamp 1586364061
transform 1 0 7268 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_71
timestamp 1586364061
transform 1 0 7636 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 130 592
use scs8hd_buf_1  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9936 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_85
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_89
timestamp 1586364061
transform 1 0 9292 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_99
timestamp 1586364061
transform 1 0 10212 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10948 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10396 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_103
timestamp 1586364061
transform 1 0 10580 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_116
timestamp 1586364061
transform 1 0 11776 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_120
timestamp 1586364061
transform 1 0 12144 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_134
timestamp 1586364061
transform 1 0 13432 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _123_
timestamp 1586364061
transform 1 0 14260 0 -1 25568
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_142
timestamp 1586364061
transform 1 0 14168 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_147
timestamp 1586364061
transform 1 0 14628 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_153
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _120_
timestamp 1586364061
transform 1 0 17112 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_165
timestamp 1586364061
transform 1 0 16284 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_170
timestamp 1586364061
transform 1 0 16744 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_6  FILLER_42_178
timestamp 1586364061
transform 1 0 17480 0 -1 25568
box -38 -48 590 592
use scs8hd_buf_2  _119_
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_191
timestamp 1586364061
transform 1 0 18676 0 -1 25568
box -38 -48 1142 592
use scs8hd_buf_2  _116_
timestamp 1586364061
transform 1 0 19964 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_203
timestamp 1586364061
transform 1 0 19780 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_209
timestamp 1586364061
transform 1 0 20332 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_213
timestamp 1586364061
transform 1 0 20700 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_4  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 22816 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 21712 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 21528 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 22632 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_228
timestamp 1586364061
transform 1 0 22080 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_232
timestamp 1586364061
transform 1 0 22448 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 23644 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_240
timestamp 1586364061
transform 1 0 23184 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_244
timestamp 1586364061
transform 1 0 23552 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_247
timestamp 1586364061
transform 1 0 23828 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_253
timestamp 1586364061
transform 1 0 24380 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_265
timestamp 1586364061
transform 1 0 25484 0 -1 25568
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 13910 0 13966 480 6 ccff_head
port 0 nsew default input
rlabel metal2 s 23202 0 23258 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 1912 480 2032 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 21904 480 22024 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 15648 480 15768 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 27520 824 28000 944 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 27520 4224 28000 4344 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 27520 20816 28000 20936 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 27520 21904 28000 22024 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 27520 15104 28000 15224 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 27520 15648 28000 15768 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 27520 16736 28000 16856 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal2 s 4894 27520 4950 28000 6 chany_top_in[0]
port 82 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_in[10]
port 83 nsew default input
rlabel metal2 s 11334 27520 11390 28000 6 chany_top_in[11]
port 84 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[12]
port 85 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[13]
port 86 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[14]
port 87 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[15]
port 88 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[16]
port 89 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[17]
port 90 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[18]
port 91 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_in[19]
port 92 nsew default input
rlabel metal2 s 5538 27520 5594 28000 6 chany_top_in[1]
port 93 nsew default input
rlabel metal2 s 6090 27520 6146 28000 6 chany_top_in[2]
port 94 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[3]
port 95 nsew default input
rlabel metal2 s 7286 27520 7342 28000 6 chany_top_in[4]
port 96 nsew default input
rlabel metal2 s 7838 27520 7894 28000 6 chany_top_in[5]
port 97 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[6]
port 98 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[7]
port 99 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chany_top_in[8]
port 100 nsew default input
rlabel metal2 s 10138 27520 10194 28000 6 chany_top_in[9]
port 101 nsew default input
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[0]
port 102 nsew default tristate
rlabel metal2 s 22374 27520 22430 28000 6 chany_top_out[10]
port 103 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[11]
port 104 nsew default tristate
rlabel metal2 s 23570 27520 23626 28000 6 chany_top_out[12]
port 105 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[13]
port 106 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[14]
port 107 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[15]
port 108 nsew default tristate
rlabel metal2 s 25870 27520 25926 28000 6 chany_top_out[16]
port 109 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[17]
port 110 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[18]
port 111 nsew default tristate
rlabel metal2 s 27618 27520 27674 28000 6 chany_top_out[19]
port 112 nsew default tristate
rlabel metal2 s 17130 27520 17186 28000 6 chany_top_out[1]
port 113 nsew default tristate
rlabel metal2 s 17774 27520 17830 28000 6 chany_top_out[2]
port 114 nsew default tristate
rlabel metal2 s 18326 27520 18382 28000 6 chany_top_out[3]
port 115 nsew default tristate
rlabel metal2 s 18878 27520 18934 28000 6 chany_top_out[4]
port 116 nsew default tristate
rlabel metal2 s 19522 27520 19578 28000 6 chany_top_out[5]
port 117 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[6]
port 118 nsew default tristate
rlabel metal2 s 20626 27520 20682 28000 6 chany_top_out[7]
port 119 nsew default tristate
rlabel metal2 s 21270 27520 21326 28000 6 chany_top_out[8]
port 120 nsew default tristate
rlabel metal2 s 21822 27520 21878 28000 6 chany_top_out[9]
port 121 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 122 nsew default input
rlabel metal3 s 0 23672 480 23792 6 left_top_grid_pin_42_
port 123 nsew default input
rlabel metal3 s 0 24216 480 24336 6 left_top_grid_pin_43_
port 124 nsew default input
rlabel metal3 s 0 24760 480 24880 6 left_top_grid_pin_44_
port 125 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_45_
port 126 nsew default input
rlabel metal3 s 0 25984 480 26104 6 left_top_grid_pin_46_
port 127 nsew default input
rlabel metal3 s 0 26528 480 26648 6 left_top_grid_pin_47_
port 128 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_48_
port 129 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_49_
port 130 nsew default input
rlabel metal2 s 4618 0 4674 480 6 prog_clk
port 131 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_1_
port 132 nsew default input
rlabel metal3 s 27520 23672 28000 23792 6 right_top_grid_pin_42_
port 133 nsew default input
rlabel metal3 s 27520 24216 28000 24336 6 right_top_grid_pin_43_
port 134 nsew default input
rlabel metal3 s 27520 24760 28000 24880 6 right_top_grid_pin_44_
port 135 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_top_grid_pin_45_
port 136 nsew default input
rlabel metal3 s 27520 25984 28000 26104 6 right_top_grid_pin_46_
port 137 nsew default input
rlabel metal3 s 27520 26528 28000 26648 6 right_top_grid_pin_47_
port 138 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_top_grid_pin_48_
port 139 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_49_
port 140 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_34_
port 141 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_35_
port 142 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_36_
port 143 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 top_left_grid_pin_37_
port 144 nsew default input
rlabel metal2 s 2594 27520 2650 28000 6 top_left_grid_pin_38_
port 145 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_39_
port 146 nsew default input
rlabel metal2 s 3790 27520 3846 28000 6 top_left_grid_pin_40_
port 147 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 top_left_grid_pin_41_
port 148 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 149 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
