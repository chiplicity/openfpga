* NGSPICE file created from sb_1__8_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt sb_1__8_ bottom_left_grid_pin_42_ bottom_left_grid_pin_43_ bottom_left_grid_pin_44_
+ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_ bottom_left_grid_pin_48_
+ bottom_left_grid_pin_49_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ left_top_grid_pin_1_ prog_clk right_bottom_grid_pin_34_
+ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_
+ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ right_top_grid_pin_1_
+ VPWR VGND
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_0.mux_l4_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_9.mux_l4_in_0_/S mux_left_track_17.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_3.mux_l1_in_3_/S mux_bottom_track_3.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_062_ chanx_right_in[12] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_114_ _114_/A chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l3_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_0_ bottom_left_grid_pin_46_ chanx_right_in[13] mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_028_ _028_/HI _028_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X _114_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[4] mux_bottom_track_3.mux_l1_in_3_/S
+ mux_bottom_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_061_ chanx_right_in[13] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_4.mux_l4_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X _071_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_113_ _113_/A chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l2_in_1_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_3_ _042_/HI chanx_left_in[16] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X _063_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_3.mux_l2_in_0_/S
+ mux_bottom_track_3.mux_l3_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S mux_right_track_8.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_060_ chanx_right_in[14] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_112_ _112_/A chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_1_/S mux_right_track_8.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_23.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_2_ chanx_left_in[6] chany_bottom_in[16] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_3.mux_l1_in_3_/S
+ mux_bottom_track_3.mux_l2_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_9.mux_l2_in_1_/S
+ mux_bottom_track_9.mux_l3_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_111_ _111_/A chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_1_/S mux_right_track_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_1_ chany_bottom_in[9] chany_bottom_in[2] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_1.mux_l3_in_0_/S
+ mux_bottom_track_3.mux_l1_in_3_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_11.mux_l2_in_1_/S
+ mux_bottom_track_11.mux_l3_in_0_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l2_in_1_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_110_ _110_/A chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_11.mux_l3_in_0_/X
+ _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_0_ right_bottom_grid_pin_41_ mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l2_in_1_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_7.mux_l3_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_13.mux_l2_in_0_ mux_bottom_track_13.mux_l1_in_1_/X mux_bottom_track_13.mux_l1_in_0_/X
+ mux_bottom_track_13.mux_l2_in_0_/S mux_bottom_track_13.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S mux_bottom_track_25.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_9.mux_l3_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_8.mux_l1_in_0_ right_bottom_grid_pin_37_ right_top_grid_pin_1_ mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_2_0_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_27.mux_l2_in_0_/X
+ _102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X _091_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_25.mux_l2_in_1_ _051_/HI chanx_left_in[18] mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_13.mux_l1_in_1_ _045_/HI chanx_left_in[10] mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S mux_bottom_track_9.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l2_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_099_ chanx_right_in[3] chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l2_in_1_ _028_/HI chanx_left_in[15] mux_bottom_track_9.mux_l2_in_1_/S
+ mux_bottom_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X _079_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_6_ chanx_left_in[14] chanx_left_in[5] mux_right_track_4.mux_l1_in_4_/S
+ mux_right_track_4.mux_l1_in_6_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_3.mux_l2_in_3_ _032_/HI left_bottom_grid_pin_40_ mux_left_track_3.mux_l2_in_1_/S
+ mux_left_track_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_13.mux_l1_in_0_ bottom_left_grid_pin_44_ chanx_right_in[10] mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l2_in_0_ bottom_left_grid_pin_42_ mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S mux_bottom_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_15.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_098_ chanx_right_in[1] chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S mux_left_track_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_0_ chanx_left_in[8] mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_1_/S mux_bottom_track_9.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_4.mux_l1_in_5_ chany_bottom_in[17] chany_bottom_in[10] mux_right_track_4.mux_l1_in_4_/S
+ mux_right_track_4.mux_l1_in_5_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l4_in_0_/X _073_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l2_in_2_ left_bottom_grid_pin_38_ left_bottom_grid_pin_36_ mux_left_track_3.mux_l2_in_1_/S
+ mux_left_track_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_1.mux_l2_in_1_/S mux_left_track_1.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l2_in_3_ _041_/HI mux_right_track_4.mux_l1_in_6_/X mux_right_track_4.mux_l2_in_2_/S
+ mux_right_track_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_097_ chanx_right_in[0] chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l1_in_0_ chanx_right_in[19] chanx_right_in[18] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_4_ chany_bottom_in[3] right_bottom_grid_pin_41_ mux_right_track_4.mux_l1_in_4_/S
+ mux_right_track_4.mux_l1_in_4_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l1_in_0_ bottom_left_grid_pin_42_ chanx_right_in[8] mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S mux_right_track_4.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X _111_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_1.mux_l1_in_1_/S mux_left_track_1.mux_l2_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_1_ left_bottom_grid_pin_34_ chany_bottom_in[14] mux_left_track_3.mux_l2_in_1_/S
+ mux_left_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_1_/S mux_right_track_4.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_4.mux_l3_in_1_/S mux_right_track_4.mux_l4_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l2_in_2_ mux_right_track_4.mux_l1_in_5_/X mux_right_track_4.mux_l1_in_4_/X
+ mux_right_track_4.mux_l2_in_2_/S mux_right_track_4.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_096_ chanx_left_in[0] chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_079_ _079_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_16.mux_l1_in_3_ _037_/HI chanx_left_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_3_ right_bottom_grid_pin_40_ right_bottom_grid_pin_39_
+ mux_right_track_4.mux_l1_in_4_/S mux_right_track_4.mux_l1_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_27.mux_l2_in_0_/S mux_left_track_1.mux_l1_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_1_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_4.mux_l2_in_2_/S mux_right_track_4.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l1_in_1_ chany_bottom_in[7] chany_bottom_in[0] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_095_ _095_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_2_/S mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_078_ chanx_left_in[16] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.mux_l1_in_2_ chanx_left_in[8] chany_bottom_in[15] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_38_ right_bottom_grid_pin_37_
+ mux_right_track_4.mux_l1_in_4_/S mux_right_track_4.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_4.mux_l1_in_4_/S mux_right_track_4.mux_l2_in_2_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l1_in_0_ chanx_right_in[13] chanx_right_in[4] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_094_ _094_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_2_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_077_ chanx_left_in[17] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_1_ chany_bottom_in[8] chany_bottom_in[1] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_36_ right_bottom_grid_pin_35_
+ mux_right_track_4.mux_l1_in_4_/S mux_right_track_4.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_2.mux_l4_in_0_/S mux_right_track_4.mux_l1_in_4_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_093_ _093_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l2_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
Xmux_bottom_track_5.mux_l1_in_3_ _054_/HI chanx_left_in[7] mux_bottom_track_5.mux_l1_in_2_/S
+ mux_bottom_track_5.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_076_ chanx_left_in[18] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_23.mux_l2_in_0_/X
+ _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_0_ right_bottom_grid_pin_38_ right_bottom_grid_pin_34_
+ mux_right_track_16.mux_l1_in_3_/S mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_0_ right_bottom_grid_pin_34_ right_top_grid_pin_1_ mux_right_track_4.mux_l1_in_4_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l4_in_0_/X _093_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ _059_/A chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l2_in_0_/X
+ _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_092_ chanx_left_in[2] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_19.mux_l2_in_0_/S
+ mux_bottom_track_21.mux_l1_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l1_in_2_ chanx_left_in[5] bottom_left_grid_pin_48_ mux_bottom_track_5.mux_l1_in_2_/S
+ mux_bottom_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_075_ _075_/A chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X _087_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_058_ chanx_right_in[16] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_19.mux_l2_in_0_ mux_bottom_track_19.mux_l1_in_1_/X mux_bottom_track_19.mux_l1_in_0_/X
+ mux_bottom_track_19.mux_l2_in_0_/S mux_bottom_track_19.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_21.mux_l2_in_0_ mux_bottom_track_21.mux_l1_in_1_/X mux_bottom_track_21.mux_l1_in_0_/X
+ mux_bottom_track_21.mux_l2_in_0_/S mux_bottom_track_21.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_19.mux_l1_in_1_ _048_/HI chanx_left_in[14] mux_bottom_track_19.mux_l1_in_0_/S
+ mux_bottom_track_19.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_21.mux_l1_in_1_ _049_/HI chanx_left_in[16] mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X _075_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_5.mux_l2_in_1_/S
+ mux_bottom_track_5.mux_l3_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_091_ _091_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_074_ _074_/A chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_46_ bottom_left_grid_pin_44_
+ mux_bottom_track_5.mux_l1_in_2_/S mux_bottom_track_5.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_057_ chanx_right_in[17] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_25.mux_l3_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_9.mux_l2_in_3_ _035_/HI left_bottom_grid_pin_41_ mux_left_track_9.mux_l2_in_2_/S
+ mux_left_track_9.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_109_ _109_/A chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_3_ _036_/HI chanx_left_in[12] mux_right_track_0.mux_l2_in_3_/S
+ mux_right_track_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_19.mux_l1_in_0_ bottom_left_grid_pin_47_ chanx_right_in[14] mux_bottom_track_19.mux_l1_in_0_/S
+ mux_bottom_track_19.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_21.mux_l1_in_0_ bottom_left_grid_pin_48_ chanx_right_in[16] mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_5.mux_l1_in_2_/S
+ mux_bottom_track_5.mux_l2_in_1_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S mux_left_track_9.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_090_ chanx_left_in[4] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X _113_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S mux_right_track_0.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_42_ chanx_right_in[5] mux_bottom_track_5.mux_l1_in_2_/S
+ mux_bottom_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_073_ _073_/A chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_056_ chanx_right_in[18] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_3_ _030_/HI left_bottom_grid_pin_38_ mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_108_ _108_/A chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l2_in_2_ left_bottom_grid_pin_37_ left_top_grid_pin_1_ mux_left_track_9.mux_l2_in_2_/S
+ mux_left_track_9.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_2_ chanx_left_in[2] chany_bottom_in[19] mux_right_track_0.mux_l2_in_3_/S
+ mux_right_track_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X _059_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_3.mux_l3_in_0_/S
+ mux_bottom_track_5.mux_l1_in_2_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S mux_left_track_17.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ chanx_right_in[2] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l1_in_2_ left_bottom_grid_pin_34_ chany_bottom_in[17] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_107_ _107_/A chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l2_in_1_ chany_bottom_in[16] chany_bottom_in[9] mux_left_track_9.mux_l2_in_2_/S
+ mux_left_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_0.mux_l2_in_1_ chany_bottom_in[12] mux_right_track_0.mux_l1_in_2_/X
+ mux_right_track_0.mux_l2_in_3_/S mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l1_in_2_ chany_bottom_in[5] right_bottom_grid_pin_41_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l2_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_071_ _071_/A chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l1_in_3_ _039_/HI chanx_left_in[18] mux_right_track_24.mux_l1_in_3_/S
+ mux_right_track_24.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_17.mux_l1_in_1_ chany_bottom_in[10] chany_bottom_in[3] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_106_ _106_/A chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_9.mux_l2_in_0_ chany_bottom_in[2] mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_2_/S mux_left_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_3_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_39_ right_bottom_grid_pin_37_
+ mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l1_in_3_/X mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_1_/S mux_right_track_24.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_11.mux_l3_in_0_/S
+ mux_bottom_track_13.mux_l1_in_1_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_070_ chanx_right_in[4] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.mux_l1_in_2_ chanx_left_in[9] chany_bottom_in[14] mux_right_track_24.mux_l1_in_3_/S
+ mux_right_track_24.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_19.mux_l1_in_0_/S
+ mux_bottom_track_19.mux_l2_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l3_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_105_ _105_/A chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ chanx_right_in[17] chanx_right_in[8] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X _095_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_3_ _043_/HI chanx_left_in[2] mux_bottom_track_1.mux_l1_in_3_/S
+ mux_bottom_track_1.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l1_in_0_ chanx_right_in[16] chanx_right_in[6] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_35_ right_top_grid_pin_1_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_13.mux_l2_in_0_/X
+ _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_1_/S mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.mux_l1_in_1_ chany_bottom_in[7] chany_bottom_in[0] mux_right_track_24.mux_l1_in_3_/S
+ mux_right_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_1.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_19.mux_l1_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_6_ left_bottom_grid_pin_41_ left_bottom_grid_pin_40_ mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_6_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_104_ _104_/A chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l1_in_3_/X mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_1_/S mux_bottom_track_1.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_1.mux_l1_in_2_ chanx_left_in[1] bottom_left_grid_pin_48_ mux_bottom_track_1.mux_l1_in_3_/S
+ mux_bottom_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l3_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_15.mux_l2_in_0_ mux_bottom_track_15.mux_l1_in_1_/X mux_bottom_track_15.mux_l1_in_0_/X
+ mux_bottom_track_15.mux_l2_in_0_/S mux_bottom_track_15.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_39_ right_bottom_grid_pin_35_
+ mux_right_track_24.mux_l1_in_3_/S mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_24.mux_l3_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_15.mux_l1_in_1_ _046_/HI chanx_left_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_5_ left_bottom_grid_pin_39_ left_bottom_grid_pin_38_ mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_5_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_034_ _034_/HI _034_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S mux_bottom_track_1.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_103_ _103_/A chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_46_ bottom_left_grid_pin_44_
+ mux_bottom_track_1.mux_l1_in_3_/S mux_bottom_track_1.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_0.mux_l2_in_3_/S mux_right_track_0.mux_l3_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_3.mux_l1_in_0_/S mux_left_track_3.mux_l2_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_5.mux_l2_in_3_ _034_/HI mux_left_track_5.mux_l1_in_6_/X mux_left_track_5.mux_l2_in_1_/S
+ mux_left_track_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_15.mux_l1_in_0_ bottom_left_grid_pin_45_ chanx_right_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_9.mux_l2_in_2_/S mux_left_track_9.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_27.mux_l2_in_0_ _052_/HI mux_bottom_track_27.mux_l1_in_0_/X mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_033_ _033_/HI _033_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X _115_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_102_ _102_/A chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l1_in_4_ left_bottom_grid_pin_37_ left_bottom_grid_pin_36_ mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_4_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S mux_left_track_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_42_ chanx_right_in[2] mux_bottom_track_1.mux_l1_in_3_/S
+ mux_bottom_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l2_in_3_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_1_/S mux_left_track_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_1.mux_l4_in_0_/S mux_left_track_3.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.mux_l2_in_2_ mux_left_track_5.mux_l1_in_5_/X mux_left_track_5.mux_l1_in_4_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_2_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_2_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_032_ _032_/HI _032_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_101_ chanx_right_in[11] chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l1_in_3_ left_bottom_grid_pin_35_ left_bottom_grid_pin_34_ mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_27.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[15] mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X _067_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_right_track_0.mux_l1_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_1_/S mux_left_track_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_24.mux_l2_in_1_/S
+ mux_right_track_24.mux_l3_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_5.mux_l4_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_031_ _031_/HI _031_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ chanx_right_in[7] chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l1_in_3_ _031_/HI left_bottom_grid_pin_39_ mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l1_in_2_ left_top_grid_pin_1_ chany_bottom_in[15] mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_33.mux_l2_in_0_/S ccff_tail
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_24.mux_l1_in_3_/S
+ mux_right_track_24.mux_l2_in_1_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l2_in_1_ mux_left_track_25.mux_l1_in_3_/X mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l2_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_030_ _030_/HI _030_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_5.mux_l1_in_1_ chany_bottom_in[8] chany_bottom_in[1] mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_2_ left_bottom_grid_pin_35_ chany_bottom_in[18] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l2_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_1.mux_l2_in_1_/S
+ mux_bottom_track_1.mux_l3_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_16.mux_l3_in_0_/S
+ mux_right_track_24.mux_l1_in_3_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_21.mux_l2_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_11.mux_l3_in_0_ mux_bottom_track_11.mux_l2_in_1_/X mux_bottom_track_11.mux_l2_in_0_/X
+ mux_bottom_track_11.mux_l3_in_0_/S mux_bottom_track_11.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l1_in_0_ chanx_right_in[14] chanx_right_in[5] mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_089_ chanx_left_in[5] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l1_in_1_ chany_bottom_in[11] chany_bottom_in[4] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_25.mux_l3_in_0_/S mux_left_track_33.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S mux_right_track_32.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_11.mux_l2_in_1_ _044_/HI chanx_left_in[19] mux_bottom_track_11.mux_l2_in_1_/S
+ mux_bottom_track_11.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_1.mux_l1_in_3_/S
+ mux_bottom_track_1.mux_l2_in_1_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_prog_clk clkbuf_2_3_0_prog_clk/X clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_32.mux_l2_in_1_ _040_/HI chanx_left_in[10] mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_7.mux_l2_in_1_/S
+ mux_bottom_track_7.mux_l3_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_088_ chanx_left_in[6] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_25.mux_l1_in_0_ chanx_right_in[18] chanx_right_in[9] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_11.mux_l2_in_0_ chanx_left_in[9] mux_bottom_track_11.mux_l1_in_0_/X
+ mux_bottom_track_11.mux_l2_in_1_/S mux_bottom_track_11.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_7.mux_l1_in_3_ _055_/HI chanx_left_in[11] mux_bottom_track_7.mux_l1_in_3_/S
+ mux_bottom_track_7.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_32.mux_l3_in_0_/S
+ mux_bottom_track_1.mux_l1_in_3_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_7.mux_l3_in_0_ mux_bottom_track_7.mux_l2_in_1_/X mux_bottom_track_7.mux_l2_in_0_/X
+ mux_bottom_track_7.mux_l3_in_0_/S mux_bottom_track_7.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_19.mux_l2_in_0_/X
+ _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_7.mux_l1_in_3_/S
+ mux_bottom_track_7.mux_l2_in_1_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_32.mux_l1_in_1_ chany_bottom_in[13] chany_bottom_in[6] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l2_in_1_ mux_bottom_track_7.mux_l1_in_3_/X mux_bottom_track_7.mux_l1_in_2_/X
+ mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_087_ _087_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _083_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_7.mux_l1_in_2_ chanx_left_in[6] bottom_left_grid_pin_49_ mux_bottom_track_7.mux_l1_in_3_/S
+ mux_bottom_track_7.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_3_ _029_/HI left_bottom_grid_pin_41_ mux_left_track_1.mux_l2_in_1_/S
+ mux_left_track_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_11.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[9] mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_23.mux_l2_in_0_ mux_bottom_track_23.mux_l1_in_1_/X mux_bottom_track_23.mux_l1_in_0_/X
+ mux_bottom_track_23.mux_l2_in_0_/S mux_bottom_track_23.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_16.mux_l2_in_1_/S
+ mux_right_track_16.mux_l3_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_5.mux_l3_in_0_/S
+ mux_bottom_track_7.mux_l1_in_3_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_32.mux_l1_in_0_ right_bottom_grid_pin_40_ right_bottom_grid_pin_36_
+ mux_right_track_32.mux_l1_in_0_/S mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_23.mux_l1_in_1_ _050_/HI chanx_left_in[17] mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S mux_left_track_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l2_in_0_ mux_bottom_track_7.mux_l1_in_1_/X mux_bottom_track_7.mux_l1_in_0_/X
+ mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_086_ chanx_left_in[8] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X _074_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l3_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_069_ chanx_right_in[5] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_7.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_7.mux_l1_in_3_/S mux_bottom_track_7.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l2_in_2_ left_bottom_grid_pin_39_ left_bottom_grid_pin_37_ mux_left_track_1.mux_l2_in_1_/S
+ mux_left_track_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l2_in_1_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_prog_clk clkbuf_2_3_0_prog_clk/X clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_2.mux_l2_in_3_ _038_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_3_/S
+ mux_right_track_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_23.mux_l1_in_0_ bottom_left_grid_pin_49_ chanx_right_in[17] mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l2_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_085_ chanx_left_in[9] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_25.mux_l1_in_0_/S mux_left_track_25.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_068_ chanx_right_in[6] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_7.mux_l3_in_0_/X _112_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S mux_right_track_2.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_7.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[6] mux_bottom_track_7.mux_l1_in_3_/S
+ mux_bottom_track_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_1_ left_bottom_grid_pin_35_ left_top_grid_pin_1_ mux_left_track_1.mux_l2_in_1_/S
+ mux_left_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_1_/S mux_right_track_2.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_8.mux_l4_in_0_/S mux_right_track_16.mux_l1_in_3_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] chany_bottom_in[18] mux_right_track_2.mux_l2_in_3_/S
+ mux_right_track_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_13.mux_l2_in_0_/S
+ mux_bottom_track_15.mux_l1_in_1_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_17.mux_l3_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_084_ chanx_left_in[10] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_067_ _067_/A chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_1_/S mux_left_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_1_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_0 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l1_in_1_ chany_bottom_in[13] chany_bottom_in[6] mux_left_track_1.mux_l1_in_1_/S
+ mux_left_track_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l2_in_1_ chany_bottom_in[11] chany_bottom_in[4] mux_right_track_2.mux_l2_in_3_/S
+ mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_083_ _083_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_5.mux_l3_in_1_/S mux_left_track_5.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_066_ chanx_right_in[8] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_2_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_2_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail mux_left_track_33.mux_l3_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l1_in_0_ chanx_right_in[12] chanx_right_in[2] mux_left_track_1.mux_l1_in_1_/S
+ mux_left_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_1_ _033_/HI mux_left_track_33.mux_l1_in_2_/X mux_left_track_33.mux_l2_in_0_/S
+ mux_left_track_33.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_3_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_2.mux_l3_in_1_/S mux_right_track_2.mux_l4_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_082_ chanx_left_in[12] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l3_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_33.mux_l1_in_2_ left_bottom_grid_pin_40_ left_bottom_grid_pin_36_
+ mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ chanx_right_in[9] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_21_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_0_/S mux_left_track_33.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_21.mux_l2_in_0_/X
+ _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_2.mux_l2_in_3_/S mux_right_track_2.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_3.mux_l1_in_3_ _053_/HI chanx_left_in[4] mux_bottom_track_3.mux_l1_in_3_/S
+ mux_bottom_track_3.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_081_ chanx_left_in[13] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X _094_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_5.mux_l1_in_4_/S mux_left_track_5.mux_l2_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_33.mux_l1_in_1_ chany_bottom_in[19] chany_bottom_in[12] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l1_in_0_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_15.mux_l2_in_0_/X
+ _108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_064_ chanx_right_in[10] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_8.mux_l3_in_1_/S mux_right_track_8.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l1_in_3_/X mux_bottom_track_3.mux_l1_in_2_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_3_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_17.mux_l1_in_0_/S mux_left_track_17.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_2_ chanx_left_in[3] bottom_left_grid_pin_49_ mux_bottom_track_3.mux_l1_in_3_/S
+ mux_bottom_track_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_080_ chanx_left_in[14] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_3.mux_l4_in_0_/S mux_left_track_5.mux_l1_in_4_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l1_in_0_ chany_bottom_in[5] chanx_right_in[10] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_063_ _063_/A chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_0_/S mux_bottom_track_17.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l3_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_115_ _115_/A chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l1_in_1_ _047_/HI chanx_left_in[13] mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_029_ _029_/HI _029_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

