magic
tech sky130A
magscale 1 2
timestamp 1605120382
<< locali >>
rect 9045 16983 9079 17153
rect 6377 14875 6411 15113
rect 9137 14943 9171 15113
rect 17693 14875 17727 15045
rect 21683 13685 21741 13719
rect 11253 10523 11287 10625
<< viali >>
rect 21373 20553 21407 20587
rect 25789 20349 25823 20383
rect 25973 20213 26007 20247
rect 26433 20213 26467 20247
rect 2053 19125 2087 19159
rect 2329 19125 2363 19159
rect 2421 18853 2455 18887
rect 1869 18785 1903 18819
rect 2329 18785 2363 18819
rect 10129 18785 10163 18819
rect 18880 18785 18914 18819
rect 22273 18785 22307 18819
rect 24492 18785 24526 18819
rect 2605 18717 2639 18751
rect 9873 18717 9907 18751
rect 18613 18717 18647 18751
rect 22017 18717 22051 18751
rect 24225 18717 24259 18751
rect 8217 18649 8251 18683
rect 23397 18649 23431 18683
rect 1961 18581 1995 18615
rect 11253 18581 11287 18615
rect 12633 18581 12667 18615
rect 15117 18581 15151 18615
rect 19993 18581 20027 18615
rect 21097 18581 21131 18615
rect 25605 18581 25639 18615
rect 20913 18377 20947 18411
rect 3525 18309 3559 18343
rect 14013 18309 14047 18343
rect 20453 18309 20487 18343
rect 2605 18241 2639 18275
rect 3617 18241 3651 18275
rect 12633 18241 12667 18275
rect 15577 18241 15611 18275
rect 19165 18241 19199 18275
rect 19625 18241 19659 18275
rect 19993 18241 20027 18275
rect 21097 18241 21131 18275
rect 24317 18241 24351 18275
rect 2513 18173 2547 18207
rect 8125 18173 8159 18207
rect 12889 18173 12923 18207
rect 18981 18173 19015 18207
rect 21353 18173 21387 18207
rect 25237 18173 25271 18207
rect 1961 18105 1995 18139
rect 8033 18105 8067 18139
rect 8370 18105 8404 18139
rect 10241 18105 10275 18139
rect 12173 18105 12207 18139
rect 14933 18105 14967 18139
rect 15485 18105 15519 18139
rect 19073 18105 19107 18139
rect 25482 18105 25516 18139
rect 2053 18037 2087 18071
rect 2421 18037 2455 18071
rect 3065 18037 3099 18071
rect 9505 18037 9539 18071
rect 9873 18037 9907 18071
rect 15025 18037 15059 18071
rect 15393 18037 15427 18071
rect 17785 18037 17819 18071
rect 18429 18037 18463 18071
rect 18613 18037 18647 18071
rect 22477 18037 22511 18071
rect 22753 18037 22787 18071
rect 24593 18037 24627 18071
rect 25145 18037 25179 18071
rect 26617 18037 26651 18071
rect 13001 17833 13035 17867
rect 14381 17833 14415 17867
rect 18613 17833 18647 17867
rect 21281 17833 21315 17867
rect 25237 17833 25271 17867
rect 26525 17833 26559 17867
rect 19073 17765 19107 17799
rect 1941 17697 1975 17731
rect 4885 17697 4919 17731
rect 7021 17697 7055 17731
rect 8401 17697 8435 17731
rect 11877 17697 11911 17731
rect 15557 17697 15591 17731
rect 18981 17697 19015 17731
rect 26893 17697 26927 17731
rect 1685 17629 1719 17663
rect 4629 17629 4663 17663
rect 8493 17629 8527 17663
rect 8585 17629 8619 17663
rect 11621 17629 11655 17663
rect 15301 17629 15335 17663
rect 17601 17629 17635 17663
rect 19257 17629 19291 17663
rect 21373 17629 21407 17663
rect 21557 17629 21591 17663
rect 25329 17629 25363 17663
rect 25513 17629 25547 17663
rect 26985 17629 27019 17663
rect 27077 17629 27111 17663
rect 18521 17561 18555 17595
rect 22109 17561 22143 17595
rect 25881 17561 25915 17595
rect 3065 17493 3099 17527
rect 6009 17493 6043 17527
rect 8033 17493 8067 17527
rect 9045 17493 9079 17527
rect 10057 17493 10091 17527
rect 10333 17493 10367 17527
rect 15117 17493 15151 17527
rect 16681 17493 16715 17527
rect 20913 17493 20947 17527
rect 24869 17493 24903 17527
rect 3801 17289 3835 17323
rect 4445 17289 4479 17323
rect 7757 17289 7791 17323
rect 11989 17289 12023 17323
rect 17877 17289 17911 17323
rect 18429 17289 18463 17323
rect 19533 17289 19567 17323
rect 20361 17289 20395 17323
rect 20913 17289 20947 17323
rect 22293 17289 22327 17323
rect 22661 17289 22695 17323
rect 24225 17289 24259 17323
rect 24593 17289 24627 17323
rect 25789 17289 25823 17323
rect 3065 17221 3099 17255
rect 5917 17221 5951 17255
rect 7389 17221 7423 17255
rect 9873 17221 9907 17255
rect 11621 17221 11655 17255
rect 14289 17221 14323 17255
rect 20821 17221 20855 17255
rect 24961 17221 24995 17255
rect 26801 17221 26835 17255
rect 2513 17153 2547 17187
rect 2697 17153 2731 17187
rect 4813 17153 4847 17187
rect 5549 17153 5583 17187
rect 8861 17153 8895 17187
rect 9045 17153 9079 17187
rect 10425 17153 10459 17187
rect 10517 17153 10551 17187
rect 14197 17153 14231 17187
rect 14933 17153 14967 17187
rect 15853 17153 15887 17187
rect 18337 17153 18371 17187
rect 18889 17153 18923 17187
rect 19073 17153 19107 17187
rect 21465 17153 21499 17187
rect 26341 17153 26375 17187
rect 2421 17085 2455 17119
rect 3433 17085 3467 17119
rect 8585 17085 8619 17119
rect 5273 17017 5307 17051
rect 14657 17085 14691 17119
rect 20085 17085 20119 17119
rect 21373 17085 21407 17119
rect 25329 17085 25363 17119
rect 10333 17017 10367 17051
rect 21281 17017 21315 17051
rect 21925 17017 21959 17051
rect 26249 17017 26283 17051
rect 1777 16949 1811 16983
rect 2053 16949 2087 16983
rect 4905 16949 4939 16983
rect 5365 16949 5399 16983
rect 8033 16949 8067 16983
rect 8217 16949 8251 16983
rect 8677 16949 8711 16983
rect 9045 16949 9079 16983
rect 9321 16949 9355 16983
rect 9965 16949 9999 16983
rect 14749 16949 14783 16983
rect 15301 16949 15335 16983
rect 15761 16949 15795 16983
rect 18797 16949 18831 16983
rect 25697 16949 25731 16983
rect 26157 16949 26191 16983
rect 27169 16949 27203 16983
rect 2421 16745 2455 16779
rect 4905 16745 4939 16779
rect 8033 16745 8067 16779
rect 9045 16745 9079 16779
rect 9689 16745 9723 16779
rect 11253 16745 11287 16779
rect 11621 16745 11655 16779
rect 14381 16745 14415 16779
rect 15301 16745 15335 16779
rect 15761 16745 15795 16779
rect 18429 16745 18463 16779
rect 18889 16745 18923 16779
rect 21189 16745 21223 16779
rect 26525 16745 26559 16779
rect 1777 16677 1811 16711
rect 2789 16677 2823 16711
rect 5273 16677 5307 16711
rect 5702 16677 5736 16711
rect 9505 16677 9539 16711
rect 10149 16677 10183 16711
rect 15669 16677 15703 16711
rect 23756 16677 23790 16711
rect 2881 16609 2915 16643
rect 5457 16609 5491 16643
rect 8401 16609 8435 16643
rect 8493 16609 8527 16643
rect 10057 16609 10091 16643
rect 11713 16609 11747 16643
rect 21557 16609 21591 16643
rect 22201 16609 22235 16643
rect 2973 16541 3007 16575
rect 8585 16541 8619 16575
rect 10333 16541 10367 16575
rect 11897 16541 11931 16575
rect 15853 16541 15887 16575
rect 21649 16541 21683 16575
rect 21741 16541 21775 16575
rect 23489 16541 23523 16575
rect 2145 16473 2179 16507
rect 25789 16473 25823 16507
rect 6837 16405 6871 16439
rect 13369 16405 13403 16439
rect 24869 16405 24903 16439
rect 27077 16405 27111 16439
rect 1869 16201 1903 16235
rect 2697 16201 2731 16235
rect 4077 16201 4111 16235
rect 5549 16201 5583 16235
rect 8769 16201 8803 16235
rect 9505 16201 9539 16235
rect 10885 16201 10919 16235
rect 11345 16201 11379 16235
rect 15025 16201 15059 16235
rect 20637 16201 20671 16235
rect 21465 16201 21499 16235
rect 23489 16201 23523 16235
rect 2145 16133 2179 16167
rect 5825 16133 5859 16167
rect 8493 16133 8527 16167
rect 3249 16065 3283 16099
rect 10057 16065 10091 16099
rect 10517 16065 10551 16099
rect 11989 16065 12023 16099
rect 13737 16065 13771 16099
rect 13829 16065 13863 16099
rect 22017 16065 22051 16099
rect 23949 16065 23983 16099
rect 24685 16065 24719 16099
rect 25145 16065 25179 16099
rect 26249 16065 26283 16099
rect 13185 15997 13219 16031
rect 15761 15997 15795 16031
rect 16017 15997 16051 16031
rect 19257 15997 19291 16031
rect 24409 15997 24443 16031
rect 25973 15997 26007 16031
rect 2605 15929 2639 15963
rect 3065 15929 3099 15963
rect 12817 15929 12851 15963
rect 13645 15929 13679 15963
rect 19165 15929 19199 15963
rect 19502 15929 19536 15963
rect 21833 15929 21867 15963
rect 3157 15861 3191 15895
rect 3709 15861 3743 15895
rect 8125 15861 8159 15895
rect 9413 15861 9447 15895
rect 9873 15861 9907 15895
rect 9965 15861 9999 15895
rect 11713 15861 11747 15895
rect 13277 15861 13311 15895
rect 15393 15861 15427 15895
rect 17141 15861 17175 15895
rect 21281 15861 21315 15895
rect 21925 15861 21959 15895
rect 22477 15861 22511 15895
rect 22845 15861 22879 15895
rect 24041 15861 24075 15895
rect 24501 15861 24535 15895
rect 25421 15861 25455 15895
rect 25605 15861 25639 15895
rect 26065 15861 26099 15895
rect 26617 15861 26651 15895
rect 2421 15657 2455 15691
rect 9137 15657 9171 15691
rect 9505 15657 9539 15691
rect 11069 15657 11103 15691
rect 13369 15657 13403 15691
rect 15853 15657 15887 15691
rect 19349 15657 19383 15691
rect 21189 15657 21223 15691
rect 21557 15657 21591 15691
rect 21741 15657 21775 15691
rect 24133 15657 24167 15691
rect 24869 15657 24903 15691
rect 25329 15657 25363 15691
rect 26525 15657 26559 15691
rect 2789 15589 2823 15623
rect 5273 15589 5307 15623
rect 6460 15589 6494 15623
rect 17386 15589 17420 15623
rect 25237 15589 25271 15623
rect 26893 15589 26927 15623
rect 2329 15521 2363 15555
rect 2881 15521 2915 15555
rect 6193 15521 6227 15555
rect 9945 15521 9979 15555
rect 13737 15521 13771 15555
rect 22109 15521 22143 15555
rect 24501 15521 24535 15555
rect 26985 15521 27019 15555
rect 2973 15453 3007 15487
rect 9689 15453 9723 15487
rect 13829 15453 13863 15487
rect 14013 15453 14047 15487
rect 16313 15453 16347 15487
rect 17141 15453 17175 15487
rect 22201 15453 22235 15487
rect 22293 15453 22327 15487
rect 25421 15453 25455 15487
rect 27169 15453 27203 15487
rect 1685 15317 1719 15351
rect 3709 15317 3743 15351
rect 7573 15317 7607 15351
rect 15485 15317 15519 15351
rect 18521 15317 18555 15351
rect 23581 15317 23615 15351
rect 25973 15317 26007 15351
rect 2789 15113 2823 15147
rect 3065 15113 3099 15147
rect 3617 15113 3651 15147
rect 4629 15113 4663 15147
rect 6285 15113 6319 15147
rect 6377 15113 6411 15147
rect 1409 14977 1443 15011
rect 4169 14977 4203 15011
rect 5089 14977 5123 15011
rect 5641 14977 5675 15011
rect 5825 14977 5859 15011
rect 1676 14909 1710 14943
rect 9137 15113 9171 15147
rect 9781 15113 9815 15147
rect 12909 15113 12943 15147
rect 16773 15113 16807 15147
rect 17141 15113 17175 15147
rect 21189 15113 21223 15147
rect 21649 15113 21683 15147
rect 22753 15113 22787 15147
rect 24593 15113 24627 15147
rect 25329 15113 25363 15147
rect 25881 15113 25915 15147
rect 7389 14977 7423 15011
rect 13737 15045 13771 15079
rect 15209 15045 15243 15079
rect 17693 15045 17727 15079
rect 17785 15045 17819 15079
rect 24961 15045 24995 15079
rect 10333 14977 10367 15011
rect 11345 14977 11379 15011
rect 14289 14977 14323 15011
rect 7849 14909 7883 14943
rect 9137 14909 9171 14943
rect 13645 14909 13679 14943
rect 14105 14909 14139 14943
rect 18613 14977 18647 15011
rect 19073 14977 19107 15011
rect 22293 14977 22327 15011
rect 26433 14977 26467 15011
rect 18429 14909 18463 14943
rect 22017 14909 22051 14943
rect 3525 14841 3559 14875
rect 4077 14841 4111 14875
rect 6377 14841 6411 14875
rect 6653 14841 6687 14875
rect 7297 14841 7331 14875
rect 10609 14841 10643 14875
rect 11253 14841 11287 14875
rect 14749 14841 14783 14875
rect 17693 14841 17727 14875
rect 18521 14841 18555 14875
rect 21557 14841 21591 14875
rect 26341 14841 26375 14875
rect 3985 14773 4019 14807
rect 5181 14773 5215 14807
rect 5549 14773 5583 14807
rect 6837 14773 6871 14807
rect 7205 14773 7239 14807
rect 9321 14773 9355 14807
rect 10793 14773 10827 14807
rect 11161 14773 11195 14807
rect 13277 14773 13311 14807
rect 14197 14773 14231 14807
rect 17417 14773 17451 14807
rect 18061 14773 18095 14807
rect 20729 14773 20763 14807
rect 22109 14773 22143 14807
rect 23121 14773 23155 14807
rect 23397 14773 23431 14807
rect 25697 14773 25731 14807
rect 26249 14773 26283 14807
rect 26985 14773 27019 14807
rect 27261 14773 27295 14807
rect 2237 14569 2271 14603
rect 2421 14569 2455 14603
rect 5825 14569 5859 14603
rect 6929 14569 6963 14603
rect 9689 14569 9723 14603
rect 10885 14569 10919 14603
rect 13001 14569 13035 14603
rect 16681 14569 16715 14603
rect 16773 14569 16807 14603
rect 19349 14569 19383 14603
rect 21649 14569 21683 14603
rect 26801 14569 26835 14603
rect 2881 14501 2915 14535
rect 5917 14501 5951 14535
rect 13461 14501 13495 14535
rect 2789 14433 2823 14467
rect 4353 14433 4387 14467
rect 6469 14433 6503 14467
rect 9505 14433 9539 14467
rect 10057 14433 10091 14467
rect 13369 14433 13403 14467
rect 18245 14433 18279 14467
rect 18705 14433 18739 14467
rect 22017 14433 22051 14467
rect 2973 14365 3007 14399
rect 3709 14365 3743 14399
rect 6009 14365 6043 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 13645 14365 13679 14399
rect 16865 14365 16899 14399
rect 18797 14365 18831 14399
rect 18889 14365 18923 14399
rect 22109 14365 22143 14399
rect 22293 14365 22327 14399
rect 5273 14297 5307 14331
rect 18061 14297 18095 14331
rect 1685 14229 1719 14263
rect 4905 14229 4939 14263
rect 5457 14229 5491 14263
rect 8953 14229 8987 14263
rect 9321 14229 9355 14263
rect 12541 14229 12575 14263
rect 14105 14229 14139 14263
rect 15577 14229 15611 14263
rect 16313 14229 16347 14263
rect 18337 14229 18371 14263
rect 24317 14229 24351 14263
rect 25973 14229 26007 14263
rect 1593 14025 1627 14059
rect 2513 14025 2547 14059
rect 4721 14025 4755 14059
rect 6561 14025 6595 14059
rect 8861 14025 8895 14059
rect 10333 14025 10367 14059
rect 10609 14025 10643 14059
rect 14105 14025 14139 14059
rect 16313 14025 16347 14059
rect 17141 14025 17175 14059
rect 19073 14025 19107 14059
rect 20545 14025 20579 14059
rect 21281 14025 21315 14059
rect 24225 14025 24259 14059
rect 3617 13957 3651 13991
rect 5089 13957 5123 13991
rect 12173 13957 12207 13991
rect 13829 13957 13863 13991
rect 15117 13957 15151 13991
rect 15301 13957 15335 13991
rect 18337 13957 18371 13991
rect 26709 13957 26743 13991
rect 2421 13889 2455 13923
rect 3157 13889 3191 13923
rect 3893 13889 3927 13923
rect 4353 13889 4387 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 12449 13889 12483 13923
rect 14841 13889 14875 13923
rect 15761 13889 15795 13923
rect 15853 13889 15887 13923
rect 17509 13889 17543 13923
rect 21833 13889 21867 13923
rect 1409 13821 1443 13855
rect 2053 13821 2087 13855
rect 8953 13821 8987 13855
rect 12705 13821 12739 13855
rect 15669 13821 15703 13855
rect 17877 13821 17911 13855
rect 19165 13821 19199 13855
rect 21557 13821 21591 13855
rect 22293 13821 22327 13855
rect 24317 13821 24351 13855
rect 24573 13821 24607 13855
rect 26525 13821 26559 13855
rect 27077 13821 27111 13855
rect 2881 13753 2915 13787
rect 5549 13753 5583 13787
rect 9198 13753 9232 13787
rect 11805 13753 11839 13787
rect 16681 13753 16715 13787
rect 19410 13753 19444 13787
rect 2973 13685 3007 13719
rect 5181 13685 5215 13719
rect 6193 13685 6227 13719
rect 21373 13685 21407 13719
rect 21649 13685 21683 13719
rect 21741 13685 21775 13719
rect 25697 13685 25731 13719
rect 2973 13481 3007 13515
rect 5733 13481 5767 13515
rect 8217 13481 8251 13515
rect 9413 13481 9447 13515
rect 13645 13481 13679 13515
rect 17233 13481 17267 13515
rect 18429 13481 18463 13515
rect 21373 13481 21407 13515
rect 23121 13481 23155 13515
rect 25237 13481 25271 13515
rect 12256 13413 12290 13447
rect 1593 13345 1627 13379
rect 1860 13345 1894 13379
rect 5641 13345 5675 13379
rect 7021 13345 7055 13379
rect 8401 13345 8435 13379
rect 11989 13345 12023 13379
rect 15117 13345 15151 13379
rect 15669 13345 15703 13379
rect 15761 13345 15795 13379
rect 19165 13345 19199 13379
rect 21741 13345 21775 13379
rect 21997 13345 22031 13379
rect 5089 13277 5123 13311
rect 5917 13277 5951 13311
rect 15853 13277 15887 13311
rect 17325 13277 17359 13311
rect 17417 13277 17451 13311
rect 19257 13277 19291 13311
rect 19441 13277 19475 13311
rect 25329 13277 25363 13311
rect 25513 13277 25547 13311
rect 6837 13209 6871 13243
rect 16865 13209 16899 13243
rect 18797 13209 18831 13243
rect 3249 13141 3283 13175
rect 5273 13141 5307 13175
rect 9045 13141 9079 13175
rect 9965 13141 9999 13175
rect 13369 13141 13403 13175
rect 15301 13141 15335 13175
rect 24317 13141 24351 13175
rect 24869 13141 24903 13175
rect 25881 13141 25915 13175
rect 2053 12937 2087 12971
rect 2329 12937 2363 12971
rect 4813 12937 4847 12971
rect 4997 12937 5031 12971
rect 6009 12937 6043 12971
rect 6377 12937 6411 12971
rect 7113 12937 7147 12971
rect 9781 12937 9815 12971
rect 12081 12937 12115 12971
rect 13737 12937 13771 12971
rect 15485 12937 15519 12971
rect 16589 12937 16623 12971
rect 17325 12937 17359 12971
rect 18797 12937 18831 12971
rect 21833 12937 21867 12971
rect 25329 12937 25363 12971
rect 4537 12869 4571 12903
rect 12633 12869 12667 12903
rect 15393 12869 15427 12903
rect 17601 12869 17635 12903
rect 19809 12869 19843 12903
rect 22109 12869 22143 12903
rect 25605 12869 25639 12903
rect 4169 12801 4203 12835
rect 5457 12801 5491 12835
rect 5549 12801 5583 12835
rect 8125 12801 8159 12835
rect 14473 12801 14507 12835
rect 15945 12801 15979 12835
rect 16129 12801 16163 12835
rect 16957 12801 16991 12835
rect 19441 12801 19475 12835
rect 20177 12801 20211 12835
rect 24041 12801 24075 12835
rect 24777 12801 24811 12835
rect 1409 12733 1443 12767
rect 5365 12733 5399 12767
rect 13461 12733 13495 12767
rect 14289 12733 14323 12767
rect 14381 12733 14415 12767
rect 24593 12733 24627 12767
rect 24685 12733 24719 12767
rect 25789 12733 25823 12767
rect 2697 12665 2731 12699
rect 8033 12665 8067 12699
rect 8370 12665 8404 12699
rect 15025 12665 15059 12699
rect 15853 12665 15887 12699
rect 18705 12665 18739 12699
rect 19257 12665 19291 12699
rect 26034 12665 26068 12699
rect 1593 12597 1627 12631
rect 7665 12597 7699 12631
rect 9505 12597 9539 12631
rect 13921 12597 13955 12631
rect 18337 12597 18371 12631
rect 19165 12597 19199 12631
rect 24225 12597 24259 12631
rect 27169 12597 27203 12631
rect 6377 12393 6411 12427
rect 12817 12393 12851 12427
rect 14013 12393 14047 12427
rect 15577 12393 15611 12427
rect 16037 12393 16071 12427
rect 17601 12393 17635 12427
rect 19073 12393 19107 12427
rect 19533 12393 19567 12427
rect 24869 12393 24903 12427
rect 25513 12393 25547 12427
rect 26249 12393 26283 12427
rect 15117 12325 15151 12359
rect 1409 12257 1443 12291
rect 1676 12257 1710 12291
rect 4997 12257 5031 12291
rect 5264 12257 5298 12291
rect 8401 12257 8435 12291
rect 10057 12257 10091 12291
rect 17509 12257 17543 12291
rect 19257 12257 19291 12291
rect 21649 12257 21683 12291
rect 21916 12257 21950 12291
rect 24225 12257 24259 12291
rect 24777 12257 24811 12291
rect 8493 12189 8527 12223
rect 8677 12189 8711 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 17693 12189 17727 12223
rect 24961 12189 24995 12223
rect 26525 12189 26559 12223
rect 9505 12121 9539 12155
rect 23949 12121 23983 12155
rect 24409 12121 24443 12155
rect 2789 12053 2823 12087
rect 7941 12053 7975 12087
rect 8033 12053 8067 12087
rect 9689 12053 9723 12087
rect 16497 12053 16531 12087
rect 17141 12053 17175 12087
rect 18889 12053 18923 12087
rect 23029 12053 23063 12087
rect 25881 12053 25915 12087
rect 2789 11849 2823 11883
rect 5457 11849 5491 11883
rect 7297 11849 7331 11883
rect 7757 11849 7791 11883
rect 8953 11849 8987 11883
rect 17509 11849 17543 11883
rect 17785 11849 17819 11883
rect 21741 11849 21775 11883
rect 24869 11849 24903 11883
rect 25237 11849 25271 11883
rect 4813 11781 4847 11815
rect 9413 11781 9447 11815
rect 22017 11781 22051 11815
rect 23489 11781 23523 11815
rect 3433 11713 3467 11747
rect 5181 11713 5215 11747
rect 8401 11713 8435 11747
rect 9965 11713 9999 11747
rect 10793 11713 10827 11747
rect 12817 11713 12851 11747
rect 15945 11713 15979 11747
rect 17049 11713 17083 11747
rect 18061 11713 18095 11747
rect 18613 11713 18647 11747
rect 19441 11713 19475 11747
rect 24317 11713 24351 11747
rect 24501 11713 24535 11747
rect 26249 11713 26283 11747
rect 26341 11713 26375 11747
rect 1409 11645 1443 11679
rect 1961 11645 1995 11679
rect 8217 11645 8251 11679
rect 8309 11645 8343 11679
rect 16865 11645 16899 11679
rect 24225 11645 24259 11679
rect 3678 11577 3712 11611
rect 9321 11577 9355 11611
rect 9873 11577 9907 11611
rect 12725 11577 12759 11611
rect 13084 11577 13118 11611
rect 16313 11577 16347 11611
rect 19349 11577 19383 11611
rect 19708 11577 19742 11611
rect 26157 11577 26191 11611
rect 1593 11509 1627 11543
rect 2513 11509 2547 11543
rect 3341 11509 3375 11543
rect 7849 11509 7883 11543
rect 9781 11509 9815 11543
rect 10517 11509 10551 11543
rect 10977 11509 11011 11543
rect 14197 11509 14231 11543
rect 16405 11509 16439 11543
rect 16773 11509 16807 11543
rect 18889 11509 18923 11543
rect 20821 11509 20855 11543
rect 23857 11509 23891 11543
rect 25605 11509 25639 11543
rect 25789 11509 25823 11543
rect 1685 11305 1719 11339
rect 2789 11305 2823 11339
rect 2881 11305 2915 11339
rect 4721 11305 4755 11339
rect 7941 11305 7975 11339
rect 8309 11305 8343 11339
rect 9505 11305 9539 11339
rect 10517 11305 10551 11339
rect 19993 11305 20027 11339
rect 23305 11305 23339 11339
rect 23949 11305 23983 11339
rect 24409 11305 24443 11339
rect 25329 11305 25363 11339
rect 26525 11305 26559 11339
rect 26985 11305 27019 11339
rect 2329 11237 2363 11271
rect 3433 11237 3467 11271
rect 8769 11237 8803 11271
rect 16282 11237 16316 11271
rect 18880 11237 18914 11271
rect 22192 11237 22226 11271
rect 25237 11237 25271 11271
rect 26893 11237 26927 11271
rect 4629 11169 4663 11203
rect 5089 11169 5123 11203
rect 13073 11169 13107 11203
rect 18613 11169 18647 11203
rect 21925 11169 21959 11203
rect 25881 11169 25915 11203
rect 2973 11101 3007 11135
rect 5181 11101 5215 11135
rect 5273 11101 5307 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 12817 11101 12851 11135
rect 16037 11101 16071 11135
rect 25421 11101 25455 11135
rect 27077 11101 27111 11135
rect 2421 11033 2455 11067
rect 9965 11033 9999 11067
rect 14197 11033 14231 11067
rect 17785 11033 17819 11067
rect 24869 11033 24903 11067
rect 5733 10965 5767 10999
rect 10149 10965 10183 10999
rect 17417 10965 17451 10999
rect 1869 10761 1903 10795
rect 2421 10761 2455 10795
rect 4169 10761 4203 10795
rect 4997 10761 5031 10795
rect 5181 10761 5215 10795
rect 11437 10761 11471 10795
rect 12265 10761 12299 10795
rect 12909 10761 12943 10795
rect 16037 10761 16071 10795
rect 18981 10761 19015 10795
rect 22017 10761 22051 10795
rect 22293 10761 22327 10795
rect 23489 10761 23523 10795
rect 24961 10761 24995 10795
rect 25329 10761 25363 10795
rect 25881 10761 25915 10795
rect 26341 10761 26375 10795
rect 27353 10761 27387 10795
rect 2329 10693 2363 10727
rect 14933 10693 14967 10727
rect 18705 10693 18739 10727
rect 26617 10693 26651 10727
rect 3065 10625 3099 10659
rect 5733 10625 5767 10659
rect 9229 10625 9263 10659
rect 10701 10625 10735 10659
rect 11253 10625 11287 10659
rect 15761 10625 15795 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 24133 10625 24167 10659
rect 24225 10625 24259 10659
rect 3985 10557 4019 10591
rect 4629 10557 4663 10591
rect 5641 10557 5675 10591
rect 6193 10557 6227 10591
rect 9965 10557 9999 10591
rect 16773 10557 16807 10591
rect 23121 10557 23155 10591
rect 24041 10557 24075 10591
rect 26433 10557 26467 10591
rect 26985 10557 27019 10591
rect 2881 10489 2915 10523
rect 3433 10489 3467 10523
rect 3893 10489 3927 10523
rect 10517 10489 10551 10523
rect 11253 10489 11287 10523
rect 13645 10489 13679 10523
rect 2789 10421 2823 10455
rect 5549 10421 5583 10455
rect 9505 10421 9539 10455
rect 10057 10421 10091 10455
rect 10425 10421 10459 10455
rect 11161 10421 11195 10455
rect 13461 10421 13495 10455
rect 16405 10421 16439 10455
rect 17417 10421 17451 10455
rect 23673 10421 23707 10455
rect 2329 10217 2363 10251
rect 4997 10217 5031 10251
rect 5365 10217 5399 10251
rect 6929 10217 6963 10251
rect 10425 10217 10459 10251
rect 12633 10217 12667 10251
rect 13093 10217 13127 10251
rect 15301 10217 15335 10251
rect 15761 10217 15795 10251
rect 16865 10217 16899 10251
rect 19349 10217 19383 10251
rect 23029 10217 23063 10251
rect 23765 10217 23799 10251
rect 25513 10217 25547 10251
rect 26709 10217 26743 10251
rect 4813 10149 4847 10183
rect 10333 10149 10367 10183
rect 13921 10149 13955 10183
rect 16497 10149 16531 10183
rect 24777 10149 24811 10183
rect 2789 10081 2823 10115
rect 11069 10081 11103 10115
rect 15669 10081 15703 10115
rect 18613 10081 18647 10115
rect 21916 10081 21950 10115
rect 26525 10081 26559 10115
rect 2881 10013 2915 10047
rect 2973 10013 3007 10047
rect 5457 10013 5491 10047
rect 5641 10013 5675 10047
rect 7021 10013 7055 10047
rect 7113 10013 7147 10047
rect 10609 10013 10643 10047
rect 13185 10013 13219 10047
rect 13369 10013 13403 10047
rect 14013 10013 14047 10047
rect 14105 10013 14139 10047
rect 15853 10013 15887 10047
rect 18705 10013 18739 10047
rect 18889 10013 18923 10047
rect 21649 10013 21683 10047
rect 24869 10013 24903 10047
rect 25053 10013 25087 10047
rect 2421 9945 2455 9979
rect 9965 9945 9999 9979
rect 13553 9945 13587 9979
rect 14657 9945 14691 9979
rect 1685 9877 1719 9911
rect 3433 9877 3467 9911
rect 6561 9877 6595 9911
rect 9321 9877 9355 9911
rect 12265 9877 12299 9911
rect 12725 9877 12759 9911
rect 18245 9877 18279 9911
rect 24409 9877 24443 9911
rect 2789 9673 2823 9707
rect 5825 9673 5859 9707
rect 10977 9673 11011 9707
rect 11897 9673 11931 9707
rect 21741 9673 21775 9707
rect 22017 9673 22051 9707
rect 27353 9673 27387 9707
rect 2513 9605 2547 9639
rect 6285 9605 6319 9639
rect 15393 9605 15427 9639
rect 17877 9605 17911 9639
rect 18337 9605 18371 9639
rect 20085 9605 20119 9639
rect 25329 9605 25363 9639
rect 26617 9605 26651 9639
rect 2145 9537 2179 9571
rect 3249 9537 3283 9571
rect 3433 9537 3467 9571
rect 13001 9537 13035 9571
rect 14565 9537 14599 9571
rect 16037 9537 16071 9571
rect 19625 9537 19659 9571
rect 25697 9537 25731 9571
rect 1409 9469 1443 9503
rect 4261 9469 4295 9503
rect 6837 9469 6871 9503
rect 9229 9469 9263 9503
rect 9321 9469 9355 9503
rect 9588 9469 9622 9503
rect 12265 9469 12299 9503
rect 12909 9469 12943 9503
rect 14381 9469 14415 9503
rect 18981 9469 19015 9503
rect 19441 9469 19475 9503
rect 23489 9469 23523 9503
rect 23673 9469 23707 9503
rect 26433 9469 26467 9503
rect 26985 9469 27019 9503
rect 3157 9401 3191 9435
rect 3893 9401 3927 9435
rect 4353 9401 4387 9435
rect 5457 9401 5491 9435
rect 7082 9401 7116 9435
rect 8953 9401 8987 9435
rect 18705 9401 18739 9435
rect 23940 9401 23974 9435
rect 1593 9333 1627 9367
rect 5089 9333 5123 9367
rect 6561 9333 6595 9367
rect 8217 9333 8251 9367
rect 9045 9333 9079 9367
rect 10701 9333 10735 9367
rect 12449 9333 12483 9367
rect 12817 9333 12851 9367
rect 13553 9333 13587 9367
rect 14013 9333 14047 9367
rect 14473 9333 14507 9367
rect 15669 9333 15703 9367
rect 18797 9333 18831 9367
rect 19073 9333 19107 9367
rect 19533 9333 19567 9367
rect 25053 9333 25087 9367
rect 2697 9129 2731 9163
rect 9137 9129 9171 9163
rect 10333 9129 10367 9163
rect 11713 9129 11747 9163
rect 12449 9129 12483 9163
rect 13369 9129 13403 9163
rect 14749 9129 14783 9163
rect 15761 9129 15795 9163
rect 16313 9129 16347 9163
rect 18613 9129 18647 9163
rect 18889 9129 18923 9163
rect 24869 9129 24903 9163
rect 25237 9129 25271 9163
rect 25329 9129 25363 9163
rect 26709 9129 26743 9163
rect 12725 9061 12759 9095
rect 17417 9061 17451 9095
rect 17877 9061 17911 9095
rect 24501 9061 24535 9095
rect 1409 8993 1443 9027
rect 2513 8993 2547 9027
rect 10057 8993 10091 9027
rect 13277 8993 13311 9027
rect 19441 8993 19475 9027
rect 21925 8993 21959 9027
rect 26525 8993 26559 9027
rect 4077 8925 4111 8959
rect 7297 8925 7331 8959
rect 11805 8925 11839 8959
rect 11897 8925 11931 8959
rect 13461 8925 13495 8959
rect 16405 8925 16439 8959
rect 16497 8925 16531 8959
rect 17969 8925 18003 8959
rect 18061 8925 18095 8959
rect 19533 8925 19567 8959
rect 19717 8925 19751 8959
rect 22017 8925 22051 8959
rect 22109 8925 22143 8959
rect 23857 8925 23891 8959
rect 25513 8925 25547 8959
rect 12909 8857 12943 8891
rect 19073 8857 19107 8891
rect 1593 8789 1627 8823
rect 3065 8789 3099 8823
rect 3709 8789 3743 8823
rect 6653 8789 6687 8823
rect 7021 8789 7055 8823
rect 11345 8789 11379 8823
rect 14105 8789 14139 8823
rect 14473 8789 14507 8823
rect 15945 8789 15979 8823
rect 17509 8789 17543 8823
rect 21557 8789 21591 8823
rect 23765 8789 23799 8823
rect 25881 8789 25915 8823
rect 2053 8585 2087 8619
rect 8217 8585 8251 8619
rect 12265 8585 12299 8619
rect 13645 8585 13679 8619
rect 15209 8585 15243 8619
rect 17601 8585 17635 8619
rect 18429 8585 18463 8619
rect 18981 8585 19015 8619
rect 19993 8585 20027 8619
rect 20545 8585 20579 8619
rect 21649 8585 21683 8619
rect 21925 8585 21959 8619
rect 23397 8585 23431 8619
rect 24501 8585 24535 8619
rect 24961 8585 24995 8619
rect 25421 8585 25455 8619
rect 26525 8585 26559 8619
rect 27169 8585 27203 8619
rect 1593 8517 1627 8551
rect 9873 8517 9907 8551
rect 13001 8517 13035 8551
rect 17049 8517 17083 8551
rect 27537 8517 27571 8551
rect 4261 8449 4295 8483
rect 19441 8449 19475 8483
rect 19533 8449 19567 8483
rect 22477 8449 22511 8483
rect 25329 8449 25363 8483
rect 26065 8449 26099 8483
rect 1409 8381 1443 8415
rect 3985 8381 4019 8415
rect 6837 8381 6871 8415
rect 10057 8381 10091 8415
rect 10149 8381 10183 8415
rect 15669 8381 15703 8415
rect 18889 8381 18923 8415
rect 19349 8381 19383 8415
rect 20729 8381 20763 8415
rect 21281 8381 21315 8415
rect 22385 8381 22419 8415
rect 25789 8381 25823 8415
rect 26985 8381 27019 8415
rect 2605 8313 2639 8347
rect 3525 8313 3559 8347
rect 6561 8313 6595 8347
rect 7082 8313 7116 8347
rect 9781 8313 9815 8347
rect 10416 8313 10450 8347
rect 14841 8313 14875 8347
rect 15485 8313 15519 8347
rect 15936 8313 15970 8347
rect 20361 8313 20395 8347
rect 3617 8245 3651 8279
rect 4077 8245 4111 8279
rect 6285 8245 6319 8279
rect 11529 8245 11563 8279
rect 11897 8245 11931 8279
rect 22293 8245 22327 8279
rect 22937 8245 22971 8279
rect 25881 8245 25915 8279
rect 1685 8041 1719 8075
rect 2329 8041 2363 8075
rect 2789 8041 2823 8075
rect 3709 8041 3743 8075
rect 4445 8041 4479 8075
rect 11437 8041 11471 8075
rect 11713 8041 11747 8075
rect 12541 8041 12575 8075
rect 12909 8041 12943 8075
rect 16129 8041 16163 8075
rect 17233 8041 17267 8075
rect 17693 8041 17727 8075
rect 18337 8041 18371 8075
rect 19073 8041 19107 8075
rect 19441 8041 19475 8075
rect 19717 8041 19751 8075
rect 21649 8041 21683 8075
rect 22385 8041 22419 8075
rect 23765 8041 23799 8075
rect 25881 8041 25915 8075
rect 26709 8041 26743 8075
rect 4537 7973 4571 8007
rect 10333 7973 10367 8007
rect 17601 7973 17635 8007
rect 21925 7973 21959 8007
rect 24961 7973 24995 8007
rect 7113 7905 7147 7939
rect 9873 7905 9907 7939
rect 17141 7905 17175 7939
rect 22753 7905 22787 7939
rect 25329 7905 25363 7939
rect 26525 7905 26559 7939
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 4721 7837 4755 7871
rect 17785 7837 17819 7871
rect 22845 7837 22879 7871
rect 23029 7837 23063 7871
rect 4077 7769 4111 7803
rect 2421 7701 2455 7735
rect 6929 7701 6963 7735
rect 7389 7701 7423 7735
rect 15761 7701 15795 7735
rect 16957 7701 16991 7735
rect 24133 7701 24167 7735
rect 25513 7701 25547 7735
rect 4261 7497 4295 7531
rect 6285 7497 6319 7531
rect 8217 7497 8251 7531
rect 16957 7497 16991 7531
rect 18521 7497 18555 7531
rect 22017 7497 22051 7531
rect 25053 7497 25087 7531
rect 26893 7497 26927 7531
rect 27629 7497 27663 7531
rect 17233 7429 17267 7463
rect 23673 7429 23707 7463
rect 26617 7429 26651 7463
rect 4629 7361 4663 7395
rect 6837 7361 6871 7395
rect 12449 7361 12483 7395
rect 16221 7361 16255 7395
rect 19165 7361 19199 7395
rect 19349 7361 19383 7395
rect 19717 7361 19751 7395
rect 21925 7361 21959 7395
rect 22661 7361 22695 7395
rect 24225 7361 24259 7395
rect 1409 7293 1443 7327
rect 2513 7293 2547 7327
rect 9045 7293 9079 7327
rect 15577 7293 15611 7327
rect 16037 7293 16071 7327
rect 24041 7293 24075 7327
rect 25237 7293 25271 7327
rect 27445 7293 27479 7327
rect 27997 7293 28031 7327
rect 2053 7225 2087 7259
rect 2421 7225 2455 7259
rect 2780 7225 2814 7259
rect 6653 7225 6687 7259
rect 7082 7225 7116 7259
rect 8953 7225 8987 7259
rect 9312 7225 9346 7259
rect 12265 7225 12299 7259
rect 12694 7225 12728 7259
rect 16129 7225 16163 7259
rect 17877 7225 17911 7259
rect 19073 7225 19107 7259
rect 21557 7225 21591 7259
rect 22385 7225 22419 7259
rect 23489 7225 23523 7259
rect 25482 7225 25516 7259
rect 1593 7157 1627 7191
rect 3893 7157 3927 7191
rect 4905 7157 4939 7191
rect 10425 7157 10459 7191
rect 13829 7157 13863 7191
rect 15209 7157 15243 7191
rect 15669 7157 15703 7191
rect 18705 7157 18739 7191
rect 22477 7157 22511 7191
rect 23121 7157 23155 7191
rect 24133 7157 24167 7191
rect 24685 7157 24719 7191
rect 9137 6953 9171 6987
rect 10057 6953 10091 6987
rect 11253 6953 11287 6987
rect 17601 6953 17635 6987
rect 17785 6953 17819 6987
rect 19165 6953 19199 6987
rect 19901 6953 19935 6987
rect 22109 6953 22143 6987
rect 23029 6953 23063 6987
rect 23397 6953 23431 6987
rect 17325 6885 17359 6919
rect 22385 6885 22419 6919
rect 22845 6885 22879 6919
rect 1409 6817 1443 6851
rect 2513 6817 2547 6851
rect 6837 6817 6871 6851
rect 11621 6817 11655 6851
rect 11713 6817 11747 6851
rect 13737 6817 13771 6851
rect 15557 6817 15591 6851
rect 19257 6817 19291 6851
rect 23489 6817 23523 6851
rect 24133 6817 24167 6851
rect 26525 6817 26559 6851
rect 2421 6749 2455 6783
rect 6929 6749 6963 6783
rect 7021 6749 7055 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 11897 6749 11931 6783
rect 13829 6749 13863 6783
rect 13921 6749 13955 6783
rect 15301 6749 15335 6783
rect 19441 6749 19475 6783
rect 23581 6749 23615 6783
rect 2697 6681 2731 6715
rect 9689 6681 9723 6715
rect 12633 6681 12667 6715
rect 13369 6681 13403 6715
rect 26709 6681 26743 6715
rect 1593 6613 1627 6647
rect 1961 6613 1995 6647
rect 3157 6613 3191 6647
rect 6469 6613 6503 6647
rect 7481 6613 7515 6647
rect 13001 6613 13035 6647
rect 16681 6613 16715 6647
rect 18797 6613 18831 6647
rect 25237 6613 25271 6647
rect 2053 6409 2087 6443
rect 2421 6409 2455 6443
rect 5825 6409 5859 6443
rect 7021 6409 7055 6443
rect 8861 6409 8895 6443
rect 10057 6409 10091 6443
rect 11345 6409 11379 6443
rect 11989 6409 12023 6443
rect 14289 6409 14323 6443
rect 14841 6409 14875 6443
rect 19165 6409 19199 6443
rect 19441 6409 19475 6443
rect 22753 6409 22787 6443
rect 23673 6409 23707 6443
rect 27353 6409 27387 6443
rect 6561 6341 6595 6375
rect 17877 6341 17911 6375
rect 22385 6341 22419 6375
rect 24685 6341 24719 6375
rect 26617 6341 26651 6375
rect 7573 6273 7607 6307
rect 9597 6273 9631 6307
rect 10701 6273 10735 6307
rect 13369 6273 13403 6307
rect 13461 6273 13495 6307
rect 13921 6273 13955 6307
rect 16313 6273 16347 6307
rect 16773 6273 16807 6307
rect 18521 6273 18555 6307
rect 18613 6273 18647 6307
rect 19625 6273 19659 6307
rect 23121 6273 23155 6307
rect 24225 6273 24259 6307
rect 1409 6205 1443 6239
rect 2513 6205 2547 6239
rect 3157 6205 3191 6239
rect 3985 6205 4019 6239
rect 7389 6205 7423 6239
rect 9137 6205 9171 6239
rect 9873 6205 9907 6239
rect 10425 6205 10459 6239
rect 15577 6205 15611 6239
rect 16221 6205 16255 6239
rect 17509 6205 17543 6239
rect 18429 6205 18463 6239
rect 23489 6205 23523 6239
rect 24133 6205 24167 6239
rect 26433 6205 26467 6239
rect 26985 6205 27019 6239
rect 3433 6137 3467 6171
rect 3893 6137 3927 6171
rect 4252 6137 4286 6171
rect 6193 6137 6227 6171
rect 7481 6137 7515 6171
rect 10517 6137 10551 6171
rect 12817 6137 12851 6171
rect 15301 6137 15335 6171
rect 16129 6137 16163 6171
rect 19870 6137 19904 6171
rect 24041 6137 24075 6171
rect 1593 6069 1627 6103
rect 2697 6069 2731 6103
rect 5365 6069 5399 6103
rect 11621 6069 11655 6103
rect 12909 6069 12943 6103
rect 13277 6069 13311 6103
rect 15761 6069 15795 6103
rect 18061 6069 18095 6103
rect 21005 6069 21039 6103
rect 1593 5865 1627 5899
rect 2329 5865 2363 5899
rect 2789 5865 2823 5899
rect 2881 5865 2915 5899
rect 4077 5865 4111 5899
rect 6561 5865 6595 5899
rect 7021 5865 7055 5899
rect 7757 5865 7791 5899
rect 8125 5865 8159 5899
rect 9505 5865 9539 5899
rect 10241 5865 10275 5899
rect 12265 5865 12299 5899
rect 12909 5865 12943 5899
rect 15761 5865 15795 5899
rect 18153 5865 18187 5899
rect 19441 5865 19475 5899
rect 19809 5865 19843 5899
rect 24133 5865 24167 5899
rect 18797 5797 18831 5831
rect 22998 5797 23032 5831
rect 4445 5729 4479 5763
rect 12817 5729 12851 5763
rect 15669 5729 15703 5763
rect 26525 5729 26559 5763
rect 3065 5661 3099 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 8217 5661 8251 5695
rect 8401 5661 8435 5695
rect 10057 5661 10091 5695
rect 13093 5661 13127 5695
rect 15853 5661 15887 5695
rect 18889 5661 18923 5695
rect 19073 5661 19107 5695
rect 22753 5661 22787 5695
rect 7665 5593 7699 5627
rect 26709 5593 26743 5627
rect 2421 5525 2455 5559
rect 12449 5525 12483 5559
rect 13461 5525 13495 5559
rect 15025 5525 15059 5559
rect 15301 5525 15335 5559
rect 18429 5525 18463 5559
rect 2421 5321 2455 5355
rect 3985 5321 4019 5355
rect 4997 5321 5031 5355
rect 5733 5321 5767 5355
rect 7573 5321 7607 5355
rect 8585 5321 8619 5355
rect 9045 5321 9079 5355
rect 12173 5321 12207 5355
rect 15025 5321 15059 5355
rect 15393 5321 15427 5355
rect 15669 5321 15703 5355
rect 17877 5321 17911 5355
rect 18889 5321 18923 5355
rect 22753 5321 22787 5355
rect 23029 5321 23063 5355
rect 23397 5321 23431 5355
rect 27353 5321 27387 5355
rect 13829 5253 13863 5287
rect 18521 5253 18555 5287
rect 3525 5185 3559 5219
rect 4629 5185 4663 5219
rect 8217 5185 8251 5219
rect 12449 5185 12483 5219
rect 15945 5185 15979 5219
rect 19441 5185 19475 5219
rect 19901 5185 19935 5219
rect 21189 5185 21223 5219
rect 1409 5117 1443 5151
rect 3893 5117 3927 5151
rect 4353 5117 4387 5151
rect 19349 5117 19383 5151
rect 20269 5117 20303 5151
rect 21373 5117 21407 5151
rect 26433 5117 26467 5151
rect 26985 5117 27019 5151
rect 2053 5049 2087 5083
rect 3157 5049 3191 5083
rect 4445 5049 4479 5083
rect 5365 5049 5399 5083
rect 8033 5049 8067 5083
rect 9321 5049 9355 5083
rect 11897 5049 11931 5083
rect 12694 5049 12728 5083
rect 14105 5049 14139 5083
rect 19257 5049 19291 5083
rect 20729 5049 20763 5083
rect 21618 5049 21652 5083
rect 1593 4981 1627 5015
rect 7021 4981 7055 5015
rect 7481 4981 7515 5015
rect 7941 4981 7975 5015
rect 26617 4981 26651 5015
rect 2513 4777 2547 4811
rect 4077 4777 4111 4811
rect 11069 4777 11103 4811
rect 12541 4777 12575 4811
rect 12633 4777 12667 4811
rect 13093 4777 13127 4811
rect 15669 4777 15703 4811
rect 18521 4777 18555 4811
rect 19257 4777 19291 4811
rect 19625 4777 19659 4811
rect 21373 4777 21407 4811
rect 2053 4709 2087 4743
rect 13001 4709 13035 4743
rect 19165 4709 19199 4743
rect 1409 4641 1443 4675
rect 2789 4641 2823 4675
rect 4445 4641 4479 4675
rect 7104 4641 7138 4675
rect 9689 4641 9723 4675
rect 9945 4641 9979 4675
rect 15761 4641 15795 4675
rect 26525 4641 26559 4675
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 6837 4573 6871 4607
rect 13277 4573 13311 4607
rect 15945 4573 15979 4607
rect 19717 4573 19751 4607
rect 19809 4573 19843 4607
rect 3341 4505 3375 4539
rect 1593 4437 1627 4471
rect 2973 4437 3007 4471
rect 3893 4437 3927 4471
rect 8217 4437 8251 4471
rect 15301 4437 15335 4471
rect 26709 4437 26743 4471
rect 2881 4233 2915 4267
rect 4169 4233 4203 4267
rect 4629 4233 4663 4267
rect 7113 4233 7147 4267
rect 8033 4233 8067 4267
rect 9781 4233 9815 4267
rect 10149 4233 10183 4267
rect 12725 4233 12759 4267
rect 13001 4233 13035 4267
rect 14381 4233 14415 4267
rect 16221 4233 16255 4267
rect 19073 4233 19107 4267
rect 20085 4233 20119 4267
rect 27353 4233 27387 4267
rect 7573 4165 7607 4199
rect 15945 4165 15979 4199
rect 5181 4097 5215 4131
rect 5641 4097 5675 4131
rect 8677 4097 8711 4131
rect 13369 4097 13403 4131
rect 18613 4097 18647 4131
rect 19625 4097 19659 4131
rect 20453 4097 20487 4131
rect 1501 4029 1535 4063
rect 3249 4029 3283 4063
rect 4997 4029 5031 4063
rect 7941 4029 7975 4063
rect 8493 4029 8527 4063
rect 14565 4029 14599 4063
rect 14821 4029 14855 4063
rect 26433 4029 26467 4063
rect 26985 4029 27019 4063
rect 27537 4029 27571 4063
rect 28089 4029 28123 4063
rect 1768 3961 1802 3995
rect 3709 3961 3743 3995
rect 8401 3961 8435 3995
rect 19533 3961 19567 3995
rect 20821 3961 20855 3995
rect 4537 3893 4571 3927
rect 5089 3893 5123 3927
rect 6561 3893 6595 3927
rect 18889 3893 18923 3927
rect 19441 3893 19475 3927
rect 26617 3893 26651 3927
rect 27721 3893 27755 3927
rect 2329 3689 2363 3723
rect 3157 3689 3191 3723
rect 3893 3689 3927 3723
rect 4077 3689 4111 3723
rect 8125 3689 8159 3723
rect 15853 3689 15887 3723
rect 19901 3689 19935 3723
rect 2053 3621 2087 3655
rect 1409 3553 1443 3587
rect 2513 3553 2547 3587
rect 4445 3553 4479 3587
rect 5641 3553 5675 3587
rect 15577 3553 15611 3587
rect 16304 3553 16338 3587
rect 18777 3553 18811 3587
rect 26525 3553 26559 3587
rect 4537 3485 4571 3519
rect 4629 3485 4663 3519
rect 5917 3485 5951 3519
rect 14657 3485 14691 3519
rect 16037 3485 16071 3519
rect 18521 3485 18555 3519
rect 1593 3349 1627 3383
rect 2697 3349 2731 3383
rect 17417 3349 17451 3383
rect 26709 3349 26743 3383
rect 2513 3145 2547 3179
rect 4077 3145 4111 3179
rect 6193 3145 6227 3179
rect 13277 3145 13311 3179
rect 14473 3145 14507 3179
rect 16129 3145 16163 3179
rect 17785 3145 17819 3179
rect 18797 3145 18831 3179
rect 18981 3145 19015 3179
rect 21373 3145 21407 3179
rect 27261 3145 27295 3179
rect 3985 3077 4019 3111
rect 5181 3077 5215 3111
rect 16497 3077 16531 3111
rect 19993 3077 20027 3111
rect 4629 3009 4663 3043
rect 5457 3009 5491 3043
rect 5825 3009 5859 3043
rect 19533 3009 19567 3043
rect 1593 2941 1627 2975
rect 2697 2941 2731 2975
rect 3617 2941 3651 2975
rect 4537 2941 4571 2975
rect 8677 2941 8711 2975
rect 9413 2941 9447 2975
rect 12449 2941 12483 2975
rect 13737 2941 13771 2975
rect 18521 2941 18555 2975
rect 19349 2941 19383 2975
rect 19441 2941 19475 2975
rect 20545 2941 20579 2975
rect 23673 2941 23707 2975
rect 24409 2941 24443 2975
rect 26341 2941 26375 2975
rect 26893 2941 26927 2975
rect 27445 2941 27479 2975
rect 27997 2941 28031 2975
rect 2237 2873 2271 2907
rect 8953 2873 8987 2907
rect 12725 2873 12759 2907
rect 14013 2873 14047 2907
rect 20821 2873 20855 2907
rect 23949 2873 23983 2907
rect 1777 2805 1811 2839
rect 2881 2805 2915 2839
rect 4445 2805 4479 2839
rect 26525 2805 26559 2839
rect 27629 2805 27663 2839
rect 3801 2601 3835 2635
rect 4905 2601 4939 2635
rect 11161 2601 11195 2635
rect 18061 2601 18095 2635
rect 19073 2601 19107 2635
rect 21925 2601 21959 2635
rect 23489 2601 23523 2635
rect 5825 2533 5859 2567
rect 13461 2533 13495 2567
rect 18613 2533 18647 2567
rect 1501 2465 1535 2499
rect 1768 2465 1802 2499
rect 3157 2465 3191 2499
rect 4077 2465 4111 2499
rect 5549 2465 5583 2499
rect 6285 2465 6319 2499
rect 6929 2465 6963 2499
rect 7665 2465 7699 2499
rect 10333 2465 10367 2499
rect 13185 2465 13219 2499
rect 13921 2465 13955 2499
rect 15761 2465 15795 2499
rect 16497 2465 16531 2499
rect 18337 2465 18371 2499
rect 19625 2465 19659 2499
rect 20361 2465 20395 2499
rect 21189 2465 21223 2499
rect 22661 2465 22695 2499
rect 25697 2465 25731 2499
rect 26249 2465 26283 2499
rect 4353 2397 4387 2431
rect 7113 2397 7147 2431
rect 10609 2397 10643 2431
rect 16037 2397 16071 2431
rect 19809 2397 19843 2431
rect 21465 2397 21499 2431
rect 22937 2397 22971 2431
rect 2881 2329 2915 2363
rect 5181 2261 5215 2295
rect 25881 2261 25915 2295
rect 27077 2261 27111 2295
<< metal1 >>
rect 3418 22176 3424 22228
rect 3476 22216 3482 22228
rect 8294 22216 8300 22228
rect 3476 22188 8300 22216
rect 3476 22176 3482 22188
rect 8294 22176 8300 22188
rect 8352 22176 8358 22228
rect 3050 22108 3056 22160
rect 3108 22148 3114 22160
rect 15654 22148 15660 22160
rect 3108 22120 15660 22148
rect 3108 22108 3114 22120
rect 15654 22108 15660 22120
rect 15712 22108 15718 22160
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 2958 20748 2964 20800
rect 3016 20788 3022 20800
rect 17954 20788 17960 20800
rect 3016 20760 17960 20788
rect 3016 20748 3022 20760
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 21361 20587 21419 20593
rect 21361 20553 21373 20587
rect 21407 20584 21419 20587
rect 22462 20584 22468 20596
rect 21407 20556 22468 20584
rect 21407 20553 21419 20556
rect 21361 20547 21419 20553
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 25777 20383 25835 20389
rect 25777 20349 25789 20383
rect 25823 20380 25835 20383
rect 25823 20352 26464 20380
rect 25823 20349 25835 20352
rect 25777 20343 25835 20349
rect 25958 20244 25964 20256
rect 25919 20216 25964 20244
rect 25958 20204 25964 20216
rect 26016 20204 26022 20256
rect 26436 20253 26464 20352
rect 26421 20247 26479 20253
rect 26421 20213 26433 20247
rect 26467 20244 26479 20247
rect 27798 20244 27804 20256
rect 26467 20216 27804 20244
rect 26467 20213 26479 20216
rect 26421 20207 26479 20213
rect 27798 20204 27804 20216
rect 27856 20204 27862 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 2317 19159 2375 19165
rect 2317 19156 2329 19159
rect 2087 19128 2329 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2317 19125 2329 19128
rect 2363 19156 2375 19159
rect 2590 19156 2596 19168
rect 2363 19128 2596 19156
rect 2363 19125 2375 19128
rect 2317 19119 2375 19125
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 2130 18844 2136 18896
rect 2188 18884 2194 18896
rect 2409 18887 2467 18893
rect 2409 18884 2421 18887
rect 2188 18856 2421 18884
rect 2188 18844 2194 18856
rect 2409 18853 2421 18856
rect 2455 18884 2467 18887
rect 3510 18884 3516 18896
rect 2455 18856 3516 18884
rect 2455 18853 2467 18856
rect 2409 18847 2467 18853
rect 3510 18844 3516 18856
rect 3568 18844 3574 18896
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 2317 18819 2375 18825
rect 2317 18816 2329 18819
rect 1903 18788 2329 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 2317 18785 2329 18788
rect 2363 18816 2375 18819
rect 3602 18816 3608 18828
rect 2363 18788 3608 18816
rect 2363 18785 2375 18788
rect 2317 18779 2375 18785
rect 3602 18776 3608 18788
rect 3660 18776 3666 18828
rect 9582 18776 9588 18828
rect 9640 18816 9646 18828
rect 10117 18819 10175 18825
rect 10117 18816 10129 18819
rect 9640 18788 10129 18816
rect 9640 18776 9646 18788
rect 10117 18785 10129 18788
rect 10163 18785 10175 18819
rect 10117 18779 10175 18785
rect 18868 18819 18926 18825
rect 18868 18785 18880 18819
rect 18914 18816 18926 18819
rect 19150 18816 19156 18828
rect 18914 18788 19156 18816
rect 18914 18785 18926 18788
rect 18868 18779 18926 18785
rect 19150 18776 19156 18788
rect 19208 18776 19214 18828
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 24486 18825 24492 18828
rect 22261 18819 22319 18825
rect 22261 18816 22273 18819
rect 22152 18788 22273 18816
rect 22152 18776 22158 18788
rect 22261 18785 22273 18788
rect 22307 18785 22319 18819
rect 24480 18816 24492 18825
rect 22261 18779 22319 18785
rect 23400 18788 24492 18816
rect 2590 18748 2596 18760
rect 2551 18720 2596 18748
rect 2590 18708 2596 18720
rect 2648 18708 2654 18760
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9824 18720 9873 18748
rect 9824 18708 9830 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 18598 18748 18604 18760
rect 18559 18720 18604 18748
rect 9861 18711 9919 18717
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 22005 18751 22063 18757
rect 22005 18717 22017 18751
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 8202 18680 8208 18692
rect 8163 18652 8208 18680
rect 8202 18640 8208 18652
rect 8260 18640 8266 18692
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 11241 18615 11299 18621
rect 11241 18581 11253 18615
rect 11287 18612 11299 18615
rect 11698 18612 11704 18624
rect 11287 18584 11704 18612
rect 11287 18581 11299 18584
rect 11241 18575 11299 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 12618 18612 12624 18624
rect 12579 18584 12624 18612
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 15105 18615 15163 18621
rect 15105 18581 15117 18615
rect 15151 18612 15163 18615
rect 15286 18612 15292 18624
rect 15151 18584 15292 18612
rect 15151 18581 15163 18584
rect 15105 18575 15163 18581
rect 15286 18572 15292 18584
rect 15344 18572 15350 18624
rect 19978 18612 19984 18624
rect 19939 18584 19984 18612
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 21082 18612 21088 18624
rect 21043 18584 21088 18612
rect 21082 18572 21088 18584
rect 21140 18612 21146 18624
rect 22020 18612 22048 18711
rect 23400 18689 23428 18788
rect 24480 18779 24492 18788
rect 24486 18776 24492 18779
rect 24544 18776 24550 18828
rect 24213 18751 24271 18757
rect 24213 18717 24225 18751
rect 24259 18717 24271 18751
rect 24213 18711 24271 18717
rect 23385 18683 23443 18689
rect 23385 18649 23397 18683
rect 23431 18649 23443 18683
rect 23385 18643 23443 18649
rect 22186 18612 22192 18624
rect 21140 18584 22192 18612
rect 21140 18572 21146 18584
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 24228 18612 24256 18711
rect 24578 18612 24584 18624
rect 24228 18584 24584 18612
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 25590 18612 25596 18624
rect 25551 18584 25596 18612
rect 25590 18572 25596 18584
rect 25648 18572 25654 18624
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 20346 18408 20352 18420
rect 20036 18380 20352 18408
rect 20036 18368 20042 18380
rect 20346 18368 20352 18380
rect 20404 18408 20410 18420
rect 20901 18411 20959 18417
rect 20901 18408 20913 18411
rect 20404 18380 20913 18408
rect 20404 18368 20410 18380
rect 20901 18377 20913 18380
rect 20947 18377 20959 18411
rect 20901 18371 20959 18377
rect 3510 18340 3516 18352
rect 3471 18312 3516 18340
rect 3510 18300 3516 18312
rect 3568 18300 3574 18352
rect 14001 18343 14059 18349
rect 14001 18309 14013 18343
rect 14047 18340 14059 18343
rect 15286 18340 15292 18352
rect 14047 18312 15292 18340
rect 14047 18309 14059 18312
rect 14001 18303 14059 18309
rect 15286 18300 15292 18312
rect 15344 18340 15350 18352
rect 15344 18312 15608 18340
rect 15344 18300 15350 18312
rect 1762 18232 1768 18284
rect 1820 18272 1826 18284
rect 2590 18272 2596 18284
rect 1820 18244 2596 18272
rect 1820 18232 1826 18244
rect 2590 18232 2596 18244
rect 2648 18232 2654 18284
rect 3602 18272 3608 18284
rect 3563 18244 3608 18272
rect 3602 18232 3608 18244
rect 3660 18232 3666 18284
rect 11514 18232 11520 18284
rect 11572 18272 11578 18284
rect 12618 18272 12624 18284
rect 11572 18244 12624 18272
rect 11572 18232 11578 18244
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 15580 18281 15608 18312
rect 18598 18300 18604 18352
rect 18656 18340 18662 18352
rect 19334 18340 19340 18352
rect 18656 18312 19340 18340
rect 18656 18300 18662 18312
rect 19334 18300 19340 18312
rect 19392 18340 19398 18352
rect 20441 18343 20499 18349
rect 20441 18340 20453 18343
rect 19392 18312 20453 18340
rect 19392 18300 19398 18312
rect 20441 18309 20453 18312
rect 20487 18309 20499 18343
rect 20441 18303 20499 18309
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 19150 18272 19156 18284
rect 19111 18244 19156 18272
rect 15565 18235 15623 18241
rect 19150 18232 19156 18244
rect 19208 18272 19214 18284
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 19208 18244 19625 18272
rect 19208 18232 19214 18244
rect 19613 18241 19625 18244
rect 19659 18272 19671 18275
rect 19981 18275 20039 18281
rect 19981 18272 19993 18275
rect 19659 18244 19993 18272
rect 19659 18241 19671 18244
rect 19613 18235 19671 18241
rect 19981 18241 19993 18244
rect 20027 18241 20039 18275
rect 19981 18235 20039 18241
rect 2501 18207 2559 18213
rect 2501 18173 2513 18207
rect 2547 18204 2559 18207
rect 3050 18204 3056 18216
rect 2547 18176 3056 18204
rect 2547 18173 2559 18176
rect 2501 18167 2559 18173
rect 3050 18164 3056 18176
rect 3108 18164 3114 18216
rect 8113 18207 8171 18213
rect 8113 18173 8125 18207
rect 8159 18204 8171 18207
rect 8202 18204 8208 18216
rect 8159 18176 8208 18204
rect 8159 18173 8171 18176
rect 8113 18167 8171 18173
rect 8202 18164 8208 18176
rect 8260 18164 8266 18216
rect 12894 18213 12900 18216
rect 12877 18207 12900 18213
rect 12877 18204 12889 18207
rect 12176 18176 12889 18204
rect 12176 18148 12204 18176
rect 12877 18173 12889 18176
rect 12952 18204 12958 18216
rect 12952 18176 13025 18204
rect 12877 18167 12900 18173
rect 12894 18164 12900 18167
rect 12952 18164 12958 18176
rect 18322 18164 18328 18216
rect 18380 18204 18386 18216
rect 18969 18207 19027 18213
rect 18969 18204 18981 18207
rect 18380 18176 18981 18204
rect 18380 18164 18386 18176
rect 18969 18173 18981 18176
rect 19015 18173 19027 18207
rect 20916 18204 20944 18371
rect 21082 18272 21088 18284
rect 21043 18244 21088 18272
rect 21082 18232 21088 18244
rect 21140 18232 21146 18284
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18272 24363 18275
rect 24486 18272 24492 18284
rect 24351 18244 24492 18272
rect 24351 18241 24363 18244
rect 24305 18235 24363 18241
rect 24486 18232 24492 18244
rect 24544 18272 24550 18284
rect 25038 18272 25044 18284
rect 24544 18244 25044 18272
rect 24544 18232 24550 18244
rect 25038 18232 25044 18244
rect 25096 18232 25102 18284
rect 21341 18207 21399 18213
rect 21341 18204 21353 18207
rect 20916 18176 21353 18204
rect 18969 18167 19027 18173
rect 21341 18173 21353 18176
rect 21387 18173 21399 18207
rect 25225 18207 25283 18213
rect 25225 18204 25237 18207
rect 21341 18167 21399 18173
rect 24872 18176 25237 18204
rect 1949 18139 2007 18145
rect 1949 18105 1961 18139
rect 1995 18136 2007 18139
rect 8021 18139 8079 18145
rect 1995 18108 2452 18136
rect 1995 18105 2007 18108
rect 1949 18099 2007 18105
rect 2038 18068 2044 18080
rect 1999 18040 2044 18068
rect 2038 18028 2044 18040
rect 2096 18028 2102 18080
rect 2424 18077 2452 18108
rect 8021 18105 8033 18139
rect 8067 18136 8079 18139
rect 8358 18139 8416 18145
rect 8358 18136 8370 18139
rect 8067 18108 8370 18136
rect 8067 18105 8079 18108
rect 8021 18099 8079 18105
rect 8358 18105 8370 18108
rect 8404 18136 8416 18139
rect 8570 18136 8576 18148
rect 8404 18108 8576 18136
rect 8404 18105 8416 18108
rect 8358 18099 8416 18105
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 9766 18096 9772 18148
rect 9824 18136 9830 18148
rect 10229 18139 10287 18145
rect 10229 18136 10241 18139
rect 9824 18108 10241 18136
rect 9824 18096 9830 18108
rect 10229 18105 10241 18108
rect 10275 18105 10287 18139
rect 12158 18136 12164 18148
rect 12119 18108 12164 18136
rect 10229 18099 10287 18105
rect 12158 18096 12164 18108
rect 12216 18096 12222 18148
rect 14274 18096 14280 18148
rect 14332 18136 14338 18148
rect 14921 18139 14979 18145
rect 14921 18136 14933 18139
rect 14332 18108 14933 18136
rect 14332 18096 14338 18108
rect 14921 18105 14933 18108
rect 14967 18136 14979 18139
rect 15470 18136 15476 18148
rect 14967 18108 15476 18136
rect 14967 18105 14979 18108
rect 14921 18099 14979 18105
rect 15470 18096 15476 18108
rect 15528 18096 15534 18148
rect 19058 18136 19064 18148
rect 17788 18108 19064 18136
rect 2409 18071 2467 18077
rect 2409 18037 2421 18071
rect 2455 18068 2467 18071
rect 2590 18068 2596 18080
rect 2455 18040 2596 18068
rect 2455 18037 2467 18040
rect 2409 18031 2467 18037
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 3050 18068 3056 18080
rect 3011 18040 3056 18068
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 9493 18071 9551 18077
rect 9493 18037 9505 18071
rect 9539 18068 9551 18071
rect 9582 18068 9588 18080
rect 9539 18040 9588 18068
rect 9539 18037 9551 18040
rect 9493 18031 9551 18037
rect 9582 18028 9588 18040
rect 9640 18068 9646 18080
rect 9861 18071 9919 18077
rect 9861 18068 9873 18071
rect 9640 18040 9873 18068
rect 9640 18028 9646 18040
rect 9861 18037 9873 18040
rect 9907 18037 9919 18071
rect 15010 18068 15016 18080
rect 14971 18040 15016 18068
rect 9861 18031 9919 18037
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 15194 18028 15200 18080
rect 15252 18068 15258 18080
rect 15381 18071 15439 18077
rect 15381 18068 15393 18071
rect 15252 18040 15393 18068
rect 15252 18028 15258 18040
rect 15381 18037 15393 18040
rect 15427 18037 15439 18071
rect 15381 18031 15439 18037
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 17788 18077 17816 18108
rect 19058 18096 19064 18108
rect 19116 18096 19122 18148
rect 17773 18071 17831 18077
rect 17773 18068 17785 18071
rect 16632 18040 17785 18068
rect 16632 18028 16638 18040
rect 17773 18037 17785 18040
rect 17819 18037 17831 18071
rect 17773 18031 17831 18037
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 18417 18071 18475 18077
rect 18417 18068 18429 18071
rect 18380 18040 18429 18068
rect 18380 18028 18386 18040
rect 18417 18037 18429 18040
rect 18463 18037 18475 18071
rect 18417 18031 18475 18037
rect 18601 18071 18659 18077
rect 18601 18037 18613 18071
rect 18647 18068 18659 18071
rect 18874 18068 18880 18080
rect 18647 18040 18880 18068
rect 18647 18037 18659 18040
rect 18601 18031 18659 18037
rect 18874 18028 18880 18040
rect 18932 18028 18938 18080
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 22465 18071 22523 18077
rect 22465 18068 22477 18071
rect 22152 18040 22477 18068
rect 22152 18028 22158 18040
rect 22465 18037 22477 18040
rect 22511 18068 22523 18071
rect 22741 18071 22799 18077
rect 22741 18068 22753 18071
rect 22511 18040 22753 18068
rect 22511 18037 22523 18040
rect 22465 18031 22523 18037
rect 22741 18037 22753 18040
rect 22787 18037 22799 18071
rect 24578 18068 24584 18080
rect 24539 18040 24584 18068
rect 22741 18031 22799 18037
rect 24578 18028 24584 18040
rect 24636 18068 24642 18080
rect 24872 18068 24900 18176
rect 25225 18173 25237 18176
rect 25271 18173 25283 18207
rect 25225 18167 25283 18173
rect 25470 18139 25528 18145
rect 25470 18136 25482 18139
rect 25148 18108 25482 18136
rect 25148 18080 25176 18108
rect 25470 18105 25482 18108
rect 25516 18136 25528 18139
rect 25590 18136 25596 18148
rect 25516 18108 25596 18136
rect 25516 18105 25528 18108
rect 25470 18099 25528 18105
rect 25590 18096 25596 18108
rect 25648 18096 25654 18148
rect 25130 18068 25136 18080
rect 24636 18040 24900 18068
rect 25091 18040 25136 18068
rect 24636 18028 24642 18040
rect 25130 18028 25136 18040
rect 25188 18028 25194 18080
rect 26234 18028 26240 18080
rect 26292 18068 26298 18080
rect 26605 18071 26663 18077
rect 26605 18068 26617 18071
rect 26292 18040 26617 18068
rect 26292 18028 26298 18040
rect 26605 18037 26617 18040
rect 26651 18037 26663 18071
rect 26605 18031 26663 18037
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 12894 17824 12900 17876
rect 12952 17864 12958 17876
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 12952 17836 13001 17864
rect 12952 17824 12958 17836
rect 12989 17833 13001 17836
rect 13035 17833 13047 17867
rect 12989 17827 13047 17833
rect 14369 17867 14427 17873
rect 14369 17833 14381 17867
rect 14415 17864 14427 17867
rect 14642 17864 14648 17876
rect 14415 17836 14648 17864
rect 14415 17833 14427 17836
rect 14369 17827 14427 17833
rect 14642 17824 14648 17836
rect 14700 17864 14706 17876
rect 15010 17864 15016 17876
rect 14700 17836 15016 17864
rect 14700 17824 14706 17836
rect 15010 17824 15016 17836
rect 15068 17824 15074 17876
rect 18601 17867 18659 17873
rect 18601 17833 18613 17867
rect 18647 17864 18659 17867
rect 21269 17867 21327 17873
rect 21269 17864 21281 17867
rect 18647 17836 21281 17864
rect 18647 17833 18659 17836
rect 18601 17827 18659 17833
rect 21269 17833 21281 17836
rect 21315 17833 21327 17867
rect 21269 17827 21327 17833
rect 18874 17756 18880 17808
rect 18932 17796 18938 17808
rect 19061 17799 19119 17805
rect 19061 17796 19073 17799
rect 18932 17768 19073 17796
rect 18932 17756 18938 17768
rect 19061 17765 19073 17768
rect 19107 17765 19119 17799
rect 19061 17759 19119 17765
rect 1762 17688 1768 17740
rect 1820 17728 1826 17740
rect 1929 17731 1987 17737
rect 1929 17728 1941 17731
rect 1820 17700 1941 17728
rect 1820 17688 1826 17700
rect 1929 17697 1941 17700
rect 1975 17697 1987 17731
rect 1929 17691 1987 17697
rect 4430 17688 4436 17740
rect 4488 17728 4494 17740
rect 4873 17731 4931 17737
rect 4873 17728 4885 17731
rect 4488 17700 4885 17728
rect 4488 17688 4494 17700
rect 4873 17697 4885 17700
rect 4919 17697 4931 17731
rect 4873 17691 4931 17697
rect 7009 17731 7067 17737
rect 7009 17697 7021 17731
rect 7055 17728 7067 17731
rect 7742 17728 7748 17740
rect 7055 17700 7748 17728
rect 7055 17697 7067 17700
rect 7009 17691 7067 17697
rect 7742 17688 7748 17700
rect 7800 17728 7806 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7800 17700 8401 17728
rect 7800 17688 7806 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 11865 17731 11923 17737
rect 11865 17728 11877 17731
rect 11756 17700 11877 17728
rect 11756 17688 11762 17700
rect 11865 17697 11877 17700
rect 11911 17697 11923 17731
rect 11865 17691 11923 17697
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 15545 17731 15603 17737
rect 15545 17728 15557 17731
rect 15252 17700 15557 17728
rect 15252 17688 15258 17700
rect 15545 17697 15557 17700
rect 15591 17697 15603 17731
rect 15545 17691 15603 17697
rect 18414 17688 18420 17740
rect 18472 17728 18478 17740
rect 18969 17731 19027 17737
rect 18969 17728 18981 17731
rect 18472 17700 18981 17728
rect 18472 17688 18478 17700
rect 18969 17697 18981 17700
rect 19015 17697 19027 17731
rect 21284 17728 21312 17827
rect 24210 17824 24216 17876
rect 24268 17864 24274 17876
rect 25225 17867 25283 17873
rect 25225 17864 25237 17867
rect 24268 17836 25237 17864
rect 24268 17824 24274 17836
rect 25225 17833 25237 17836
rect 25271 17864 25283 17867
rect 26513 17867 26571 17873
rect 26513 17864 26525 17867
rect 25271 17836 26525 17864
rect 25271 17833 25283 17836
rect 25225 17827 25283 17833
rect 26513 17833 26525 17836
rect 26559 17833 26571 17867
rect 26513 17827 26571 17833
rect 22646 17728 22652 17740
rect 21284 17700 22652 17728
rect 18969 17691 19027 17697
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 24946 17688 24952 17740
rect 25004 17728 25010 17740
rect 26881 17731 26939 17737
rect 25004 17700 25544 17728
rect 25004 17688 25010 17700
rect 1670 17660 1676 17672
rect 1631 17632 1676 17660
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 3786 17620 3792 17672
rect 3844 17660 3850 17672
rect 4617 17663 4675 17669
rect 4617 17660 4629 17663
rect 3844 17632 4629 17660
rect 3844 17620 3850 17632
rect 4617 17629 4629 17632
rect 4663 17629 4675 17663
rect 4617 17623 4675 17629
rect 7650 17620 7656 17672
rect 7708 17660 7714 17672
rect 8481 17663 8539 17669
rect 8481 17660 8493 17663
rect 7708 17632 8493 17660
rect 7708 17620 7714 17632
rect 8481 17629 8493 17632
rect 8527 17629 8539 17663
rect 8481 17623 8539 17629
rect 8496 17592 8524 17623
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 8628 17632 8673 17660
rect 8628 17620 8634 17632
rect 9766 17620 9772 17672
rect 9824 17660 9830 17672
rect 11514 17660 11520 17672
rect 9824 17632 11520 17660
rect 9824 17620 9830 17632
rect 11514 17620 11520 17632
rect 11572 17660 11578 17672
rect 11609 17663 11667 17669
rect 11609 17660 11621 17663
rect 11572 17632 11621 17660
rect 11572 17620 11578 17632
rect 11609 17629 11621 17632
rect 11655 17629 11667 17663
rect 15286 17660 15292 17672
rect 15247 17632 15292 17660
rect 11609 17623 11667 17629
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 17586 17660 17592 17672
rect 17547 17632 17592 17660
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 19242 17660 19248 17672
rect 19203 17632 19248 17660
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 21358 17660 21364 17672
rect 21319 17632 21364 17660
rect 21358 17620 21364 17632
rect 21416 17620 21422 17672
rect 21542 17660 21548 17672
rect 21455 17632 21548 17660
rect 21542 17620 21548 17632
rect 21600 17660 21606 17672
rect 22002 17660 22008 17672
rect 21600 17632 22008 17660
rect 21600 17620 21606 17632
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 25314 17660 25320 17672
rect 25275 17632 25320 17660
rect 25314 17620 25320 17632
rect 25372 17620 25378 17672
rect 25516 17669 25544 17700
rect 26881 17697 26893 17731
rect 26927 17728 26939 17731
rect 27154 17728 27160 17740
rect 26927 17700 27160 17728
rect 26927 17697 26939 17700
rect 26881 17691 26939 17697
rect 27154 17688 27160 17700
rect 27212 17688 27218 17740
rect 25501 17663 25559 17669
rect 25501 17629 25513 17663
rect 25547 17660 25559 17663
rect 26142 17660 26148 17672
rect 25547 17632 26148 17660
rect 25547 17629 25559 17632
rect 25501 17623 25559 17629
rect 26142 17620 26148 17632
rect 26200 17620 26206 17672
rect 26786 17620 26792 17672
rect 26844 17660 26850 17672
rect 26973 17663 27031 17669
rect 26973 17660 26985 17663
rect 26844 17632 26985 17660
rect 26844 17620 26850 17632
rect 26973 17629 26985 17632
rect 27019 17629 27031 17663
rect 26973 17623 27031 17629
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17629 27123 17663
rect 27065 17623 27123 17629
rect 9490 17592 9496 17604
rect 8496 17564 9496 17592
rect 9490 17552 9496 17564
rect 9548 17552 9554 17604
rect 18509 17595 18567 17601
rect 18509 17561 18521 17595
rect 18555 17592 18567 17595
rect 19150 17592 19156 17604
rect 18555 17564 19156 17592
rect 18555 17561 18567 17564
rect 18509 17555 18567 17561
rect 19150 17552 19156 17564
rect 19208 17552 19214 17604
rect 22097 17595 22155 17601
rect 22097 17561 22109 17595
rect 22143 17592 22155 17595
rect 22186 17592 22192 17604
rect 22143 17564 22192 17592
rect 22143 17561 22155 17564
rect 22097 17555 22155 17561
rect 22186 17552 22192 17564
rect 22244 17592 22250 17604
rect 23566 17592 23572 17604
rect 22244 17564 23572 17592
rect 22244 17552 22250 17564
rect 23566 17552 23572 17564
rect 23624 17592 23630 17604
rect 24578 17592 24584 17604
rect 23624 17564 24584 17592
rect 23624 17552 23630 17564
rect 24578 17552 24584 17564
rect 24636 17592 24642 17604
rect 25869 17595 25927 17601
rect 25869 17592 25881 17595
rect 24636 17564 25881 17592
rect 24636 17552 24642 17564
rect 25869 17561 25881 17564
rect 25915 17561 25927 17595
rect 25869 17555 25927 17561
rect 26326 17552 26332 17604
rect 26384 17592 26390 17604
rect 27080 17592 27108 17623
rect 26384 17564 27108 17592
rect 26384 17552 26390 17564
rect 2682 17484 2688 17536
rect 2740 17524 2746 17536
rect 3053 17527 3111 17533
rect 3053 17524 3065 17527
rect 2740 17496 3065 17524
rect 2740 17484 2746 17496
rect 3053 17493 3065 17496
rect 3099 17524 3111 17527
rect 4430 17524 4436 17536
rect 3099 17496 4436 17524
rect 3099 17493 3111 17496
rect 3053 17487 3111 17493
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 5997 17527 6055 17533
rect 5997 17524 6009 17527
rect 5592 17496 6009 17524
rect 5592 17484 5598 17496
rect 5997 17493 6009 17496
rect 6043 17493 6055 17527
rect 5997 17487 6055 17493
rect 8021 17527 8079 17533
rect 8021 17493 8033 17527
rect 8067 17524 8079 17527
rect 8570 17524 8576 17536
rect 8067 17496 8576 17524
rect 8067 17493 8079 17496
rect 8021 17487 8079 17493
rect 8570 17484 8576 17496
rect 8628 17524 8634 17536
rect 9033 17527 9091 17533
rect 9033 17524 9045 17527
rect 8628 17496 9045 17524
rect 8628 17484 8634 17496
rect 9033 17493 9045 17496
rect 9079 17493 9091 17527
rect 10042 17524 10048 17536
rect 10003 17496 10048 17524
rect 9033 17487 9091 17493
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 10318 17524 10324 17536
rect 10279 17496 10324 17524
rect 10318 17484 10324 17496
rect 10376 17484 10382 17536
rect 15102 17524 15108 17536
rect 15063 17496 15108 17524
rect 15102 17484 15108 17496
rect 15160 17484 15166 17536
rect 16666 17524 16672 17536
rect 16627 17496 16672 17524
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 20901 17527 20959 17533
rect 20901 17493 20913 17527
rect 20947 17524 20959 17527
rect 21450 17524 21456 17536
rect 20947 17496 21456 17524
rect 20947 17493 20959 17496
rect 20901 17487 20959 17493
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 24854 17524 24860 17536
rect 24815 17496 24860 17524
rect 24854 17484 24860 17496
rect 24912 17484 24918 17536
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 1670 17320 1676 17332
rect 1452 17292 1676 17320
rect 1452 17280 1458 17292
rect 1670 17280 1676 17292
rect 1728 17320 1734 17332
rect 3786 17320 3792 17332
rect 1728 17292 3792 17320
rect 1728 17280 1734 17292
rect 3786 17280 3792 17292
rect 3844 17280 3850 17332
rect 4430 17320 4436 17332
rect 4391 17292 4436 17320
rect 4430 17280 4436 17292
rect 4488 17280 4494 17332
rect 7742 17320 7748 17332
rect 7703 17292 7748 17320
rect 7742 17280 7748 17292
rect 7800 17280 7806 17332
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 11977 17323 12035 17329
rect 11977 17320 11989 17323
rect 11572 17292 11989 17320
rect 11572 17280 11578 17292
rect 11977 17289 11989 17292
rect 12023 17289 12035 17323
rect 11977 17283 12035 17289
rect 17865 17323 17923 17329
rect 17865 17289 17877 17323
rect 17911 17320 17923 17323
rect 18414 17320 18420 17332
rect 17911 17292 18420 17320
rect 17911 17289 17923 17292
rect 17865 17283 17923 17289
rect 18414 17280 18420 17292
rect 18472 17280 18478 17332
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 19521 17323 19579 17329
rect 19521 17320 19533 17323
rect 19300 17292 19533 17320
rect 19300 17280 19306 17292
rect 19521 17289 19533 17292
rect 19567 17320 19579 17323
rect 20346 17320 20352 17332
rect 19567 17292 20352 17320
rect 19567 17289 19579 17292
rect 19521 17283 19579 17289
rect 20346 17280 20352 17292
rect 20404 17280 20410 17332
rect 20901 17323 20959 17329
rect 20901 17289 20913 17323
rect 20947 17320 20959 17323
rect 21358 17320 21364 17332
rect 20947 17292 21364 17320
rect 20947 17289 20959 17292
rect 20901 17283 20959 17289
rect 21358 17280 21364 17292
rect 21416 17320 21422 17332
rect 22281 17323 22339 17329
rect 22281 17320 22293 17323
rect 21416 17292 22293 17320
rect 21416 17280 21422 17292
rect 22281 17289 22293 17292
rect 22327 17289 22339 17323
rect 22646 17320 22652 17332
rect 22607 17292 22652 17320
rect 22281 17283 22339 17289
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 24210 17320 24216 17332
rect 24171 17292 24216 17320
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 24581 17323 24639 17329
rect 24581 17289 24593 17323
rect 24627 17320 24639 17323
rect 25314 17320 25320 17332
rect 24627 17292 25320 17320
rect 24627 17289 24639 17292
rect 24581 17283 24639 17289
rect 25314 17280 25320 17292
rect 25372 17320 25378 17332
rect 25777 17323 25835 17329
rect 25777 17320 25789 17323
rect 25372 17292 25789 17320
rect 25372 17280 25378 17292
rect 25777 17289 25789 17292
rect 25823 17289 25835 17323
rect 25777 17283 25835 17289
rect 3053 17255 3111 17261
rect 3053 17252 3065 17255
rect 2516 17224 3065 17252
rect 2038 17144 2044 17196
rect 2096 17184 2102 17196
rect 2516 17193 2544 17224
rect 3053 17221 3065 17224
rect 3099 17221 3111 17255
rect 3804 17252 3832 17280
rect 5442 17252 5448 17264
rect 3804 17224 5448 17252
rect 3053 17215 3111 17221
rect 5442 17212 5448 17224
rect 5500 17252 5506 17264
rect 5905 17255 5963 17261
rect 5905 17252 5917 17255
rect 5500 17224 5917 17252
rect 5500 17212 5506 17224
rect 5905 17221 5917 17224
rect 5951 17221 5963 17255
rect 5905 17215 5963 17221
rect 7377 17255 7435 17261
rect 7377 17221 7389 17255
rect 7423 17252 7435 17255
rect 8478 17252 8484 17264
rect 7423 17224 8484 17252
rect 7423 17221 7435 17224
rect 7377 17215 7435 17221
rect 8478 17212 8484 17224
rect 8536 17212 8542 17264
rect 9861 17255 9919 17261
rect 9861 17221 9873 17255
rect 9907 17252 9919 17255
rect 11609 17255 11667 17261
rect 11609 17252 11621 17255
rect 9907 17224 11621 17252
rect 9907 17221 9919 17224
rect 9861 17215 9919 17221
rect 2501 17187 2559 17193
rect 2501 17184 2513 17187
rect 2096 17156 2513 17184
rect 2096 17144 2102 17156
rect 2501 17153 2513 17156
rect 2547 17153 2559 17187
rect 2682 17184 2688 17196
rect 2643 17156 2688 17184
rect 2501 17147 2559 17153
rect 2682 17144 2688 17156
rect 2740 17184 2746 17196
rect 2958 17184 2964 17196
rect 2740 17156 2964 17184
rect 2740 17144 2746 17156
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17184 4859 17187
rect 5534 17184 5540 17196
rect 4847 17156 5540 17184
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17184 8907 17187
rect 9033 17187 9091 17193
rect 9033 17184 9045 17187
rect 8895 17156 9045 17184
rect 8895 17153 8907 17156
rect 8849 17147 8907 17153
rect 9033 17153 9045 17156
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 10042 17144 10048 17196
rect 10100 17184 10106 17196
rect 10520 17193 10548 17224
rect 11609 17221 11621 17224
rect 11655 17252 11667 17255
rect 11698 17252 11704 17264
rect 11655 17224 11704 17252
rect 11655 17221 11667 17224
rect 11609 17215 11667 17221
rect 11698 17212 11704 17224
rect 11756 17212 11762 17264
rect 13722 17212 13728 17264
rect 13780 17252 13786 17264
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 13780 17224 14289 17252
rect 13780 17212 13786 17224
rect 14277 17221 14289 17224
rect 14323 17221 14335 17255
rect 14277 17215 14335 17221
rect 10413 17187 10471 17193
rect 10413 17184 10425 17187
rect 10100 17156 10425 17184
rect 10100 17144 10106 17156
rect 10413 17153 10425 17156
rect 10459 17153 10471 17187
rect 10413 17147 10471 17153
rect 10505 17187 10563 17193
rect 10505 17153 10517 17187
rect 10551 17153 10563 17187
rect 10505 17147 10563 17153
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17184 14243 17187
rect 14918 17184 14924 17196
rect 14231 17156 14924 17184
rect 14231 17153 14243 17156
rect 14185 17147 14243 17153
rect 14918 17144 14924 17156
rect 14976 17144 14982 17196
rect 15102 17144 15108 17196
rect 15160 17184 15166 17196
rect 15841 17187 15899 17193
rect 15841 17184 15853 17187
rect 15160 17156 15853 17184
rect 15160 17144 15166 17156
rect 15841 17153 15853 17156
rect 15887 17153 15899 17187
rect 15841 17147 15899 17153
rect 18138 17144 18144 17196
rect 18196 17184 18202 17196
rect 18325 17187 18383 17193
rect 18325 17184 18337 17187
rect 18196 17156 18337 17184
rect 18196 17144 18202 17156
rect 18325 17153 18337 17156
rect 18371 17184 18383 17187
rect 18877 17187 18935 17193
rect 18877 17184 18889 17187
rect 18371 17156 18889 17184
rect 18371 17153 18383 17156
rect 18325 17147 18383 17153
rect 18877 17153 18889 17156
rect 18923 17184 18935 17187
rect 18966 17184 18972 17196
rect 18923 17156 18972 17184
rect 18923 17153 18935 17156
rect 18877 17147 18935 17153
rect 18966 17144 18972 17156
rect 19024 17144 19030 17196
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19150 17184 19156 17196
rect 19107 17156 19156 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 19150 17144 19156 17156
rect 19208 17184 19214 17196
rect 19426 17184 19432 17196
rect 19208 17156 19432 17184
rect 19208 17144 19214 17156
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 20364 17184 20392 17280
rect 20809 17255 20867 17261
rect 20809 17221 20821 17255
rect 20855 17252 20867 17255
rect 21542 17252 21548 17264
rect 20855 17224 21548 17252
rect 20855 17221 20867 17224
rect 20809 17215 20867 17221
rect 21542 17212 21548 17224
rect 21600 17212 21606 17264
rect 24946 17252 24952 17264
rect 24907 17224 24952 17252
rect 24946 17212 24952 17224
rect 25004 17212 25010 17264
rect 26786 17252 26792 17264
rect 26747 17224 26792 17252
rect 26786 17212 26792 17224
rect 26844 17212 26850 17264
rect 21453 17187 21511 17193
rect 21453 17184 21465 17187
rect 20364 17156 21465 17184
rect 21453 17153 21465 17156
rect 21499 17153 21511 17187
rect 26326 17184 26332 17196
rect 26287 17156 26332 17184
rect 21453 17147 21511 17153
rect 26326 17144 26332 17156
rect 26384 17144 26390 17196
rect 1946 17076 1952 17128
rect 2004 17116 2010 17128
rect 2409 17119 2467 17125
rect 2409 17116 2421 17119
rect 2004 17088 2421 17116
rect 2004 17076 2010 17088
rect 2409 17085 2421 17088
rect 2455 17116 2467 17119
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 2455 17088 3433 17116
rect 2455 17085 2467 17088
rect 2409 17079 2467 17085
rect 3421 17085 3433 17088
rect 3467 17085 3479 17119
rect 8570 17116 8576 17128
rect 8531 17088 8576 17116
rect 3421 17079 3479 17085
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 14642 17116 14648 17128
rect 14603 17088 14648 17116
rect 14642 17076 14648 17088
rect 14700 17076 14706 17128
rect 20073 17119 20131 17125
rect 20073 17085 20085 17119
rect 20119 17116 20131 17119
rect 21358 17116 21364 17128
rect 20119 17088 21364 17116
rect 20119 17085 20131 17088
rect 20073 17079 20131 17085
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 25130 17076 25136 17128
rect 25188 17116 25194 17128
rect 25317 17119 25375 17125
rect 25317 17116 25329 17119
rect 25188 17088 25329 17116
rect 25188 17076 25194 17088
rect 25317 17085 25329 17088
rect 25363 17116 25375 17119
rect 26344 17116 26372 17144
rect 25363 17088 26372 17116
rect 25363 17085 25375 17088
rect 25317 17079 25375 17085
rect 5258 17048 5264 17060
rect 2056 17020 5264 17048
rect 1762 16980 1768 16992
rect 1723 16952 1768 16980
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 2056 16989 2084 17020
rect 5258 17008 5264 17020
rect 5316 17008 5322 17060
rect 10318 17048 10324 17060
rect 8220 17020 10324 17048
rect 2041 16983 2099 16989
rect 2041 16949 2053 16983
rect 2087 16949 2099 16983
rect 4890 16980 4896 16992
rect 4851 16952 4896 16980
rect 2041 16943 2099 16949
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 5350 16980 5356 16992
rect 5311 16952 5356 16980
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 7650 16940 7656 16992
rect 7708 16980 7714 16992
rect 8220 16989 8248 17020
rect 10318 17008 10324 17020
rect 10376 17008 10382 17060
rect 21266 17048 21272 17060
rect 21179 17020 21272 17048
rect 21266 17008 21272 17020
rect 21324 17048 21330 17060
rect 21913 17051 21971 17057
rect 21913 17048 21925 17051
rect 21324 17020 21925 17048
rect 21324 17008 21330 17020
rect 21913 17017 21925 17020
rect 21959 17017 21971 17051
rect 26234 17048 26240 17060
rect 26195 17020 26240 17048
rect 21913 17011 21971 17017
rect 26234 17008 26240 17020
rect 26292 17048 26298 17060
rect 29178 17048 29184 17060
rect 26292 17020 29184 17048
rect 26292 17008 26298 17020
rect 29178 17008 29184 17020
rect 29236 17008 29242 17060
rect 8021 16983 8079 16989
rect 8021 16980 8033 16983
rect 7708 16952 8033 16980
rect 7708 16940 7714 16952
rect 8021 16949 8033 16952
rect 8067 16949 8079 16983
rect 8021 16943 8079 16949
rect 8205 16983 8263 16989
rect 8205 16949 8217 16983
rect 8251 16949 8263 16983
rect 8662 16980 8668 16992
rect 8623 16952 8668 16980
rect 8205 16943 8263 16949
rect 8662 16940 8668 16952
rect 8720 16940 8726 16992
rect 9033 16983 9091 16989
rect 9033 16949 9045 16983
rect 9079 16980 9091 16983
rect 9309 16983 9367 16989
rect 9309 16980 9321 16983
rect 9079 16952 9321 16980
rect 9079 16949 9091 16952
rect 9033 16943 9091 16949
rect 9309 16949 9321 16952
rect 9355 16980 9367 16983
rect 9582 16980 9588 16992
rect 9355 16952 9588 16980
rect 9355 16949 9367 16952
rect 9309 16943 9367 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 9953 16983 10011 16989
rect 9953 16949 9965 16983
rect 9999 16980 10011 16983
rect 10686 16980 10692 16992
rect 9999 16952 10692 16980
rect 9999 16949 10011 16952
rect 9953 16943 10011 16949
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 14734 16980 14740 16992
rect 14695 16952 14740 16980
rect 14734 16940 14740 16952
rect 14792 16940 14798 16992
rect 15194 16940 15200 16992
rect 15252 16980 15258 16992
rect 15289 16983 15347 16989
rect 15289 16980 15301 16983
rect 15252 16952 15301 16980
rect 15252 16940 15258 16952
rect 15289 16949 15301 16952
rect 15335 16949 15347 16983
rect 15289 16943 15347 16949
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 15749 16983 15807 16989
rect 15749 16980 15761 16983
rect 15436 16952 15761 16980
rect 15436 16940 15442 16952
rect 15749 16949 15761 16952
rect 15795 16980 15807 16983
rect 16298 16980 16304 16992
rect 15795 16952 16304 16980
rect 15795 16949 15807 16952
rect 15749 16943 15807 16949
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 18782 16980 18788 16992
rect 18743 16952 18788 16980
rect 18782 16940 18788 16952
rect 18840 16940 18846 16992
rect 25685 16983 25743 16989
rect 25685 16949 25697 16983
rect 25731 16980 25743 16983
rect 26145 16983 26203 16989
rect 26145 16980 26157 16983
rect 25731 16952 26157 16980
rect 25731 16949 25743 16952
rect 25685 16943 25743 16949
rect 26145 16949 26157 16952
rect 26191 16980 26203 16983
rect 26418 16980 26424 16992
rect 26191 16952 26424 16980
rect 26191 16949 26203 16952
rect 26145 16943 26203 16949
rect 26418 16940 26424 16952
rect 26476 16940 26482 16992
rect 27154 16980 27160 16992
rect 27115 16952 27160 16980
rect 27154 16940 27160 16952
rect 27212 16940 27218 16992
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 4893 16779 4951 16785
rect 4893 16776 4905 16779
rect 2455 16748 4905 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 4893 16745 4905 16748
rect 4939 16776 4951 16779
rect 5350 16776 5356 16788
rect 4939 16748 5356 16776
rect 4939 16745 4951 16748
rect 4893 16739 4951 16745
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 8662 16776 8668 16788
rect 8067 16748 8668 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 8662 16736 8668 16748
rect 8720 16776 8726 16788
rect 9033 16779 9091 16785
rect 9033 16776 9045 16779
rect 8720 16748 9045 16776
rect 8720 16736 8726 16748
rect 9033 16745 9045 16748
rect 9079 16745 9091 16779
rect 9033 16739 9091 16745
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16776 9735 16779
rect 10042 16776 10048 16788
rect 9723 16748 10048 16776
rect 9723 16745 9735 16748
rect 9677 16739 9735 16745
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 11241 16779 11299 16785
rect 11241 16745 11253 16779
rect 11287 16745 11299 16779
rect 11606 16776 11612 16788
rect 11567 16748 11612 16776
rect 11241 16739 11299 16745
rect 1765 16711 1823 16717
rect 1765 16677 1777 16711
rect 1811 16708 1823 16711
rect 2682 16708 2688 16720
rect 1811 16680 2688 16708
rect 1811 16677 1823 16680
rect 1765 16671 1823 16677
rect 2682 16668 2688 16680
rect 2740 16708 2746 16720
rect 2777 16711 2835 16717
rect 2777 16708 2789 16711
rect 2740 16680 2789 16708
rect 2740 16668 2746 16680
rect 2777 16677 2789 16680
rect 2823 16677 2835 16711
rect 5258 16708 5264 16720
rect 5219 16680 5264 16708
rect 2777 16671 2835 16677
rect 5258 16668 5264 16680
rect 5316 16668 5322 16720
rect 5534 16668 5540 16720
rect 5592 16708 5598 16720
rect 5690 16711 5748 16717
rect 5690 16708 5702 16711
rect 5592 16680 5702 16708
rect 5592 16668 5598 16680
rect 5690 16677 5702 16680
rect 5736 16677 5748 16711
rect 9490 16708 9496 16720
rect 9403 16680 9496 16708
rect 5690 16671 5748 16677
rect 9490 16668 9496 16680
rect 9548 16708 9554 16720
rect 10137 16711 10195 16717
rect 10137 16708 10149 16711
rect 9548 16680 10149 16708
rect 9548 16668 9554 16680
rect 10137 16677 10149 16680
rect 10183 16677 10195 16711
rect 10137 16671 10195 16677
rect 2406 16600 2412 16652
rect 2464 16640 2470 16652
rect 2869 16643 2927 16649
rect 2869 16640 2881 16643
rect 2464 16612 2881 16640
rect 2464 16600 2470 16612
rect 2869 16609 2881 16612
rect 2915 16640 2927 16643
rect 4062 16640 4068 16652
rect 2915 16612 4068 16640
rect 2915 16609 2927 16612
rect 2869 16603 2927 16609
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 8294 16640 8300 16652
rect 8207 16612 8300 16640
rect 2958 16572 2964 16584
rect 2919 16544 2964 16572
rect 2958 16532 2964 16544
rect 3016 16532 3022 16584
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 8220 16572 8248 16612
rect 8294 16600 8300 16612
rect 8352 16640 8358 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 8352 16612 8401 16640
rect 8352 16600 8358 16612
rect 8389 16609 8401 16612
rect 8435 16609 8447 16643
rect 8389 16603 8447 16609
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 8662 16640 8668 16652
rect 8527 16612 8668 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9600 16612 10057 16640
rect 8570 16572 8576 16584
rect 8168 16544 8248 16572
rect 8531 16544 8576 16572
rect 8168 16532 8174 16544
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 9122 16532 9128 16584
rect 9180 16572 9186 16584
rect 9600 16572 9628 16612
rect 10045 16609 10057 16612
rect 10091 16640 10103 16643
rect 11256 16640 11284 16739
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 14369 16779 14427 16785
rect 14369 16745 14381 16779
rect 14415 16776 14427 16779
rect 14734 16776 14740 16788
rect 14415 16748 14740 16776
rect 14415 16745 14427 16748
rect 14369 16739 14427 16745
rect 14734 16736 14740 16748
rect 14792 16776 14798 16788
rect 15289 16779 15347 16785
rect 15289 16776 15301 16779
rect 14792 16748 15301 16776
rect 14792 16736 14798 16748
rect 15289 16745 15301 16748
rect 15335 16745 15347 16779
rect 15289 16739 15347 16745
rect 15749 16779 15807 16785
rect 15749 16745 15761 16779
rect 15795 16776 15807 16779
rect 15930 16776 15936 16788
rect 15795 16748 15936 16776
rect 15795 16745 15807 16748
rect 15749 16739 15807 16745
rect 15654 16708 15660 16720
rect 15615 16680 15660 16708
rect 15654 16668 15660 16680
rect 15712 16668 15718 16720
rect 11698 16640 11704 16652
rect 10091 16612 11284 16640
rect 11659 16612 11704 16640
rect 10091 16609 10103 16612
rect 10045 16603 10103 16609
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 15764 16640 15792 16739
rect 15930 16736 15936 16748
rect 15988 16736 15994 16788
rect 17586 16736 17592 16788
rect 17644 16776 17650 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 17644 16748 18429 16776
rect 17644 16736 17650 16748
rect 18417 16745 18429 16748
rect 18463 16776 18475 16779
rect 18782 16776 18788 16788
rect 18463 16748 18788 16776
rect 18463 16745 18475 16748
rect 18417 16739 18475 16745
rect 18782 16736 18788 16748
rect 18840 16736 18846 16788
rect 18874 16736 18880 16788
rect 18932 16776 18938 16788
rect 21177 16779 21235 16785
rect 18932 16748 18977 16776
rect 18932 16736 18938 16748
rect 21177 16745 21189 16779
rect 21223 16776 21235 16779
rect 21266 16776 21272 16788
rect 21223 16748 21272 16776
rect 21223 16745 21235 16748
rect 21177 16739 21235 16745
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 26513 16779 26571 16785
rect 26513 16745 26525 16779
rect 26559 16776 26571 16779
rect 27154 16776 27160 16788
rect 26559 16748 27160 16776
rect 26559 16745 26571 16748
rect 26513 16739 26571 16745
rect 27154 16736 27160 16748
rect 27212 16736 27218 16788
rect 23474 16668 23480 16720
rect 23532 16708 23538 16720
rect 23744 16711 23802 16717
rect 23744 16708 23756 16711
rect 23532 16680 23756 16708
rect 23532 16668 23538 16680
rect 23744 16677 23756 16680
rect 23790 16708 23802 16711
rect 24946 16708 24952 16720
rect 23790 16680 24952 16708
rect 23790 16677 23802 16680
rect 23744 16671 23802 16677
rect 24946 16668 24952 16680
rect 25004 16708 25010 16720
rect 25406 16708 25412 16720
rect 25004 16680 25412 16708
rect 25004 16668 25010 16680
rect 25406 16668 25412 16680
rect 25464 16668 25470 16720
rect 15120 16612 15792 16640
rect 9180 16544 9628 16572
rect 9180 16532 9186 16544
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 10318 16572 10324 16584
rect 9732 16544 10324 16572
rect 9732 16532 9738 16544
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 11885 16575 11943 16581
rect 11885 16541 11897 16575
rect 11931 16572 11943 16575
rect 11974 16572 11980 16584
rect 11931 16544 11980 16572
rect 11931 16541 11943 16544
rect 11885 16535 11943 16541
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 15010 16532 15016 16584
rect 15068 16572 15074 16584
rect 15120 16572 15148 16612
rect 20806 16600 20812 16652
rect 20864 16640 20870 16652
rect 21266 16640 21272 16652
rect 20864 16612 21272 16640
rect 20864 16600 20870 16612
rect 21266 16600 21272 16612
rect 21324 16640 21330 16652
rect 21545 16643 21603 16649
rect 21545 16640 21557 16643
rect 21324 16612 21557 16640
rect 21324 16600 21330 16612
rect 21545 16609 21557 16612
rect 21591 16609 21603 16643
rect 22189 16643 22247 16649
rect 22189 16640 22201 16643
rect 21545 16603 21603 16609
rect 22112 16612 22201 16640
rect 15068 16544 15148 16572
rect 15841 16575 15899 16581
rect 15068 16532 15074 16544
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 21634 16572 21640 16584
rect 21595 16544 21640 16572
rect 15841 16535 15899 16541
rect 1854 16464 1860 16516
rect 1912 16504 1918 16516
rect 2133 16507 2191 16513
rect 2133 16504 2145 16507
rect 1912 16476 2145 16504
rect 1912 16464 1918 16476
rect 2133 16473 2145 16476
rect 2179 16504 2191 16507
rect 2976 16504 3004 16532
rect 2179 16476 3004 16504
rect 2179 16473 2191 16476
rect 2133 16467 2191 16473
rect 15194 16464 15200 16516
rect 15252 16504 15258 16516
rect 15856 16504 15884 16535
rect 21634 16532 21640 16544
rect 21692 16532 21698 16584
rect 21729 16575 21787 16581
rect 21729 16541 21741 16575
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 15252 16476 15884 16504
rect 15252 16464 15258 16476
rect 21542 16464 21548 16516
rect 21600 16504 21606 16516
rect 21744 16504 21772 16535
rect 21818 16532 21824 16584
rect 21876 16572 21882 16584
rect 22112 16572 22140 16612
rect 22189 16609 22201 16612
rect 22235 16609 22247 16643
rect 23566 16640 23572 16652
rect 22189 16603 22247 16609
rect 23492 16612 23572 16640
rect 23492 16581 23520 16612
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 21876 16544 22140 16572
rect 23477 16575 23535 16581
rect 21876 16532 21882 16544
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 25777 16507 25835 16513
rect 25777 16504 25789 16507
rect 21600 16476 21772 16504
rect 24412 16476 25789 16504
rect 21600 16464 21606 16476
rect 6822 16436 6828 16448
rect 6783 16408 6828 16436
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 13354 16436 13360 16448
rect 13315 16408 13360 16436
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 19702 16396 19708 16448
rect 19760 16436 19766 16448
rect 24412 16436 24440 16476
rect 25777 16473 25789 16476
rect 25823 16504 25835 16507
rect 26234 16504 26240 16516
rect 25823 16476 26240 16504
rect 25823 16473 25835 16476
rect 25777 16467 25835 16473
rect 26234 16464 26240 16476
rect 26292 16464 26298 16516
rect 19760 16408 24440 16436
rect 19760 16396 19766 16408
rect 24670 16396 24676 16448
rect 24728 16436 24734 16448
rect 24857 16439 24915 16445
rect 24857 16436 24869 16439
rect 24728 16408 24869 16436
rect 24728 16396 24734 16408
rect 24857 16405 24869 16408
rect 24903 16405 24915 16439
rect 24857 16399 24915 16405
rect 27065 16439 27123 16445
rect 27065 16405 27077 16439
rect 27111 16436 27123 16439
rect 27154 16436 27160 16448
rect 27111 16408 27160 16436
rect 27111 16405 27123 16408
rect 27065 16399 27123 16405
rect 27154 16396 27160 16408
rect 27212 16396 27218 16448
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 1854 16232 1860 16244
rect 1815 16204 1860 16232
rect 1854 16192 1860 16204
rect 1912 16192 1918 16244
rect 2682 16232 2688 16244
rect 2643 16204 2688 16232
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 4062 16232 4068 16244
rect 4023 16204 4068 16232
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 5534 16232 5540 16244
rect 5495 16204 5540 16232
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 8628 16204 8769 16232
rect 8628 16192 8634 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 9490 16232 9496 16244
rect 9451 16204 9496 16232
rect 8757 16195 8815 16201
rect 1762 16124 1768 16176
rect 1820 16164 1826 16176
rect 2133 16167 2191 16173
rect 2133 16164 2145 16167
rect 1820 16136 2145 16164
rect 1820 16124 1826 16136
rect 2133 16133 2145 16136
rect 2179 16164 2191 16167
rect 2958 16164 2964 16176
rect 2179 16136 2964 16164
rect 2179 16133 2191 16136
rect 2133 16127 2191 16133
rect 2958 16124 2964 16136
rect 3016 16164 3022 16176
rect 3016 16136 3280 16164
rect 3016 16124 3022 16136
rect 3252 16105 3280 16136
rect 5442 16124 5448 16176
rect 5500 16164 5506 16176
rect 5813 16167 5871 16173
rect 5813 16164 5825 16167
rect 5500 16136 5825 16164
rect 5500 16124 5506 16136
rect 5813 16133 5825 16136
rect 5859 16133 5871 16167
rect 5813 16127 5871 16133
rect 8481 16167 8539 16173
rect 8481 16133 8493 16167
rect 8527 16164 8539 16167
rect 8662 16164 8668 16176
rect 8527 16136 8668 16164
rect 8527 16133 8539 16136
rect 8481 16127 8539 16133
rect 8662 16124 8668 16136
rect 8720 16124 8726 16176
rect 3237 16099 3295 16105
rect 3237 16065 3249 16099
rect 3283 16065 3295 16099
rect 8772 16096 8800 16195
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10873 16235 10931 16241
rect 10873 16232 10885 16235
rect 10376 16204 10885 16232
rect 10376 16192 10382 16204
rect 10873 16201 10885 16204
rect 10919 16201 10931 16235
rect 10873 16195 10931 16201
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16232 11391 16235
rect 11606 16232 11612 16244
rect 11379 16204 11612 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 15010 16232 15016 16244
rect 14971 16204 15016 16232
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 20622 16232 20628 16244
rect 19484 16204 20628 16232
rect 19484 16192 19490 16204
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 21358 16192 21364 16244
rect 21416 16232 21422 16244
rect 21453 16235 21511 16241
rect 21453 16232 21465 16235
rect 21416 16204 21465 16232
rect 21416 16192 21422 16204
rect 21453 16201 21465 16204
rect 21499 16201 21511 16235
rect 23474 16232 23480 16244
rect 23435 16204 23480 16232
rect 21453 16195 21511 16201
rect 23474 16192 23480 16204
rect 23532 16192 23538 16244
rect 24946 16124 24952 16176
rect 25004 16164 25010 16176
rect 25590 16164 25596 16176
rect 25004 16136 25596 16164
rect 25004 16124 25010 16136
rect 25590 16124 25596 16136
rect 25648 16124 25654 16176
rect 10045 16099 10103 16105
rect 10045 16096 10057 16099
rect 8772 16068 10057 16096
rect 3237 16059 3295 16065
rect 10045 16065 10057 16068
rect 10091 16096 10103 16099
rect 10502 16096 10508 16108
rect 10091 16068 10508 16096
rect 10091 16065 10103 16068
rect 10045 16059 10103 16065
rect 10502 16056 10508 16068
rect 10560 16096 10566 16108
rect 11974 16096 11980 16108
rect 10560 16068 11980 16096
rect 10560 16056 10566 16068
rect 11974 16056 11980 16068
rect 12032 16056 12038 16108
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13412 16068 13737 16096
rect 13412 16056 13418 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 13817 16099 13875 16105
rect 13817 16065 13829 16099
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 3142 15988 3148 16040
rect 3200 16028 3206 16040
rect 4982 16028 4988 16040
rect 3200 16000 4988 16028
rect 3200 15988 3206 16000
rect 4982 15988 4988 16000
rect 5040 16028 5046 16040
rect 10870 16028 10876 16040
rect 5040 16000 10876 16028
rect 5040 15988 5046 16000
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 16028 13231 16031
rect 13538 16028 13544 16040
rect 13219 16000 13544 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 13538 15988 13544 16000
rect 13596 16028 13602 16040
rect 13832 16028 13860 16059
rect 21542 16056 21548 16108
rect 21600 16096 21606 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21600 16068 22017 16096
rect 21600 16056 21606 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 23937 16099 23995 16105
rect 23937 16065 23949 16099
rect 23983 16096 23995 16099
rect 24210 16096 24216 16108
rect 23983 16068 24216 16096
rect 23983 16065 23995 16068
rect 23937 16059 23995 16065
rect 24210 16056 24216 16068
rect 24268 16096 24274 16108
rect 24670 16096 24676 16108
rect 24268 16068 24676 16096
rect 24268 16056 24274 16068
rect 24670 16056 24676 16068
rect 24728 16056 24734 16108
rect 25133 16099 25191 16105
rect 25133 16065 25145 16099
rect 25179 16096 25191 16099
rect 26237 16099 26295 16105
rect 26237 16096 26249 16099
rect 25179 16068 26249 16096
rect 25179 16065 25191 16068
rect 25133 16059 25191 16065
rect 26237 16065 26249 16068
rect 26283 16096 26295 16099
rect 26326 16096 26332 16108
rect 26283 16068 26332 16096
rect 26283 16065 26295 16068
rect 26237 16059 26295 16065
rect 26326 16056 26332 16068
rect 26384 16096 26390 16108
rect 27154 16096 27160 16108
rect 26384 16068 27160 16096
rect 26384 16056 26390 16068
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 13596 16000 13860 16028
rect 15749 16031 15807 16037
rect 13596 15988 13602 16000
rect 15749 15997 15761 16031
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 2593 15963 2651 15969
rect 2593 15929 2605 15963
rect 2639 15960 2651 15963
rect 2866 15960 2872 15972
rect 2639 15932 2872 15960
rect 2639 15929 2651 15932
rect 2593 15923 2651 15929
rect 2866 15920 2872 15932
rect 2924 15960 2930 15972
rect 3053 15963 3111 15969
rect 3053 15960 3065 15963
rect 2924 15932 3065 15960
rect 2924 15920 2930 15932
rect 3053 15929 3065 15932
rect 3099 15960 3111 15963
rect 3510 15960 3516 15972
rect 3099 15932 3516 15960
rect 3099 15929 3111 15932
rect 3053 15923 3111 15929
rect 3510 15920 3516 15932
rect 3568 15920 3574 15972
rect 12805 15963 12863 15969
rect 12805 15929 12817 15963
rect 12851 15960 12863 15963
rect 13633 15963 13691 15969
rect 13633 15960 13645 15963
rect 12851 15932 13645 15960
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 13633 15929 13645 15932
rect 13679 15960 13691 15963
rect 13722 15960 13728 15972
rect 13679 15932 13728 15960
rect 13679 15929 13691 15932
rect 13633 15923 13691 15929
rect 13722 15920 13728 15932
rect 13780 15920 13786 15972
rect 15764 15960 15792 15991
rect 15838 15988 15844 16040
rect 15896 16028 15902 16040
rect 16005 16031 16063 16037
rect 16005 16028 16017 16031
rect 15896 16000 16017 16028
rect 15896 15988 15902 16000
rect 16005 15997 16017 16000
rect 16051 15997 16063 16031
rect 16005 15991 16063 15997
rect 19245 16031 19303 16037
rect 19245 15997 19257 16031
rect 19291 16028 19303 16031
rect 19334 16028 19340 16040
rect 19291 16000 19340 16028
rect 19291 15997 19303 16000
rect 19245 15991 19303 15997
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 24397 16031 24455 16037
rect 24397 15997 24409 16031
rect 24443 16028 24455 16031
rect 24762 16028 24768 16040
rect 24443 16000 24768 16028
rect 24443 15997 24455 16000
rect 24397 15991 24455 15997
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 25961 16031 26019 16037
rect 25961 16028 25973 16031
rect 25424 16000 25973 16028
rect 16298 15960 16304 15972
rect 15764 15932 16304 15960
rect 16298 15920 16304 15932
rect 16356 15920 16362 15972
rect 17494 15960 17500 15972
rect 16408 15932 17500 15960
rect 3145 15895 3203 15901
rect 3145 15861 3157 15895
rect 3191 15892 3203 15895
rect 3602 15892 3608 15904
rect 3191 15864 3608 15892
rect 3191 15861 3203 15864
rect 3145 15855 3203 15861
rect 3602 15852 3608 15864
rect 3660 15892 3666 15904
rect 3697 15895 3755 15901
rect 3697 15892 3709 15895
rect 3660 15864 3709 15892
rect 3660 15852 3666 15864
rect 3697 15861 3709 15864
rect 3743 15861 3755 15895
rect 8110 15892 8116 15904
rect 8071 15864 8116 15892
rect 3697 15855 3755 15861
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 9401 15895 9459 15901
rect 9401 15892 9413 15895
rect 8352 15864 9413 15892
rect 8352 15852 8358 15864
rect 9401 15861 9413 15864
rect 9447 15892 9459 15895
rect 9861 15895 9919 15901
rect 9861 15892 9873 15895
rect 9447 15864 9873 15892
rect 9447 15861 9459 15864
rect 9401 15855 9459 15861
rect 9861 15861 9873 15864
rect 9907 15861 9919 15895
rect 9861 15855 9919 15861
rect 9950 15852 9956 15904
rect 10008 15892 10014 15904
rect 11698 15892 11704 15904
rect 10008 15864 10053 15892
rect 11659 15864 11704 15892
rect 10008 15852 10014 15864
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 13262 15892 13268 15904
rect 13223 15864 13268 15892
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 15381 15895 15439 15901
rect 15381 15861 15393 15895
rect 15427 15892 15439 15895
rect 15654 15892 15660 15904
rect 15427 15864 15660 15892
rect 15427 15861 15439 15864
rect 15381 15855 15439 15861
rect 15654 15852 15660 15864
rect 15712 15892 15718 15904
rect 16408 15892 16436 15932
rect 17494 15920 17500 15932
rect 17552 15920 17558 15972
rect 19153 15963 19211 15969
rect 19153 15929 19165 15963
rect 19199 15960 19211 15963
rect 19490 15963 19548 15969
rect 19490 15960 19502 15963
rect 19199 15932 19502 15960
rect 19199 15929 19211 15932
rect 19153 15923 19211 15929
rect 19490 15929 19502 15932
rect 19536 15960 19548 15963
rect 20714 15960 20720 15972
rect 19536 15932 20720 15960
rect 19536 15929 19548 15932
rect 19490 15923 19548 15929
rect 20714 15920 20720 15932
rect 20772 15920 20778 15972
rect 21818 15960 21824 15972
rect 21779 15932 21824 15960
rect 21818 15920 21824 15932
rect 21876 15920 21882 15972
rect 17126 15892 17132 15904
rect 15712 15864 16436 15892
rect 17087 15864 17132 15892
rect 15712 15852 15718 15864
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 21269 15895 21327 15901
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21358 15892 21364 15904
rect 21315 15864 21364 15892
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 21910 15892 21916 15904
rect 21871 15864 21916 15892
rect 21910 15852 21916 15864
rect 21968 15892 21974 15904
rect 22465 15895 22523 15901
rect 22465 15892 22477 15895
rect 21968 15864 22477 15892
rect 21968 15852 21974 15864
rect 22465 15861 22477 15864
rect 22511 15861 22523 15895
rect 22830 15892 22836 15904
rect 22791 15864 22836 15892
rect 22465 15855 22523 15861
rect 22830 15852 22836 15864
rect 22888 15852 22894 15904
rect 24026 15892 24032 15904
rect 23987 15864 24032 15892
rect 24026 15852 24032 15864
rect 24084 15852 24090 15904
rect 24486 15852 24492 15904
rect 24544 15892 24550 15904
rect 24544 15864 24589 15892
rect 24544 15852 24550 15864
rect 25130 15852 25136 15904
rect 25188 15892 25194 15904
rect 25424 15901 25452 16000
rect 25961 15997 25973 16000
rect 26007 15997 26019 16031
rect 25961 15991 26019 15997
rect 25866 15920 25872 15972
rect 25924 15960 25930 15972
rect 25924 15932 26096 15960
rect 25924 15920 25930 15932
rect 25409 15895 25467 15901
rect 25409 15892 25421 15895
rect 25188 15864 25421 15892
rect 25188 15852 25194 15864
rect 25409 15861 25421 15864
rect 25455 15861 25467 15895
rect 25590 15892 25596 15904
rect 25551 15864 25596 15892
rect 25409 15855 25467 15861
rect 25590 15852 25596 15864
rect 25648 15852 25654 15904
rect 26068 15901 26096 15932
rect 26053 15895 26111 15901
rect 26053 15861 26065 15895
rect 26099 15892 26111 15895
rect 26605 15895 26663 15901
rect 26605 15892 26617 15895
rect 26099 15864 26617 15892
rect 26099 15861 26111 15864
rect 26053 15855 26111 15861
rect 26605 15861 26617 15864
rect 26651 15861 26663 15895
rect 26605 15855 26663 15861
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 2406 15688 2412 15700
rect 2367 15660 2412 15688
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 9122 15688 9128 15700
rect 9083 15660 9128 15688
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 9950 15688 9956 15700
rect 9539 15660 9956 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10502 15648 10508 15700
rect 10560 15688 10566 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 10560 15660 11069 15688
rect 10560 15648 10566 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 13354 15688 13360 15700
rect 13315 15660 13360 15688
rect 11057 15651 11115 15657
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 15838 15688 15844 15700
rect 15799 15660 15844 15688
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 19334 15688 19340 15700
rect 19295 15660 19340 15688
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 20622 15648 20628 15700
rect 20680 15688 20686 15700
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 20680 15660 21189 15688
rect 20680 15648 20686 15660
rect 21177 15657 21189 15660
rect 21223 15688 21235 15691
rect 21542 15688 21548 15700
rect 21223 15660 21548 15688
rect 21223 15657 21235 15660
rect 21177 15651 21235 15657
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 21634 15648 21640 15700
rect 21692 15688 21698 15700
rect 21729 15691 21787 15697
rect 21729 15688 21741 15691
rect 21692 15660 21741 15688
rect 21692 15648 21698 15660
rect 21729 15657 21741 15660
rect 21775 15688 21787 15691
rect 22830 15688 22836 15700
rect 21775 15660 22836 15688
rect 21775 15657 21787 15660
rect 21729 15651 21787 15657
rect 22830 15648 22836 15660
rect 22888 15648 22894 15700
rect 24121 15691 24179 15697
rect 24121 15657 24133 15691
rect 24167 15688 24179 15691
rect 24486 15688 24492 15700
rect 24167 15660 24492 15688
rect 24167 15657 24179 15660
rect 24121 15651 24179 15657
rect 24486 15648 24492 15660
rect 24544 15688 24550 15700
rect 24857 15691 24915 15697
rect 24857 15688 24869 15691
rect 24544 15660 24869 15688
rect 24544 15648 24550 15660
rect 24857 15657 24869 15660
rect 24903 15657 24915 15691
rect 24857 15651 24915 15657
rect 25317 15691 25375 15697
rect 25317 15657 25329 15691
rect 25363 15688 25375 15691
rect 25590 15688 25596 15700
rect 25363 15660 25596 15688
rect 25363 15657 25375 15660
rect 25317 15651 25375 15657
rect 25590 15648 25596 15660
rect 25648 15648 25654 15700
rect 26513 15691 26571 15697
rect 26513 15657 26525 15691
rect 26559 15657 26571 15691
rect 26513 15651 26571 15657
rect 2774 15580 2780 15632
rect 2832 15620 2838 15632
rect 4062 15620 4068 15632
rect 2832 15592 4068 15620
rect 2832 15580 2838 15592
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 5261 15623 5319 15629
rect 5261 15589 5273 15623
rect 5307 15620 5319 15623
rect 6270 15620 6276 15632
rect 5307 15592 6276 15620
rect 5307 15589 5319 15592
rect 5261 15583 5319 15589
rect 6270 15580 6276 15592
rect 6328 15620 6334 15632
rect 6448 15623 6506 15629
rect 6448 15620 6460 15623
rect 6328 15592 6460 15620
rect 6328 15580 6334 15592
rect 6448 15589 6460 15592
rect 6494 15620 6506 15623
rect 6822 15620 6828 15632
rect 6494 15592 6828 15620
rect 6494 15589 6506 15592
rect 6448 15583 6506 15589
rect 6822 15580 6828 15592
rect 6880 15580 6886 15632
rect 17126 15580 17132 15632
rect 17184 15620 17190 15632
rect 17374 15623 17432 15629
rect 17374 15620 17386 15623
rect 17184 15592 17386 15620
rect 17184 15580 17190 15592
rect 17374 15589 17386 15592
rect 17420 15589 17432 15623
rect 17374 15583 17432 15589
rect 24670 15580 24676 15632
rect 24728 15620 24734 15632
rect 25225 15623 25283 15629
rect 25225 15620 25237 15623
rect 24728 15592 25237 15620
rect 24728 15580 24734 15592
rect 25225 15589 25237 15592
rect 25271 15620 25283 15623
rect 26528 15620 26556 15651
rect 25271 15592 26556 15620
rect 26881 15623 26939 15629
rect 25271 15589 25283 15592
rect 25225 15583 25283 15589
rect 26881 15589 26893 15623
rect 26927 15620 26939 15623
rect 27062 15620 27068 15632
rect 26927 15592 27068 15620
rect 26927 15589 26939 15592
rect 26881 15583 26939 15589
rect 27062 15580 27068 15592
rect 27120 15580 27126 15632
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15552 2375 15555
rect 2406 15552 2412 15564
rect 2363 15524 2412 15552
rect 2363 15521 2375 15524
rect 2317 15515 2375 15521
rect 2406 15512 2412 15524
rect 2464 15552 2470 15564
rect 2869 15555 2927 15561
rect 2869 15552 2881 15555
rect 2464 15524 2881 15552
rect 2464 15512 2470 15524
rect 2869 15521 2881 15524
rect 2915 15521 2927 15555
rect 2869 15515 2927 15521
rect 5442 15512 5448 15564
rect 5500 15552 5506 15564
rect 6181 15555 6239 15561
rect 6181 15552 6193 15555
rect 5500 15524 6193 15552
rect 5500 15512 5506 15524
rect 6181 15521 6193 15524
rect 6227 15521 6239 15555
rect 6181 15515 6239 15521
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 9933 15555 9991 15561
rect 9933 15552 9945 15555
rect 9824 15524 9945 15552
rect 9824 15512 9830 15524
rect 9933 15521 9945 15524
rect 9979 15521 9991 15555
rect 13722 15552 13728 15564
rect 13683 15524 13728 15552
rect 9933 15515 9991 15521
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 19334 15552 19340 15564
rect 17144 15524 19340 15552
rect 2958 15484 2964 15496
rect 2919 15456 2964 15484
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 9732 15456 9777 15484
rect 9732 15444 9738 15456
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 13817 15487 13875 15493
rect 13817 15484 13829 15487
rect 13044 15456 13829 15484
rect 13044 15444 13050 15456
rect 13817 15453 13829 15456
rect 13863 15453 13875 15487
rect 13817 15447 13875 15453
rect 14001 15487 14059 15493
rect 14001 15453 14013 15487
rect 14047 15484 14059 15487
rect 15838 15484 15844 15496
rect 14047 15456 15844 15484
rect 14047 15453 14059 15456
rect 14001 15447 14059 15453
rect 12894 15376 12900 15428
rect 12952 15416 12958 15428
rect 14016 15416 14044 15447
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16298 15484 16304 15496
rect 16211 15456 16304 15484
rect 16298 15444 16304 15456
rect 16356 15484 16362 15496
rect 16758 15484 16764 15496
rect 16356 15456 16764 15484
rect 16356 15444 16362 15456
rect 16758 15444 16764 15456
rect 16816 15484 16822 15496
rect 17144 15493 17172 15524
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 22097 15555 22155 15561
rect 22097 15521 22109 15555
rect 22143 15552 22155 15555
rect 22646 15552 22652 15564
rect 22143 15524 22652 15552
rect 22143 15521 22155 15524
rect 22097 15515 22155 15521
rect 22646 15512 22652 15524
rect 22704 15512 22710 15564
rect 24489 15555 24547 15561
rect 24489 15521 24501 15555
rect 24535 15552 24547 15555
rect 24762 15552 24768 15564
rect 24535 15524 24768 15552
rect 24535 15521 24547 15524
rect 24489 15515 24547 15521
rect 24762 15512 24768 15524
rect 24820 15512 24826 15564
rect 26973 15555 27031 15561
rect 26973 15521 26985 15555
rect 27019 15552 27031 15555
rect 27246 15552 27252 15564
rect 27019 15524 27252 15552
rect 27019 15521 27031 15524
rect 26973 15515 27031 15521
rect 27246 15512 27252 15524
rect 27304 15512 27310 15564
rect 17129 15487 17187 15493
rect 17129 15484 17141 15487
rect 16816 15456 17141 15484
rect 16816 15444 16822 15456
rect 17129 15453 17141 15456
rect 17175 15453 17187 15487
rect 17129 15447 17187 15453
rect 21174 15444 21180 15496
rect 21232 15484 21238 15496
rect 22189 15487 22247 15493
rect 22189 15484 22201 15487
rect 21232 15456 22201 15484
rect 21232 15444 21238 15456
rect 22189 15453 22201 15456
rect 22235 15453 22247 15487
rect 22189 15447 22247 15453
rect 22278 15444 22284 15496
rect 22336 15484 22342 15496
rect 25406 15484 25412 15496
rect 22336 15456 22381 15484
rect 25367 15456 25412 15484
rect 22336 15444 22342 15456
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 27154 15484 27160 15496
rect 27115 15456 27160 15484
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 12952 15388 14044 15416
rect 12952 15376 12958 15388
rect 1670 15348 1676 15360
rect 1631 15320 1676 15348
rect 1670 15308 1676 15320
rect 1728 15348 1734 15360
rect 3694 15348 3700 15360
rect 1728 15320 3700 15348
rect 1728 15308 1734 15320
rect 3694 15308 3700 15320
rect 3752 15308 3758 15360
rect 7558 15348 7564 15360
rect 7519 15320 7564 15348
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15473 15351 15531 15357
rect 15473 15348 15485 15351
rect 15252 15320 15485 15348
rect 15252 15308 15258 15320
rect 15473 15317 15485 15320
rect 15519 15317 15531 15351
rect 18506 15348 18512 15360
rect 18467 15320 18512 15348
rect 15473 15311 15531 15317
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 23566 15348 23572 15360
rect 23479 15320 23572 15348
rect 23566 15308 23572 15320
rect 23624 15348 23630 15360
rect 24302 15348 24308 15360
rect 23624 15320 24308 15348
rect 23624 15308 23630 15320
rect 24302 15308 24308 15320
rect 24360 15308 24366 15360
rect 25038 15308 25044 15360
rect 25096 15348 25102 15360
rect 25961 15351 26019 15357
rect 25961 15348 25973 15351
rect 25096 15320 25973 15348
rect 25096 15308 25102 15320
rect 25961 15317 25973 15320
rect 26007 15348 26019 15351
rect 26326 15348 26332 15360
rect 26007 15320 26332 15348
rect 26007 15317 26019 15320
rect 25961 15311 26019 15317
rect 26326 15308 26332 15320
rect 26384 15308 26390 15360
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 2958 15144 2964 15156
rect 2823 15116 2964 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 2958 15104 2964 15116
rect 3016 15144 3022 15156
rect 3053 15147 3111 15153
rect 3053 15144 3065 15147
rect 3016 15116 3065 15144
rect 3016 15104 3022 15116
rect 3053 15113 3065 15116
rect 3099 15113 3111 15147
rect 3602 15144 3608 15156
rect 3563 15116 3608 15144
rect 3053 15107 3111 15113
rect 3602 15104 3608 15116
rect 3660 15104 3666 15156
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 4617 15147 4675 15153
rect 4617 15144 4629 15147
rect 4120 15116 4629 15144
rect 4120 15104 4126 15116
rect 4617 15113 4629 15116
rect 4663 15113 4675 15147
rect 6270 15144 6276 15156
rect 6231 15116 6276 15144
rect 4617 15107 4675 15113
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 6365 15147 6423 15153
rect 6365 15113 6377 15147
rect 6411 15144 6423 15147
rect 9125 15147 9183 15153
rect 9125 15144 9137 15147
rect 6411 15116 9137 15144
rect 6411 15113 6423 15116
rect 6365 15107 6423 15113
rect 9125 15113 9137 15116
rect 9171 15113 9183 15147
rect 9125 15107 9183 15113
rect 9582 15104 9588 15156
rect 9640 15104 9646 15156
rect 9766 15144 9772 15156
rect 9727 15116 9772 15144
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 12894 15144 12900 15156
rect 12855 15116 12900 15144
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 16758 15144 16764 15156
rect 13556 15116 16344 15144
rect 16719 15116 16764 15144
rect 6638 15076 6644 15088
rect 5644 15048 6644 15076
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 3694 14968 3700 15020
rect 3752 15008 3758 15020
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 3752 14980 4169 15008
rect 3752 14968 3758 14980
rect 4157 14977 4169 14980
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 4614 14968 4620 15020
rect 4672 15008 4678 15020
rect 5644 15017 5672 15048
rect 6638 15036 6644 15048
rect 6696 15076 6702 15088
rect 6696 15048 7512 15076
rect 6696 15036 6702 15048
rect 5077 15011 5135 15017
rect 5077 15008 5089 15011
rect 4672 14980 5089 15008
rect 4672 14968 4678 14980
rect 5077 14977 5089 14980
rect 5123 15008 5135 15011
rect 5629 15011 5687 15017
rect 5629 15008 5641 15011
rect 5123 14980 5641 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5629 14977 5641 14980
rect 5675 14977 5687 15011
rect 5629 14971 5687 14977
rect 5813 15011 5871 15017
rect 5813 14977 5825 15011
rect 5859 15008 5871 15011
rect 6270 15008 6276 15020
rect 5859 14980 6276 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 6270 14968 6276 14980
rect 6328 15008 6334 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 6328 14980 7389 15008
rect 6328 14968 6334 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 7484 15008 7512 15048
rect 9306 15036 9312 15088
rect 9364 15076 9370 15088
rect 9600 15076 9628 15104
rect 9364 15048 9628 15076
rect 9364 15036 9370 15048
rect 9858 15036 9864 15088
rect 9916 15076 9922 15088
rect 13556 15076 13584 15116
rect 13722 15076 13728 15088
rect 9916 15048 13584 15076
rect 13635 15048 13728 15076
rect 9916 15036 9922 15048
rect 13722 15036 13728 15048
rect 13780 15076 13786 15088
rect 15197 15079 15255 15085
rect 15197 15076 15209 15079
rect 13780 15048 15209 15076
rect 13780 15036 13786 15048
rect 15197 15045 15209 15048
rect 15243 15045 15255 15079
rect 16316 15076 16344 15116
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 17126 15144 17132 15156
rect 17087 15116 17132 15144
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 19886 15104 19892 15156
rect 19944 15144 19950 15156
rect 21174 15144 21180 15156
rect 19944 15116 21180 15144
rect 19944 15104 19950 15116
rect 21174 15104 21180 15116
rect 21232 15104 21238 15156
rect 21637 15147 21695 15153
rect 21637 15113 21649 15147
rect 21683 15144 21695 15147
rect 21910 15144 21916 15156
rect 21683 15116 21916 15144
rect 21683 15113 21695 15116
rect 21637 15107 21695 15113
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 22738 15144 22744 15156
rect 22699 15116 22744 15144
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 24581 15147 24639 15153
rect 24581 15113 24593 15147
rect 24627 15144 24639 15147
rect 24670 15144 24676 15156
rect 24627 15116 24676 15144
rect 24627 15113 24639 15116
rect 24581 15107 24639 15113
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 25317 15147 25375 15153
rect 25317 15113 25329 15147
rect 25363 15144 25375 15147
rect 25590 15144 25596 15156
rect 25363 15116 25596 15144
rect 25363 15113 25375 15116
rect 25317 15107 25375 15113
rect 25590 15104 25596 15116
rect 25648 15104 25654 15156
rect 25866 15144 25872 15156
rect 25827 15116 25872 15144
rect 25866 15104 25872 15116
rect 25924 15104 25930 15156
rect 17681 15079 17739 15085
rect 17681 15076 17693 15079
rect 16316 15048 17693 15076
rect 15197 15039 15255 15045
rect 17681 15045 17693 15048
rect 17727 15076 17739 15079
rect 17773 15079 17831 15085
rect 17773 15076 17785 15079
rect 17727 15048 17785 15076
rect 17727 15045 17739 15048
rect 17681 15039 17739 15045
rect 17773 15045 17785 15048
rect 17819 15045 17831 15079
rect 17773 15039 17831 15045
rect 24949 15079 25007 15085
rect 24949 15045 24961 15079
rect 24995 15076 25007 15079
rect 25406 15076 25412 15088
rect 24995 15048 25412 15076
rect 24995 15045 25007 15048
rect 24949 15039 25007 15045
rect 25406 15036 25412 15048
rect 25464 15036 25470 15088
rect 10226 15008 10232 15020
rect 7484 14980 10232 15008
rect 7377 14971 7435 14977
rect 10226 14968 10232 14980
rect 10284 14968 10290 15020
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 11333 15011 11391 15017
rect 11333 15008 11345 15011
rect 10367 14980 11345 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 11333 14977 11345 14980
rect 11379 15008 11391 15011
rect 12158 15008 12164 15020
rect 11379 14980 12164 15008
rect 11379 14977 11391 14980
rect 11333 14971 11391 14977
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 14182 14968 14188 15020
rect 14240 15008 14246 15020
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 14240 14980 14289 15008
rect 14240 14968 14246 14980
rect 14277 14977 14289 14980
rect 14323 15008 14335 15011
rect 15102 15008 15108 15020
rect 14323 14980 15108 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 18506 14968 18512 15020
rect 18564 15008 18570 15020
rect 18601 15011 18659 15017
rect 18601 15008 18613 15011
rect 18564 14980 18613 15008
rect 18564 14968 18570 14980
rect 18601 14977 18613 14980
rect 18647 15008 18659 15011
rect 19058 15008 19064 15020
rect 18647 14980 19064 15008
rect 18647 14977 18659 14980
rect 18601 14971 18659 14977
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21266 15008 21272 15020
rect 20772 14980 21272 15008
rect 20772 14968 20778 14980
rect 21266 14968 21272 14980
rect 21324 15008 21330 15020
rect 22278 15008 22284 15020
rect 21324 14980 22284 15008
rect 21324 14968 21330 14980
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 26326 14968 26332 15020
rect 26384 15008 26390 15020
rect 26421 15011 26479 15017
rect 26421 15008 26433 15011
rect 26384 14980 26433 15008
rect 26384 14968 26390 14980
rect 26421 14977 26433 14980
rect 26467 14977 26479 15011
rect 26421 14971 26479 14977
rect 1670 14949 1676 14952
rect 1664 14940 1676 14949
rect 1631 14912 1676 14940
rect 1664 14903 1676 14912
rect 1670 14900 1676 14903
rect 1728 14900 1734 14952
rect 5442 14900 5448 14952
rect 5500 14940 5506 14952
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 5500 14912 7849 14940
rect 5500 14900 5506 14912
rect 7837 14909 7849 14912
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14940 9183 14943
rect 9398 14940 9404 14952
rect 9171 14912 9404 14940
rect 9171 14909 9183 14912
rect 9125 14903 9183 14909
rect 9398 14900 9404 14912
rect 9456 14900 9462 14952
rect 10870 14900 10876 14952
rect 10928 14940 10934 14952
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 10928 14912 13645 14940
rect 10928 14900 10934 14912
rect 13633 14909 13645 14912
rect 13679 14940 13691 14943
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 13679 14912 14105 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 14093 14909 14105 14912
rect 14139 14940 14151 14943
rect 14550 14940 14556 14952
rect 14139 14912 14556 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 18414 14940 18420 14952
rect 17420 14912 18420 14940
rect 1118 14832 1124 14884
rect 1176 14872 1182 14884
rect 3513 14875 3571 14881
rect 3513 14872 3525 14875
rect 1176 14844 3525 14872
rect 1176 14832 1182 14844
rect 3513 14841 3525 14844
rect 3559 14872 3571 14875
rect 4065 14875 4123 14881
rect 4065 14872 4077 14875
rect 3559 14844 4077 14872
rect 3559 14841 3571 14844
rect 3513 14835 3571 14841
rect 4065 14841 4077 14844
rect 4111 14872 4123 14875
rect 6365 14875 6423 14881
rect 6365 14872 6377 14875
rect 4111 14844 6377 14872
rect 4111 14841 4123 14844
rect 4065 14835 4123 14841
rect 6365 14841 6377 14844
rect 6411 14841 6423 14875
rect 6365 14835 6423 14841
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 7006 14872 7012 14884
rect 6687 14844 7012 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7006 14832 7012 14844
rect 7064 14872 7070 14884
rect 7285 14875 7343 14881
rect 7285 14872 7297 14875
rect 7064 14844 7297 14872
rect 7064 14832 7070 14844
rect 7285 14841 7297 14844
rect 7331 14872 7343 14875
rect 10597 14875 10655 14881
rect 10597 14872 10609 14875
rect 7331 14844 10609 14872
rect 7331 14841 7343 14844
rect 7285 14835 7343 14841
rect 10597 14841 10609 14844
rect 10643 14872 10655 14875
rect 11241 14875 11299 14881
rect 11241 14872 11253 14875
rect 10643 14844 11253 14872
rect 10643 14841 10655 14844
rect 10597 14835 10655 14841
rect 11241 14841 11253 14844
rect 11287 14841 11299 14875
rect 11241 14835 11299 14841
rect 12986 14832 12992 14884
rect 13044 14872 13050 14884
rect 14737 14875 14795 14881
rect 14737 14872 14749 14875
rect 13044 14844 14749 14872
rect 13044 14832 13050 14844
rect 14737 14841 14749 14844
rect 14783 14841 14795 14875
rect 14737 14835 14795 14841
rect 17420 14816 17448 14912
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 21726 14940 21732 14952
rect 20732 14912 21732 14940
rect 17681 14875 17739 14881
rect 17681 14841 17693 14875
rect 17727 14872 17739 14875
rect 18506 14872 18512 14884
rect 17727 14844 18512 14872
rect 17727 14841 17739 14844
rect 17681 14835 17739 14841
rect 18506 14832 18512 14844
rect 18564 14832 18570 14884
rect 20732 14816 20760 14912
rect 21726 14900 21732 14912
rect 21784 14940 21790 14952
rect 22005 14943 22063 14949
rect 22005 14940 22017 14943
rect 21784 14912 22017 14940
rect 21784 14900 21790 14912
rect 22005 14909 22017 14912
rect 22051 14909 22063 14943
rect 22005 14903 22063 14909
rect 21545 14875 21603 14881
rect 21545 14841 21557 14875
rect 21591 14872 21603 14875
rect 21910 14872 21916 14884
rect 21591 14844 21916 14872
rect 21591 14841 21603 14844
rect 21545 14835 21603 14841
rect 21910 14832 21916 14844
rect 21968 14872 21974 14884
rect 26329 14875 26387 14881
rect 26329 14872 26341 14875
rect 21968 14844 22048 14872
rect 21968 14832 21974 14844
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 3752 14776 3985 14804
rect 3752 14764 3758 14776
rect 3973 14773 3985 14776
rect 4019 14773 4031 14807
rect 5166 14804 5172 14816
rect 5127 14776 5172 14804
rect 3973 14767 4031 14773
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7190 14804 7196 14816
rect 7151 14776 7196 14804
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 9306 14804 9312 14816
rect 9267 14776 9312 14804
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 10778 14804 10784 14816
rect 10739 14776 10784 14804
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11149 14807 11207 14813
rect 11149 14773 11161 14807
rect 11195 14804 11207 14807
rect 11330 14804 11336 14816
rect 11195 14776 11336 14804
rect 11195 14773 11207 14776
rect 11149 14767 11207 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 13170 14764 13176 14816
rect 13228 14804 13234 14816
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 13228 14776 13277 14804
rect 13228 14764 13234 14776
rect 13265 14773 13277 14776
rect 13311 14804 13323 14807
rect 14182 14804 14188 14816
rect 13311 14776 14188 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 17402 14804 17408 14816
rect 17363 14776 17408 14804
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 18046 14804 18052 14816
rect 18007 14776 18052 14804
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 20714 14804 20720 14816
rect 20675 14776 20720 14804
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 22020 14804 22048 14844
rect 25700 14844 26341 14872
rect 25700 14816 25728 14844
rect 26329 14841 26341 14844
rect 26375 14841 26387 14875
rect 26329 14835 26387 14841
rect 22097 14807 22155 14813
rect 22097 14804 22109 14807
rect 22020 14776 22109 14804
rect 22097 14773 22109 14776
rect 22143 14773 22155 14807
rect 23106 14804 23112 14816
rect 23067 14776 23112 14804
rect 22097 14767 22155 14773
rect 23106 14764 23112 14776
rect 23164 14804 23170 14816
rect 23385 14807 23443 14813
rect 23385 14804 23397 14807
rect 23164 14776 23397 14804
rect 23164 14764 23170 14776
rect 23385 14773 23397 14776
rect 23431 14773 23443 14807
rect 25682 14804 25688 14816
rect 25643 14776 25688 14804
rect 23385 14767 23443 14773
rect 25682 14764 25688 14776
rect 25740 14764 25746 14816
rect 26237 14807 26295 14813
rect 26237 14773 26249 14807
rect 26283 14804 26295 14807
rect 26602 14804 26608 14816
rect 26283 14776 26608 14804
rect 26283 14773 26295 14776
rect 26237 14767 26295 14773
rect 26602 14764 26608 14776
rect 26660 14764 26666 14816
rect 26973 14807 27031 14813
rect 26973 14773 26985 14807
rect 27019 14804 27031 14807
rect 27062 14804 27068 14816
rect 27019 14776 27068 14804
rect 27019 14773 27031 14776
rect 26973 14767 27031 14773
rect 27062 14764 27068 14776
rect 27120 14764 27126 14816
rect 27246 14804 27252 14816
rect 27207 14776 27252 14804
rect 27246 14764 27252 14776
rect 27304 14764 27310 14816
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 2225 14603 2283 14609
rect 2225 14600 2237 14603
rect 1728 14572 2237 14600
rect 1728 14560 1734 14572
rect 2225 14569 2237 14572
rect 2271 14569 2283 14603
rect 2406 14600 2412 14612
rect 2367 14572 2412 14600
rect 2225 14563 2283 14569
rect 2240 14328 2268 14563
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 5166 14560 5172 14612
rect 5224 14600 5230 14612
rect 5813 14603 5871 14609
rect 5813 14600 5825 14603
rect 5224 14572 5825 14600
rect 5224 14560 5230 14572
rect 5813 14569 5825 14572
rect 5859 14600 5871 14603
rect 6546 14600 6552 14612
rect 5859 14572 6552 14600
rect 5859 14569 5871 14572
rect 5813 14563 5871 14569
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 6917 14603 6975 14609
rect 6917 14569 6929 14603
rect 6963 14600 6975 14603
rect 7190 14600 7196 14612
rect 6963 14572 7196 14600
rect 6963 14569 6975 14572
rect 6917 14563 6975 14569
rect 7190 14560 7196 14572
rect 7248 14560 7254 14612
rect 9677 14603 9735 14609
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 9950 14600 9956 14612
rect 9723 14572 9956 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10594 14560 10600 14612
rect 10652 14600 10658 14612
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 10652 14572 10885 14600
rect 10652 14560 10658 14572
rect 10873 14569 10885 14572
rect 10919 14600 10931 14603
rect 11330 14600 11336 14612
rect 10919 14572 11336 14600
rect 10919 14569 10931 14572
rect 10873 14563 10931 14569
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 12986 14600 12992 14612
rect 12947 14572 12992 14600
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16298 14600 16304 14612
rect 15804 14572 16304 14600
rect 15804 14560 15810 14572
rect 16298 14560 16304 14572
rect 16356 14600 16362 14612
rect 16669 14603 16727 14609
rect 16669 14600 16681 14603
rect 16356 14572 16681 14600
rect 16356 14560 16362 14572
rect 16669 14569 16681 14572
rect 16715 14569 16727 14603
rect 16669 14563 16727 14569
rect 16761 14603 16819 14609
rect 16761 14569 16773 14603
rect 16807 14600 16819 14603
rect 17126 14600 17132 14612
rect 16807 14572 17132 14600
rect 16807 14569 16819 14572
rect 16761 14563 16819 14569
rect 17126 14560 17132 14572
rect 17184 14600 17190 14612
rect 18046 14600 18052 14612
rect 17184 14572 18052 14600
rect 17184 14560 17190 14572
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 19334 14600 19340 14612
rect 19295 14572 19340 14600
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 21637 14603 21695 14609
rect 21637 14569 21649 14603
rect 21683 14600 21695 14603
rect 21818 14600 21824 14612
rect 21683 14572 21824 14600
rect 21683 14569 21695 14572
rect 21637 14563 21695 14569
rect 21818 14560 21824 14572
rect 21876 14560 21882 14612
rect 26789 14603 26847 14609
rect 26789 14569 26801 14603
rect 26835 14600 26847 14603
rect 27154 14600 27160 14612
rect 26835 14572 27160 14600
rect 26835 14569 26847 14572
rect 26789 14563 26847 14569
rect 27154 14560 27160 14572
rect 27212 14560 27218 14612
rect 2866 14532 2872 14544
rect 2827 14504 2872 14532
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 5905 14535 5963 14541
rect 5905 14532 5917 14535
rect 4764 14504 5917 14532
rect 4764 14492 4770 14504
rect 5905 14501 5917 14504
rect 5951 14532 5963 14535
rect 6822 14532 6828 14544
rect 5951 14504 6828 14532
rect 5951 14501 5963 14504
rect 5905 14495 5963 14501
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 13262 14492 13268 14544
rect 13320 14532 13326 14544
rect 13449 14535 13507 14541
rect 13449 14532 13461 14535
rect 13320 14504 13461 14532
rect 13320 14492 13326 14504
rect 13449 14501 13461 14504
rect 13495 14501 13507 14535
rect 13449 14495 13507 14501
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14464 2835 14467
rect 3602 14464 3608 14476
rect 2823 14436 3608 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 3602 14424 3608 14436
rect 3660 14424 3666 14476
rect 4341 14467 4399 14473
rect 4341 14433 4353 14467
rect 4387 14464 4399 14467
rect 5442 14464 5448 14476
rect 4387 14436 5448 14464
rect 4387 14433 4399 14436
rect 4341 14427 4399 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 6270 14424 6276 14476
rect 6328 14464 6334 14476
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 6328 14436 6469 14464
rect 6328 14424 6334 14436
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 9490 14464 9496 14476
rect 9451 14436 9496 14464
rect 6457 14427 6515 14433
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 12158 14424 12164 14476
rect 12216 14464 12222 14476
rect 13357 14467 13415 14473
rect 13357 14464 13369 14467
rect 12216 14436 13369 14464
rect 12216 14424 12222 14436
rect 13357 14433 13369 14436
rect 13403 14464 13415 14467
rect 13998 14464 14004 14476
rect 13403 14436 14004 14464
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 18230 14464 18236 14476
rect 18191 14436 18236 14464
rect 18230 14424 18236 14436
rect 18288 14424 18294 14476
rect 18690 14464 18696 14476
rect 18651 14436 18696 14464
rect 18690 14424 18696 14436
rect 18748 14424 18754 14476
rect 21818 14424 21824 14476
rect 21876 14464 21882 14476
rect 22005 14467 22063 14473
rect 22005 14464 22017 14467
rect 21876 14436 22017 14464
rect 21876 14424 21882 14436
rect 22005 14433 22017 14436
rect 22051 14433 22063 14467
rect 22005 14427 22063 14433
rect 2958 14396 2964 14408
rect 2919 14368 2964 14396
rect 2958 14356 2964 14368
rect 3016 14356 3022 14408
rect 3694 14396 3700 14408
rect 3655 14368 3700 14396
rect 3694 14356 3700 14368
rect 3752 14356 3758 14408
rect 5626 14356 5632 14408
rect 5684 14396 5690 14408
rect 5997 14399 6055 14405
rect 5997 14396 6009 14399
rect 5684 14368 6009 14396
rect 5684 14356 5690 14368
rect 5997 14365 6009 14368
rect 6043 14396 6055 14399
rect 7558 14396 7564 14408
rect 6043 14368 7564 14396
rect 6043 14365 6055 14368
rect 5997 14359 6055 14365
rect 7558 14356 7564 14368
rect 7616 14356 7622 14408
rect 10134 14396 10140 14408
rect 10095 14368 10140 14396
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14396 13691 14399
rect 16850 14396 16856 14408
rect 13679 14368 14136 14396
rect 16811 14368 16856 14396
rect 13679 14365 13691 14368
rect 13633 14359 13691 14365
rect 2976 14328 3004 14356
rect 2240 14300 3004 14328
rect 1394 14220 1400 14272
rect 1452 14260 1458 14272
rect 1673 14263 1731 14269
rect 1673 14260 1685 14263
rect 1452 14232 1685 14260
rect 1452 14220 1458 14232
rect 1673 14229 1685 14232
rect 1719 14260 1731 14263
rect 3712 14260 3740 14356
rect 5261 14331 5319 14337
rect 5261 14297 5273 14331
rect 5307 14328 5319 14331
rect 5534 14328 5540 14340
rect 5307 14300 5540 14328
rect 5307 14297 5319 14300
rect 5261 14291 5319 14297
rect 5534 14288 5540 14300
rect 5592 14328 5598 14340
rect 5810 14328 5816 14340
rect 5592 14300 5816 14328
rect 5592 14288 5598 14300
rect 5810 14288 5816 14300
rect 5868 14328 5874 14340
rect 6454 14328 6460 14340
rect 5868 14300 6460 14328
rect 5868 14288 5874 14300
rect 6454 14288 6460 14300
rect 6512 14288 6518 14340
rect 9766 14288 9772 14340
rect 9824 14328 9830 14340
rect 10244 14328 10272 14359
rect 10318 14328 10324 14340
rect 9824 14300 10324 14328
rect 9824 14288 9830 14300
rect 10318 14288 10324 14300
rect 10376 14288 10382 14340
rect 14108 14272 14136 14368
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 18782 14396 18788 14408
rect 18743 14368 18788 14396
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 18874 14356 18880 14408
rect 18932 14396 18938 14408
rect 22097 14399 22155 14405
rect 22097 14396 22109 14399
rect 18932 14368 18977 14396
rect 22020 14368 22109 14396
rect 18932 14356 18938 14368
rect 22020 14340 22048 14368
rect 22097 14365 22109 14368
rect 22143 14365 22155 14399
rect 22278 14396 22284 14408
rect 22191 14368 22284 14396
rect 22097 14359 22155 14365
rect 22278 14356 22284 14368
rect 22336 14396 22342 14408
rect 23106 14396 23112 14408
rect 22336 14368 23112 14396
rect 22336 14356 22342 14368
rect 23106 14356 23112 14368
rect 23164 14356 23170 14408
rect 18049 14331 18107 14337
rect 18049 14297 18061 14331
rect 18095 14328 18107 14331
rect 19150 14328 19156 14340
rect 18095 14300 19156 14328
rect 18095 14297 18107 14300
rect 18049 14291 18107 14297
rect 19150 14288 19156 14300
rect 19208 14328 19214 14340
rect 19334 14328 19340 14340
rect 19208 14300 19340 14328
rect 19208 14288 19214 14300
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 22002 14288 22008 14340
rect 22060 14288 22066 14340
rect 1719 14232 3740 14260
rect 4893 14263 4951 14269
rect 1719 14229 1731 14232
rect 1673 14223 1731 14229
rect 4893 14229 4905 14263
rect 4939 14260 4951 14263
rect 5074 14260 5080 14272
rect 4939 14232 5080 14260
rect 4939 14229 4951 14232
rect 4893 14223 4951 14229
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 5442 14260 5448 14272
rect 5403 14232 5448 14260
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 8110 14220 8116 14272
rect 8168 14260 8174 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8168 14232 8953 14260
rect 8168 14220 8174 14232
rect 8941 14229 8953 14232
rect 8987 14260 8999 14263
rect 9306 14260 9312 14272
rect 8987 14232 9312 14260
rect 8987 14229 8999 14232
rect 8941 14223 8999 14229
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 12526 14260 12532 14272
rect 12487 14232 12532 14260
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 14090 14260 14096 14272
rect 14051 14232 14096 14260
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 15565 14263 15623 14269
rect 15565 14229 15577 14263
rect 15611 14260 15623 14263
rect 15654 14260 15660 14272
rect 15611 14232 15660 14260
rect 15611 14229 15623 14232
rect 15565 14223 15623 14229
rect 15654 14220 15660 14232
rect 15712 14260 15718 14272
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 15712 14232 16313 14260
rect 15712 14220 15718 14232
rect 16301 14229 16313 14232
rect 16347 14229 16359 14263
rect 18322 14260 18328 14272
rect 18283 14232 18328 14260
rect 16301 14223 16359 14229
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 24302 14260 24308 14272
rect 24263 14232 24308 14260
rect 24302 14220 24308 14232
rect 24360 14220 24366 14272
rect 25961 14263 26019 14269
rect 25961 14229 25973 14263
rect 26007 14260 26019 14263
rect 26602 14260 26608 14272
rect 26007 14232 26608 14260
rect 26007 14229 26019 14232
rect 25961 14223 26019 14229
rect 26602 14220 26608 14232
rect 26660 14220 26666 14272
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 2406 14056 2412 14068
rect 1627 14028 2412 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 2682 14056 2688 14068
rect 2547 14028 2688 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 2682 14016 2688 14028
rect 2740 14016 2746 14068
rect 4706 14056 4712 14068
rect 4667 14028 4712 14056
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 6546 14056 6552 14068
rect 6507 14028 6552 14056
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 8846 14056 8852 14068
rect 8759 14028 8852 14056
rect 8846 14016 8852 14028
rect 8904 14056 8910 14068
rect 10042 14056 10048 14068
rect 8904 14028 10048 14056
rect 8904 14016 8910 14028
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10318 14056 10324 14068
rect 10279 14028 10324 14056
rect 10318 14016 10324 14028
rect 10376 14056 10382 14068
rect 10597 14059 10655 14065
rect 10597 14056 10609 14059
rect 10376 14028 10609 14056
rect 10376 14016 10382 14028
rect 10597 14025 10609 14028
rect 10643 14025 10655 14059
rect 14090 14056 14096 14068
rect 14051 14028 14096 14056
rect 10597 14019 10655 14025
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 16298 14056 16304 14068
rect 15120 14028 15884 14056
rect 16259 14028 16304 14056
rect 3602 13988 3608 14000
rect 3563 13960 3608 13988
rect 3602 13948 3608 13960
rect 3660 13948 3666 14000
rect 5077 13991 5135 13997
rect 5077 13957 5089 13991
rect 5123 13988 5135 13991
rect 5123 13960 5856 13988
rect 5123 13957 5135 13960
rect 5077 13951 5135 13957
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13920 2467 13923
rect 2866 13920 2872 13932
rect 2455 13892 2872 13920
rect 2455 13889 2467 13892
rect 2409 13883 2467 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 2958 13880 2964 13932
rect 3016 13920 3022 13932
rect 3145 13923 3203 13929
rect 3145 13920 3157 13923
rect 3016 13892 3157 13920
rect 3016 13880 3022 13892
rect 3145 13889 3157 13892
rect 3191 13920 3203 13923
rect 3881 13923 3939 13929
rect 3881 13920 3893 13923
rect 3191 13892 3893 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3881 13889 3893 13892
rect 3927 13889 3939 13923
rect 3881 13883 3939 13889
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 5442 13920 5448 13932
rect 4387 13892 5448 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 5442 13880 5448 13892
rect 5500 13920 5506 13932
rect 5828 13929 5856 13960
rect 10226 13948 10232 14000
rect 10284 13988 10290 14000
rect 12158 13988 12164 14000
rect 10284 13960 12164 13988
rect 10284 13948 10290 13960
rect 12158 13948 12164 13960
rect 12216 13948 12222 14000
rect 13814 13988 13820 14000
rect 13775 13960 13820 13988
rect 13814 13948 13820 13960
rect 13872 13988 13878 14000
rect 15120 13997 15148 14028
rect 15105 13991 15163 13997
rect 15105 13988 15117 13991
rect 13872 13960 15117 13988
rect 13872 13948 13878 13960
rect 15105 13957 15117 13960
rect 15151 13957 15163 13991
rect 15105 13951 15163 13957
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 15289 13991 15347 13997
rect 15289 13988 15301 13991
rect 15252 13960 15301 13988
rect 15252 13948 15258 13960
rect 15289 13957 15301 13960
rect 15335 13957 15347 13991
rect 15289 13951 15347 13957
rect 15856 13932 15884 14028
rect 16298 14016 16304 14028
rect 16356 14056 16362 14068
rect 16666 14056 16672 14068
rect 16356 14028 16672 14056
rect 16356 14016 16362 14028
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 17126 14056 17132 14068
rect 17087 14028 17132 14056
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 19058 14056 19064 14068
rect 19019 14028 19064 14056
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 19168 14028 20545 14056
rect 16850 13948 16856 14000
rect 16908 13988 16914 14000
rect 18325 13991 18383 13997
rect 18325 13988 18337 13991
rect 16908 13960 18337 13988
rect 16908 13948 16914 13960
rect 18325 13957 18337 13960
rect 18371 13988 18383 13991
rect 18874 13988 18880 14000
rect 18371 13960 18880 13988
rect 18371 13957 18383 13960
rect 18325 13951 18383 13957
rect 18874 13948 18880 13960
rect 18932 13988 18938 14000
rect 19168 13988 19196 14028
rect 20533 14025 20545 14028
rect 20579 14025 20591 14059
rect 21266 14056 21272 14068
rect 21227 14028 21272 14056
rect 20533 14019 20591 14025
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 21818 14016 21824 14068
rect 21876 14056 21882 14068
rect 24210 14056 24216 14068
rect 21876 14028 22324 14056
rect 24171 14028 24216 14056
rect 21876 14016 21882 14028
rect 18932 13960 19196 13988
rect 18932 13948 18938 13960
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5500 13892 5641 13920
rect 5500 13880 5506 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 6362 13920 6368 13932
rect 5859 13892 6368 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 12437 13923 12495 13929
rect 12437 13920 12449 13923
rect 11992 13892 12449 13920
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 2038 13852 2044 13864
rect 1951 13824 2044 13852
rect 2038 13812 2044 13824
rect 2096 13852 2102 13864
rect 2774 13852 2780 13864
rect 2096 13824 2780 13852
rect 2096 13812 2102 13824
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13821 8999 13855
rect 8941 13815 8999 13821
rect 2792 13716 2820 13812
rect 2869 13787 2927 13793
rect 2869 13753 2881 13787
rect 2915 13784 2927 13787
rect 3234 13784 3240 13796
rect 2915 13756 3240 13784
rect 2915 13753 2927 13756
rect 2869 13747 2927 13753
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 5074 13744 5080 13796
rect 5132 13784 5138 13796
rect 5537 13787 5595 13793
rect 5537 13784 5549 13787
rect 5132 13756 5549 13784
rect 5132 13744 5138 13756
rect 5537 13753 5549 13756
rect 5583 13753 5595 13787
rect 5537 13747 5595 13753
rect 8110 13744 8116 13796
rect 8168 13784 8174 13796
rect 8956 13784 8984 13815
rect 11992 13796 12020 13892
rect 12437 13889 12449 13892
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15746 13920 15752 13932
rect 14875 13892 15752 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 15838 13880 15844 13932
rect 15896 13920 15902 13932
rect 17497 13923 17555 13929
rect 15896 13892 15989 13920
rect 15896 13880 15902 13892
rect 17497 13889 17509 13923
rect 17543 13920 17555 13923
rect 18230 13920 18236 13932
rect 17543 13892 18236 13920
rect 17543 13889 17555 13892
rect 17497 13883 17555 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 20772 13892 21833 13920
rect 20772 13880 20778 13892
rect 21821 13889 21833 13892
rect 21867 13920 21879 13923
rect 22002 13920 22008 13932
rect 21867 13892 22008 13920
rect 21867 13889 21879 13892
rect 21821 13883 21879 13889
rect 22002 13880 22008 13892
rect 22060 13880 22066 13932
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 12693 13855 12751 13861
rect 12693 13852 12705 13855
rect 12584 13824 12705 13852
rect 12584 13812 12590 13824
rect 12693 13821 12705 13824
rect 12739 13852 12751 13855
rect 15654 13852 15660 13864
rect 12739 13824 13768 13852
rect 15615 13824 15660 13852
rect 12739 13821 12751 13824
rect 12693 13815 12751 13821
rect 8168 13756 8984 13784
rect 8168 13744 8174 13756
rect 2961 13719 3019 13725
rect 2961 13716 2973 13719
rect 2792 13688 2973 13716
rect 2961 13685 2973 13688
rect 3007 13685 3019 13719
rect 5166 13716 5172 13728
rect 5127 13688 5172 13716
rect 2961 13679 3019 13685
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 5626 13676 5632 13728
rect 5684 13716 5690 13728
rect 6181 13719 6239 13725
rect 6181 13716 6193 13719
rect 5684 13688 6193 13716
rect 5684 13676 5690 13688
rect 6181 13685 6193 13688
rect 6227 13685 6239 13719
rect 8956 13716 8984 13756
rect 9030 13744 9036 13796
rect 9088 13784 9094 13796
rect 9186 13787 9244 13793
rect 9186 13784 9198 13787
rect 9088 13756 9198 13784
rect 9088 13744 9094 13756
rect 9186 13753 9198 13756
rect 9232 13753 9244 13787
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 9186 13747 9244 13753
rect 9600 13756 11805 13784
rect 9600 13728 9628 13756
rect 11793 13753 11805 13756
rect 11839 13784 11851 13787
rect 11974 13784 11980 13796
rect 11839 13756 11980 13784
rect 11839 13753 11851 13756
rect 11793 13747 11851 13753
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 13740 13784 13768 13824
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 17865 13855 17923 13861
rect 17865 13821 17877 13855
rect 17911 13852 17923 13855
rect 18690 13852 18696 13864
rect 17911 13824 18696 13852
rect 17911 13821 17923 13824
rect 17865 13815 17923 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 19150 13852 19156 13864
rect 19111 13824 19156 13852
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 21174 13812 21180 13864
rect 21232 13852 21238 13864
rect 22296 13861 22324 14028
rect 24210 14016 24216 14028
rect 24268 14016 24274 14068
rect 24228 13920 24256 14016
rect 26697 13991 26755 13997
rect 26697 13957 26709 13991
rect 26743 13988 26755 13991
rect 26878 13988 26884 14000
rect 26743 13960 26884 13988
rect 26743 13957 26755 13960
rect 26697 13951 26755 13957
rect 26878 13948 26884 13960
rect 26936 13948 26942 14000
rect 24228 13892 24440 13920
rect 21545 13855 21603 13861
rect 21545 13852 21557 13855
rect 21232 13824 21557 13852
rect 21232 13812 21238 13824
rect 21545 13821 21557 13824
rect 21591 13821 21603 13855
rect 21545 13815 21603 13821
rect 22281 13855 22339 13861
rect 22281 13821 22293 13855
rect 22327 13852 22339 13855
rect 23382 13852 23388 13864
rect 22327 13824 23388 13852
rect 22327 13821 22339 13824
rect 22281 13815 22339 13821
rect 23382 13812 23388 13824
rect 23440 13812 23446 13864
rect 24302 13852 24308 13864
rect 23584 13824 24308 13852
rect 16669 13787 16727 13793
rect 16669 13784 16681 13787
rect 13740 13756 16681 13784
rect 16669 13753 16681 13756
rect 16715 13784 16727 13787
rect 16850 13784 16856 13796
rect 16715 13756 16856 13784
rect 16715 13753 16727 13756
rect 16669 13747 16727 13753
rect 16850 13744 16856 13756
rect 16908 13744 16914 13796
rect 19058 13744 19064 13796
rect 19116 13784 19122 13796
rect 19426 13793 19432 13796
rect 19398 13787 19432 13793
rect 19398 13784 19410 13787
rect 19116 13756 19410 13784
rect 19116 13744 19122 13756
rect 19398 13753 19410 13756
rect 19484 13784 19490 13796
rect 23584 13784 23612 13824
rect 24302 13812 24308 13824
rect 24360 13812 24366 13864
rect 24412 13852 24440 13892
rect 24561 13855 24619 13861
rect 24561 13852 24573 13855
rect 24412 13824 24573 13852
rect 24561 13821 24573 13824
rect 24607 13821 24619 13855
rect 26510 13852 26516 13864
rect 26471 13824 26516 13852
rect 24561 13815 24619 13821
rect 26510 13812 26516 13824
rect 26568 13852 26574 13864
rect 27065 13855 27123 13861
rect 27065 13852 27077 13855
rect 26568 13824 27077 13852
rect 26568 13812 26574 13824
rect 27065 13821 27077 13824
rect 27111 13821 27123 13855
rect 27065 13815 27123 13821
rect 19484 13756 19546 13784
rect 23400 13756 23612 13784
rect 19398 13747 19432 13753
rect 19426 13744 19432 13747
rect 19484 13744 19490 13756
rect 9582 13716 9588 13728
rect 8956 13688 9588 13716
rect 6181 13679 6239 13685
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 21361 13719 21419 13725
rect 21361 13685 21373 13719
rect 21407 13716 21419 13719
rect 21542 13716 21548 13728
rect 21407 13688 21548 13716
rect 21407 13685 21419 13688
rect 21361 13679 21419 13685
rect 21542 13676 21548 13688
rect 21600 13716 21606 13728
rect 21637 13719 21695 13725
rect 21637 13716 21649 13719
rect 21600 13688 21649 13716
rect 21600 13676 21606 13688
rect 21637 13685 21649 13688
rect 21683 13685 21695 13719
rect 21637 13679 21695 13685
rect 21729 13719 21787 13725
rect 21729 13685 21741 13719
rect 21775 13716 21787 13719
rect 23400 13716 23428 13756
rect 21775 13688 23428 13716
rect 25685 13719 25743 13725
rect 21775 13685 21787 13688
rect 21729 13679 21787 13685
rect 25685 13685 25697 13719
rect 25731 13716 25743 13719
rect 25866 13716 25872 13728
rect 25731 13688 25872 13716
rect 25731 13685 25743 13688
rect 25685 13679 25743 13685
rect 25866 13676 25872 13688
rect 25924 13676 25930 13728
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 2958 13512 2964 13524
rect 2919 13484 2964 13512
rect 2958 13472 2964 13484
rect 3016 13472 3022 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 8205 13515 8263 13521
rect 8205 13481 8217 13515
rect 8251 13512 8263 13515
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 8251 13484 9413 13512
rect 8251 13481 8263 13484
rect 8205 13475 8263 13481
rect 9401 13481 9413 13484
rect 9447 13512 9459 13515
rect 9490 13512 9496 13524
rect 9447 13484 9496 13512
rect 9447 13481 9459 13484
rect 9401 13475 9459 13481
rect 1486 13336 1492 13388
rect 1544 13376 1550 13388
rect 1581 13379 1639 13385
rect 1581 13376 1593 13379
rect 1544 13348 1593 13376
rect 1544 13336 1550 13348
rect 1581 13345 1593 13348
rect 1627 13345 1639 13379
rect 1581 13339 1639 13345
rect 1848 13379 1906 13385
rect 1848 13345 1860 13379
rect 1894 13376 1906 13379
rect 2314 13376 2320 13388
rect 1894 13348 2320 13376
rect 1894 13345 1906 13348
rect 1848 13339 1906 13345
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 5626 13376 5632 13388
rect 5587 13348 5632 13376
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13376 7067 13379
rect 7098 13376 7104 13388
rect 7055 13348 7104 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 7098 13336 7104 13348
rect 7156 13376 7162 13388
rect 8220 13376 8248 13475
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 13320 13484 13645 13512
rect 13320 13472 13326 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 17218 13512 17224 13524
rect 17179 13484 17224 13512
rect 13633 13475 13691 13481
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 18417 13515 18475 13521
rect 18417 13481 18429 13515
rect 18463 13512 18475 13515
rect 18782 13512 18788 13524
rect 18463 13484 18788 13512
rect 18463 13481 18475 13484
rect 18417 13475 18475 13481
rect 18782 13472 18788 13484
rect 18840 13472 18846 13524
rect 21358 13512 21364 13524
rect 21319 13484 21364 13512
rect 21358 13472 21364 13484
rect 21416 13472 21422 13524
rect 23106 13512 23112 13524
rect 23067 13484 23112 13512
rect 23106 13472 23112 13484
rect 23164 13472 23170 13524
rect 25222 13512 25228 13524
rect 25183 13484 25228 13512
rect 25222 13472 25228 13484
rect 25280 13472 25286 13524
rect 12250 13453 12256 13456
rect 12244 13444 12256 13453
rect 12211 13416 12256 13444
rect 12244 13407 12256 13416
rect 12250 13404 12256 13407
rect 12308 13404 12314 13456
rect 16850 13404 16856 13456
rect 16908 13444 16914 13456
rect 16908 13416 17356 13444
rect 16908 13404 16914 13416
rect 7156 13348 8248 13376
rect 8389 13379 8447 13385
rect 7156 13336 7162 13348
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 8478 13376 8484 13388
rect 8435 13348 8484 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8478 13336 8484 13348
rect 8536 13336 8542 13388
rect 11974 13376 11980 13388
rect 11935 13348 11980 13376
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 15105 13379 15163 13385
rect 15105 13345 15117 13379
rect 15151 13376 15163 13379
rect 15470 13376 15476 13388
rect 15151 13348 15476 13376
rect 15151 13345 15163 13348
rect 15105 13339 15163 13345
rect 15470 13336 15476 13348
rect 15528 13376 15534 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15528 13348 15669 13376
rect 15528 13336 15534 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 17328 13376 17356 13416
rect 25314 13404 25320 13456
rect 25372 13404 25378 13456
rect 19153 13379 19211 13385
rect 15804 13348 16896 13376
rect 17328 13348 17448 13376
rect 15804 13336 15810 13348
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13308 5135 13311
rect 5534 13308 5540 13320
rect 5123 13280 5540 13308
rect 5123 13277 5135 13280
rect 5077 13271 5135 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13308 5963 13311
rect 6270 13308 6276 13320
rect 5951 13280 6276 13308
rect 5951 13277 5963 13280
rect 5905 13271 5963 13277
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 15838 13308 15844 13320
rect 15799 13280 15844 13308
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 16868 13249 16896 13348
rect 17310 13308 17316 13320
rect 17271 13280 17316 13308
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 17420 13317 17448 13348
rect 19153 13345 19165 13379
rect 19199 13376 19211 13379
rect 19518 13376 19524 13388
rect 19199 13348 19524 13376
rect 19199 13345 19211 13348
rect 19153 13339 19211 13345
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 21542 13336 21548 13388
rect 21600 13376 21606 13388
rect 21729 13379 21787 13385
rect 21729 13376 21741 13379
rect 21600 13348 21741 13376
rect 21600 13336 21606 13348
rect 21729 13345 21741 13348
rect 21775 13345 21787 13379
rect 21729 13339 21787 13345
rect 21818 13336 21824 13388
rect 21876 13376 21882 13388
rect 21985 13379 22043 13385
rect 21985 13376 21997 13379
rect 21876 13348 21997 13376
rect 21876 13336 21882 13348
rect 21985 13345 21997 13348
rect 22031 13345 22043 13379
rect 25332 13376 25360 13404
rect 25332 13348 25452 13376
rect 21985 13339 22043 13345
rect 17405 13311 17463 13317
rect 17405 13277 17417 13311
rect 17451 13277 17463 13311
rect 19242 13308 19248 13320
rect 19203 13280 19248 13308
rect 17405 13271 17463 13277
rect 19242 13268 19248 13280
rect 19300 13268 19306 13320
rect 19426 13308 19432 13320
rect 19387 13280 19432 13308
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 25314 13308 25320 13320
rect 25275 13280 25320 13308
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 6825 13243 6883 13249
rect 6825 13240 6837 13243
rect 5408 13212 6837 13240
rect 5408 13200 5414 13212
rect 6825 13209 6837 13212
rect 6871 13209 6883 13243
rect 6825 13203 6883 13209
rect 16853 13243 16911 13249
rect 16853 13209 16865 13243
rect 16899 13209 16911 13243
rect 16853 13203 16911 13209
rect 18690 13200 18696 13252
rect 18748 13240 18754 13252
rect 18785 13243 18843 13249
rect 18785 13240 18797 13243
rect 18748 13212 18797 13240
rect 18748 13200 18754 13212
rect 18785 13209 18797 13212
rect 18831 13209 18843 13243
rect 25424 13240 25452 13348
rect 25501 13311 25559 13317
rect 25501 13277 25513 13311
rect 25547 13308 25559 13311
rect 25547 13280 25912 13308
rect 25547 13277 25559 13280
rect 25501 13271 25559 13277
rect 25774 13240 25780 13252
rect 25424 13212 25780 13240
rect 18785 13203 18843 13209
rect 25774 13200 25780 13212
rect 25832 13200 25838 13252
rect 25884 13184 25912 13280
rect 3234 13172 3240 13184
rect 3195 13144 3240 13172
rect 3234 13132 3240 13144
rect 3292 13132 3298 13184
rect 5261 13175 5319 13181
rect 5261 13141 5273 13175
rect 5307 13172 5319 13175
rect 5442 13172 5448 13184
rect 5307 13144 5448 13172
rect 5307 13141 5319 13144
rect 5261 13135 5319 13141
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 9030 13172 9036 13184
rect 8991 13144 9036 13172
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 9953 13175 10011 13181
rect 9953 13141 9965 13175
rect 9999 13172 10011 13175
rect 10134 13172 10140 13184
rect 9999 13144 10140 13172
rect 9999 13141 10011 13144
rect 9953 13135 10011 13141
rect 10134 13132 10140 13144
rect 10192 13172 10198 13184
rect 10778 13172 10784 13184
rect 10192 13144 10784 13172
rect 10192 13132 10198 13144
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 13354 13172 13360 13184
rect 13315 13144 13360 13172
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 15289 13175 15347 13181
rect 15289 13172 15301 13175
rect 14332 13144 15301 13172
rect 14332 13132 14338 13144
rect 15289 13141 15301 13144
rect 15335 13141 15347 13175
rect 15289 13135 15347 13141
rect 24305 13175 24363 13181
rect 24305 13141 24317 13175
rect 24351 13172 24363 13175
rect 24670 13172 24676 13184
rect 24351 13144 24676 13172
rect 24351 13141 24363 13144
rect 24305 13135 24363 13141
rect 24670 13132 24676 13144
rect 24728 13172 24734 13184
rect 24857 13175 24915 13181
rect 24857 13172 24869 13175
rect 24728 13144 24869 13172
rect 24728 13132 24734 13144
rect 24857 13141 24869 13144
rect 24903 13141 24915 13175
rect 25866 13172 25872 13184
rect 25827 13144 25872 13172
rect 24857 13135 24915 13141
rect 25866 13132 25872 13144
rect 25924 13132 25930 13184
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 2041 12971 2099 12977
rect 2041 12937 2053 12971
rect 2087 12968 2099 12971
rect 2130 12968 2136 12980
rect 2087 12940 2136 12968
rect 2087 12937 2099 12940
rect 2041 12931 2099 12937
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 2056 12764 2084 12931
rect 2130 12928 2136 12940
rect 2188 12928 2194 12980
rect 2314 12968 2320 12980
rect 2275 12940 2320 12968
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 4798 12968 4804 12980
rect 4759 12940 4804 12968
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 4985 12971 5043 12977
rect 4985 12937 4997 12971
rect 5031 12968 5043 12971
rect 5074 12968 5080 12980
rect 5031 12940 5080 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5997 12971 6055 12977
rect 5997 12968 6009 12971
rect 5776 12940 6009 12968
rect 5776 12928 5782 12940
rect 5997 12937 6009 12940
rect 6043 12937 6055 12971
rect 5997 12931 6055 12937
rect 4246 12860 4252 12912
rect 4304 12900 4310 12912
rect 4525 12903 4583 12909
rect 4525 12900 4537 12903
rect 4304 12872 4537 12900
rect 4304 12860 4310 12872
rect 4525 12869 4537 12872
rect 4571 12900 4583 12903
rect 5626 12900 5632 12912
rect 4571 12872 5632 12900
rect 4571 12869 4583 12872
rect 4525 12863 4583 12869
rect 5626 12860 5632 12872
rect 5684 12860 5690 12912
rect 6012 12900 6040 12931
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 6328 12940 6377 12968
rect 6328 12928 6334 12940
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 7098 12968 7104 12980
rect 7059 12940 7104 12968
rect 6365 12931 6423 12937
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9769 12971 9827 12977
rect 9769 12968 9781 12971
rect 9732 12940 9781 12968
rect 9732 12928 9738 12940
rect 9769 12937 9781 12940
rect 9815 12937 9827 12971
rect 9769 12931 9827 12937
rect 12069 12971 12127 12977
rect 12069 12937 12081 12971
rect 12115 12968 12127 12971
rect 12250 12968 12256 12980
rect 12115 12940 12256 12968
rect 12115 12937 12127 12940
rect 12069 12931 12127 12937
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 13722 12968 13728 12980
rect 13412 12940 13728 12968
rect 13412 12928 13418 12940
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 15470 12968 15476 12980
rect 15431 12940 15476 12968
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 16577 12971 16635 12977
rect 16577 12937 16589 12971
rect 16623 12968 16635 12971
rect 16850 12968 16856 12980
rect 16623 12940 16856 12968
rect 16623 12937 16635 12940
rect 16577 12931 16635 12937
rect 6454 12900 6460 12912
rect 6012 12872 6460 12900
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 11974 12860 11980 12912
rect 12032 12900 12038 12912
rect 12621 12903 12679 12909
rect 12621 12900 12633 12903
rect 12032 12872 12633 12900
rect 12032 12860 12038 12872
rect 12621 12869 12633 12872
rect 12667 12900 12679 12903
rect 12802 12900 12808 12912
rect 12667 12872 12808 12900
rect 12667 12869 12679 12872
rect 12621 12863 12679 12869
rect 12802 12860 12808 12872
rect 12860 12860 12866 12912
rect 15381 12903 15439 12909
rect 15381 12869 15393 12903
rect 15427 12900 15439 12903
rect 15562 12900 15568 12912
rect 15427 12872 15568 12900
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 15562 12860 15568 12872
rect 15620 12900 15626 12912
rect 15620 12872 15976 12900
rect 15620 12860 15626 12872
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12832 4215 12835
rect 5442 12832 5448 12844
rect 4203 12804 5448 12832
rect 4203 12801 4215 12804
rect 4157 12795 4215 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 5718 12832 5724 12844
rect 5592 12804 5724 12832
rect 5592 12792 5598 12804
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 8110 12832 8116 12844
rect 8071 12804 8116 12832
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 13722 12792 13728 12844
rect 13780 12832 13786 12844
rect 15948 12841 15976 12872
rect 14461 12835 14519 12841
rect 14461 12832 14473 12835
rect 13780 12804 14473 12832
rect 13780 12792 13786 12804
rect 14461 12801 14473 12804
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12801 15991 12835
rect 15933 12795 15991 12801
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12832 16175 12835
rect 16592 12832 16620 12931
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17310 12968 17316 12980
rect 17271 12940 17316 12968
rect 17310 12928 17316 12940
rect 17368 12928 17374 12980
rect 18782 12968 18788 12980
rect 18743 12940 18788 12968
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 21818 12968 21824 12980
rect 21779 12940 21824 12968
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 25314 12968 25320 12980
rect 25275 12940 25320 12968
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 16868 12900 16896 12928
rect 17589 12903 17647 12909
rect 17589 12900 17601 12903
rect 16868 12872 17601 12900
rect 17589 12869 17601 12872
rect 17635 12869 17647 12903
rect 17589 12863 17647 12869
rect 19518 12860 19524 12912
rect 19576 12900 19582 12912
rect 19797 12903 19855 12909
rect 19797 12900 19809 12903
rect 19576 12872 19809 12900
rect 19576 12860 19582 12872
rect 19797 12869 19809 12872
rect 19843 12869 19855 12903
rect 19797 12863 19855 12869
rect 21542 12860 21548 12912
rect 21600 12900 21606 12912
rect 22097 12903 22155 12909
rect 22097 12900 22109 12903
rect 21600 12872 22109 12900
rect 21600 12860 21606 12872
rect 22097 12869 22109 12872
rect 22143 12869 22155 12903
rect 22097 12863 22155 12869
rect 24302 12860 24308 12912
rect 24360 12900 24366 12912
rect 24360 12872 24900 12900
rect 24360 12860 24366 12872
rect 16163 12804 16620 12832
rect 16945 12835 17003 12841
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 16945 12801 16957 12835
rect 16991 12832 17003 12835
rect 17218 12832 17224 12844
rect 16991 12804 17224 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 17218 12792 17224 12804
rect 17276 12792 17282 12844
rect 19426 12832 19432 12844
rect 19387 12804 19432 12832
rect 19426 12792 19432 12804
rect 19484 12832 19490 12844
rect 20165 12835 20223 12841
rect 20165 12832 20177 12835
rect 19484 12804 20177 12832
rect 19484 12792 19490 12804
rect 20165 12801 20177 12804
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 23934 12792 23940 12844
rect 23992 12832 23998 12844
rect 24029 12835 24087 12841
rect 24029 12832 24041 12835
rect 23992 12804 24041 12832
rect 23992 12792 23998 12804
rect 24029 12801 24041 12804
rect 24075 12801 24087 12835
rect 24029 12795 24087 12801
rect 1443 12736 2084 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 5350 12764 5356 12776
rect 4856 12736 5356 12764
rect 4856 12724 4862 12736
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 13449 12767 13507 12773
rect 13449 12733 13461 12767
rect 13495 12764 13507 12767
rect 14274 12764 14280 12776
rect 13495 12736 14280 12764
rect 13495 12733 13507 12736
rect 13449 12727 13507 12733
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14366 12724 14372 12776
rect 14424 12764 14430 12776
rect 15102 12764 15108 12776
rect 14424 12736 15108 12764
rect 14424 12724 14430 12736
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 24044 12764 24072 12795
rect 24394 12792 24400 12844
rect 24452 12832 24458 12844
rect 24765 12835 24823 12841
rect 24765 12832 24777 12835
rect 24452 12804 24777 12832
rect 24452 12792 24458 12804
rect 24765 12801 24777 12804
rect 24811 12801 24823 12835
rect 24765 12795 24823 12801
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 24044 12736 24593 12764
rect 24581 12733 24593 12736
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 24670 12724 24676 12776
rect 24728 12764 24734 12776
rect 24872 12764 24900 12872
rect 25222 12860 25228 12912
rect 25280 12900 25286 12912
rect 25593 12903 25651 12909
rect 25593 12900 25605 12903
rect 25280 12872 25605 12900
rect 25280 12860 25286 12872
rect 25593 12869 25605 12872
rect 25639 12869 25651 12903
rect 25593 12863 25651 12869
rect 25314 12792 25320 12844
rect 25372 12832 25378 12844
rect 25498 12832 25504 12844
rect 25372 12804 25504 12832
rect 25372 12792 25378 12804
rect 25498 12792 25504 12804
rect 25556 12792 25562 12844
rect 25777 12767 25835 12773
rect 25777 12764 25789 12767
rect 24728 12736 24773 12764
rect 24872 12736 25789 12764
rect 24728 12724 24734 12736
rect 25777 12733 25789 12736
rect 25823 12764 25835 12767
rect 25823 12736 26188 12764
rect 25823 12733 25835 12736
rect 25777 12727 25835 12733
rect 26160 12708 26188 12736
rect 1486 12656 1492 12708
rect 1544 12696 1550 12708
rect 2682 12696 2688 12708
rect 1544 12668 2688 12696
rect 1544 12656 1550 12668
rect 2682 12656 2688 12668
rect 2740 12656 2746 12708
rect 7926 12656 7932 12708
rect 7984 12696 7990 12708
rect 8021 12699 8079 12705
rect 8021 12696 8033 12699
rect 7984 12668 8033 12696
rect 7984 12656 7990 12668
rect 8021 12665 8033 12668
rect 8067 12696 8079 12699
rect 8358 12699 8416 12705
rect 8358 12696 8370 12699
rect 8067 12668 8370 12696
rect 8067 12665 8079 12668
rect 8021 12659 8079 12665
rect 8358 12665 8370 12668
rect 8404 12665 8416 12699
rect 8358 12659 8416 12665
rect 8478 12656 8484 12708
rect 8536 12696 8542 12708
rect 9214 12696 9220 12708
rect 8536 12668 9220 12696
rect 8536 12656 8542 12668
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 14458 12696 14464 12708
rect 13924 12668 14464 12696
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 7653 12631 7711 12637
rect 7653 12597 7665 12631
rect 7699 12628 7711 12631
rect 8496 12628 8524 12656
rect 7699 12600 8524 12628
rect 7699 12597 7711 12600
rect 7653 12591 7711 12597
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 13924 12637 13952 12668
rect 14458 12656 14464 12668
rect 14516 12656 14522 12708
rect 15013 12699 15071 12705
rect 15013 12665 15025 12699
rect 15059 12696 15071 12699
rect 15562 12696 15568 12708
rect 15059 12668 15568 12696
rect 15059 12665 15071 12668
rect 15013 12659 15071 12665
rect 15562 12656 15568 12668
rect 15620 12696 15626 12708
rect 15841 12699 15899 12705
rect 15841 12696 15853 12699
rect 15620 12668 15853 12696
rect 15620 12656 15626 12668
rect 15841 12665 15853 12668
rect 15887 12665 15899 12699
rect 15841 12659 15899 12665
rect 18693 12699 18751 12705
rect 18693 12665 18705 12699
rect 18739 12696 18751 12699
rect 18966 12696 18972 12708
rect 18739 12668 18972 12696
rect 18739 12665 18751 12668
rect 18693 12659 18751 12665
rect 18966 12656 18972 12668
rect 19024 12696 19030 12708
rect 19245 12699 19303 12705
rect 19245 12696 19257 12699
rect 19024 12668 19257 12696
rect 19024 12656 19030 12668
rect 19245 12665 19257 12668
rect 19291 12665 19303 12699
rect 19245 12659 19303 12665
rect 25498 12656 25504 12708
rect 25556 12696 25562 12708
rect 25866 12696 25872 12708
rect 25556 12668 25872 12696
rect 25556 12656 25562 12668
rect 25866 12656 25872 12668
rect 25924 12696 25930 12708
rect 26022 12699 26080 12705
rect 26022 12696 26034 12699
rect 25924 12668 26034 12696
rect 25924 12656 25930 12668
rect 26022 12665 26034 12668
rect 26068 12665 26080 12699
rect 26022 12659 26080 12665
rect 26142 12656 26148 12708
rect 26200 12656 26206 12708
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 9088 12600 9505 12628
rect 9088 12588 9094 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 9493 12591 9551 12597
rect 13909 12631 13967 12637
rect 13909 12597 13921 12631
rect 13955 12597 13967 12631
rect 13909 12591 13967 12597
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18325 12631 18383 12637
rect 18325 12628 18337 12631
rect 18012 12600 18337 12628
rect 18012 12588 18018 12600
rect 18325 12597 18337 12600
rect 18371 12628 18383 12631
rect 19153 12631 19211 12637
rect 19153 12628 19165 12631
rect 18371 12600 19165 12628
rect 18371 12597 18383 12600
rect 18325 12591 18383 12597
rect 19153 12597 19165 12600
rect 19199 12597 19211 12631
rect 19153 12591 19211 12597
rect 24213 12631 24271 12637
rect 24213 12597 24225 12631
rect 24259 12628 24271 12631
rect 24302 12628 24308 12640
rect 24259 12600 24308 12628
rect 24259 12597 24271 12600
rect 24213 12591 24271 12597
rect 24302 12588 24308 12600
rect 24360 12588 24366 12640
rect 27154 12628 27160 12640
rect 27115 12600 27160 12628
rect 27154 12588 27160 12600
rect 27212 12588 27218 12640
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 2314 12384 2320 12436
rect 2372 12424 2378 12436
rect 6362 12424 6368 12436
rect 2372 12396 2820 12424
rect 6323 12396 6368 12424
rect 2372 12384 2378 12396
rect 2792 12368 2820 12396
rect 6362 12384 6368 12396
rect 6420 12424 6426 12436
rect 7742 12424 7748 12436
rect 6420 12396 7748 12424
rect 6420 12384 6426 12396
rect 7742 12384 7748 12396
rect 7800 12424 7806 12436
rect 7926 12424 7932 12436
rect 7800 12396 7932 12424
rect 7800 12384 7806 12396
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 12802 12424 12808 12436
rect 12763 12396 12808 12424
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 14001 12427 14059 12433
rect 14001 12393 14013 12427
rect 14047 12424 14059 12427
rect 14366 12424 14372 12436
rect 14047 12396 14372 12424
rect 14047 12393 14059 12396
rect 14001 12387 14059 12393
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 15562 12424 15568 12436
rect 15523 12396 15568 12424
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 16025 12427 16083 12433
rect 16025 12424 16037 12427
rect 15896 12396 16037 12424
rect 15896 12384 15902 12396
rect 16025 12393 16037 12396
rect 16071 12393 16083 12427
rect 16025 12387 16083 12393
rect 17589 12427 17647 12433
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 17678 12424 17684 12436
rect 17635 12396 17684 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 18230 12384 18236 12436
rect 18288 12424 18294 12436
rect 19061 12427 19119 12433
rect 19061 12424 19073 12427
rect 18288 12396 19073 12424
rect 18288 12384 18294 12396
rect 19061 12393 19073 12396
rect 19107 12393 19119 12427
rect 19061 12387 19119 12393
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19521 12427 19579 12433
rect 19521 12424 19533 12427
rect 19484 12396 19533 12424
rect 19484 12384 19490 12396
rect 19521 12393 19533 12396
rect 19567 12393 19579 12427
rect 19521 12387 19579 12393
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 24857 12427 24915 12433
rect 24857 12424 24869 12427
rect 23532 12396 24869 12424
rect 23532 12384 23538 12396
rect 24857 12393 24869 12396
rect 24903 12424 24915 12427
rect 25038 12424 25044 12436
rect 24903 12396 25044 12424
rect 24903 12393 24915 12396
rect 24857 12387 24915 12393
rect 25038 12384 25044 12396
rect 25096 12384 25102 12436
rect 25498 12424 25504 12436
rect 25459 12396 25504 12424
rect 25498 12384 25504 12396
rect 25556 12384 25562 12436
rect 25590 12384 25596 12436
rect 25648 12384 25654 12436
rect 26234 12424 26240 12436
rect 26195 12396 26240 12424
rect 26234 12384 26240 12396
rect 26292 12384 26298 12436
rect 2774 12316 2780 12368
rect 2832 12316 2838 12368
rect 15105 12359 15163 12365
rect 15105 12325 15117 12359
rect 15151 12356 15163 12359
rect 15746 12356 15752 12368
rect 15151 12328 15752 12356
rect 15151 12325 15163 12328
rect 15105 12319 15163 12325
rect 15746 12316 15752 12328
rect 15804 12316 15810 12368
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1486 12288 1492 12300
rect 1443 12260 1492 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1486 12248 1492 12260
rect 1544 12248 1550 12300
rect 1670 12297 1676 12300
rect 1664 12251 1676 12297
rect 1728 12288 1734 12300
rect 1728 12260 1764 12288
rect 1670 12248 1676 12251
rect 1728 12248 1734 12260
rect 2682 12248 2688 12300
rect 2740 12288 2746 12300
rect 4982 12288 4988 12300
rect 2740 12260 4988 12288
rect 2740 12248 2746 12260
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 5252 12291 5310 12297
rect 5252 12257 5264 12291
rect 5298 12288 5310 12291
rect 5718 12288 5724 12300
rect 5298 12260 5724 12288
rect 5298 12257 5310 12260
rect 5252 12251 5310 12257
rect 5718 12248 5724 12260
rect 5776 12288 5782 12300
rect 5776 12260 6316 12288
rect 5776 12248 5782 12260
rect 6288 12164 6316 12260
rect 7834 12248 7840 12300
rect 7892 12288 7898 12300
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 7892 12260 8401 12288
rect 7892 12248 7898 12260
rect 8389 12257 8401 12260
rect 8435 12257 8447 12291
rect 8389 12251 8447 12257
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10594 12288 10600 12300
rect 10091 12260 10600 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12288 17555 12291
rect 17770 12288 17776 12300
rect 17543 12260 17776 12288
rect 17543 12257 17555 12260
rect 17497 12251 17555 12257
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 18874 12248 18880 12300
rect 18932 12288 18938 12300
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 18932 12260 19257 12288
rect 18932 12248 18938 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 21542 12248 21548 12300
rect 21600 12288 21606 12300
rect 21910 12297 21916 12300
rect 21637 12291 21695 12297
rect 21637 12288 21649 12291
rect 21600 12260 21649 12288
rect 21600 12248 21606 12260
rect 21637 12257 21649 12260
rect 21683 12257 21695 12291
rect 21904 12288 21916 12297
rect 21823 12260 21916 12288
rect 21637 12251 21695 12257
rect 21904 12251 21916 12260
rect 21968 12288 21974 12300
rect 24213 12291 24271 12297
rect 24213 12288 24225 12291
rect 21968 12260 24225 12288
rect 21910 12248 21916 12251
rect 21968 12248 21974 12260
rect 24213 12257 24225 12260
rect 24259 12288 24271 12291
rect 24394 12288 24400 12300
rect 24259 12260 24400 12288
rect 24259 12257 24271 12260
rect 24213 12251 24271 12257
rect 24394 12248 24400 12260
rect 24452 12248 24458 12300
rect 24762 12288 24768 12300
rect 24723 12260 24768 12288
rect 24762 12248 24768 12260
rect 24820 12248 24826 12300
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 8481 12223 8539 12229
rect 8481 12220 8493 12223
rect 7340 12192 8493 12220
rect 7340 12180 7346 12192
rect 8481 12189 8493 12192
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12220 8723 12223
rect 9030 12220 9036 12232
rect 8711 12192 9036 12220
rect 8711 12189 8723 12192
rect 8665 12183 8723 12189
rect 9030 12180 9036 12192
rect 9088 12180 9094 12232
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10008 12192 10149 12220
rect 10008 12180 10014 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12220 17739 12223
rect 17862 12220 17868 12232
rect 17727 12192 17868 12220
rect 17727 12189 17739 12192
rect 17681 12183 17739 12189
rect 6270 12112 6276 12164
rect 6328 12152 6334 12164
rect 9493 12155 9551 12161
rect 9493 12152 9505 12155
rect 6328 12124 9505 12152
rect 6328 12112 6334 12124
rect 9493 12121 9505 12124
rect 9539 12152 9551 12155
rect 9582 12152 9588 12164
rect 9539 12124 9588 12152
rect 9539 12121 9551 12124
rect 9493 12115 9551 12121
rect 9582 12112 9588 12124
rect 9640 12152 9646 12164
rect 10244 12152 10272 12183
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 24412 12220 24440 12248
rect 25608 12232 25636 12384
rect 24949 12223 25007 12229
rect 24949 12220 24961 12223
rect 24412 12192 24961 12220
rect 24949 12189 24961 12192
rect 24995 12189 25007 12223
rect 24949 12183 25007 12189
rect 25590 12180 25596 12232
rect 25648 12180 25654 12232
rect 26513 12223 26571 12229
rect 26513 12189 26525 12223
rect 26559 12220 26571 12223
rect 26878 12220 26884 12232
rect 26559 12192 26884 12220
rect 26559 12189 26571 12192
rect 26513 12183 26571 12189
rect 26878 12180 26884 12192
rect 26936 12180 26942 12232
rect 9640 12124 10272 12152
rect 23937 12155 23995 12161
rect 9640 12112 9646 12124
rect 23937 12121 23949 12155
rect 23983 12152 23995 12155
rect 24118 12152 24124 12164
rect 23983 12124 24124 12152
rect 23983 12121 23995 12124
rect 23937 12115 23995 12121
rect 24118 12112 24124 12124
rect 24176 12152 24182 12164
rect 24397 12155 24455 12161
rect 24397 12152 24409 12155
rect 24176 12124 24409 12152
rect 24176 12112 24182 12124
rect 24397 12121 24409 12124
rect 24443 12121 24455 12155
rect 24397 12115 24455 12121
rect 25682 12112 25688 12164
rect 25740 12152 25746 12164
rect 26602 12152 26608 12164
rect 25740 12124 26608 12152
rect 25740 12112 25746 12124
rect 26602 12112 26608 12124
rect 26660 12112 26666 12164
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 7926 12084 7932 12096
rect 2832 12056 2877 12084
rect 7887 12056 7932 12084
rect 2832 12044 2838 12056
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 8021 12087 8079 12093
rect 8021 12053 8033 12087
rect 8067 12084 8079 12087
rect 8110 12084 8116 12096
rect 8067 12056 8116 12084
rect 8067 12053 8079 12056
rect 8021 12047 8079 12053
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 9674 12084 9680 12096
rect 9635 12056 9680 12084
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 16482 12084 16488 12096
rect 16443 12056 16488 12084
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 17126 12084 17132 12096
rect 17087 12056 17132 12084
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 18877 12087 18935 12093
rect 18877 12053 18889 12087
rect 18923 12084 18935 12087
rect 19150 12084 19156 12096
rect 18923 12056 19156 12084
rect 18923 12053 18935 12056
rect 18877 12047 18935 12053
rect 19150 12044 19156 12056
rect 19208 12044 19214 12096
rect 23014 12084 23020 12096
rect 22975 12056 23020 12084
rect 23014 12044 23020 12056
rect 23072 12044 23078 12096
rect 24946 12044 24952 12096
rect 25004 12084 25010 12096
rect 25130 12084 25136 12096
rect 25004 12056 25136 12084
rect 25004 12044 25010 12056
rect 25130 12044 25136 12056
rect 25188 12044 25194 12096
rect 25866 12084 25872 12096
rect 25827 12056 25872 12084
rect 25866 12044 25872 12056
rect 25924 12044 25930 12096
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 2777 11883 2835 11889
rect 2777 11880 2789 11883
rect 2740 11852 2789 11880
rect 2740 11840 2746 11852
rect 2777 11849 2789 11852
rect 2823 11849 2835 11883
rect 2777 11843 2835 11849
rect 2792 11744 2820 11843
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5040 11852 5457 11880
rect 5040 11840 5046 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 5445 11843 5503 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 7742 11880 7748 11892
rect 7703 11852 7748 11880
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 8941 11883 8999 11889
rect 8941 11849 8953 11883
rect 8987 11880 8999 11883
rect 9030 11880 9036 11892
rect 8987 11852 9036 11880
rect 8987 11849 8999 11852
rect 8941 11843 8999 11849
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 17497 11883 17555 11889
rect 17497 11849 17509 11883
rect 17543 11880 17555 11883
rect 17678 11880 17684 11892
rect 17543 11852 17684 11880
rect 17543 11849 17555 11852
rect 17497 11843 17555 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 17770 11840 17776 11892
rect 17828 11880 17834 11892
rect 17828 11852 18092 11880
rect 17828 11840 17834 11852
rect 4801 11815 4859 11821
rect 4801 11781 4813 11815
rect 4847 11812 4859 11815
rect 5258 11812 5264 11824
rect 4847 11784 5264 11812
rect 4847 11781 4859 11784
rect 4801 11775 4859 11781
rect 5258 11772 5264 11784
rect 5316 11772 5322 11824
rect 3418 11744 3424 11756
rect 2792 11716 3424 11744
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 6270 11744 6276 11756
rect 5215 11716 6276 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 6270 11704 6276 11716
rect 6328 11704 6334 11756
rect 7760 11744 7788 11840
rect 7926 11772 7932 11824
rect 7984 11812 7990 11824
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 7984 11784 9413 11812
rect 7984 11772 7990 11784
rect 9401 11781 9413 11784
rect 9447 11781 9459 11815
rect 9401 11775 9459 11781
rect 8389 11747 8447 11753
rect 8389 11744 8401 11747
rect 7760 11716 8401 11744
rect 8389 11713 8401 11716
rect 8435 11713 8447 11747
rect 8389 11707 8447 11713
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9640 11716 9965 11744
rect 9640 11704 9646 11716
rect 9953 11713 9965 11716
rect 9999 11744 10011 11747
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 9999 11716 10793 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 12802 11744 12808 11756
rect 12763 11716 12808 11744
rect 10781 11707 10839 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 15838 11704 15844 11756
rect 15896 11744 15902 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15896 11716 15945 11744
rect 15896 11704 15902 11716
rect 15933 11713 15945 11716
rect 15979 11744 15991 11747
rect 17037 11747 17095 11753
rect 17037 11744 17049 11747
rect 15979 11716 17049 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 17037 11713 17049 11716
rect 17083 11744 17095 11747
rect 17862 11744 17868 11756
rect 17083 11716 17868 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 18064 11753 18092 11852
rect 19426 11840 19432 11892
rect 19484 11880 19490 11892
rect 19610 11880 19616 11892
rect 19484 11852 19616 11880
rect 19484 11840 19490 11852
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 21729 11883 21787 11889
rect 21729 11849 21741 11883
rect 21775 11880 21787 11883
rect 21910 11880 21916 11892
rect 21775 11852 21916 11880
rect 21775 11849 21787 11852
rect 21729 11843 21787 11849
rect 21910 11840 21916 11852
rect 21968 11840 21974 11892
rect 24762 11840 24768 11892
rect 24820 11880 24826 11892
rect 24857 11883 24915 11889
rect 24857 11880 24869 11883
rect 24820 11852 24869 11880
rect 24820 11840 24826 11852
rect 24857 11849 24869 11852
rect 24903 11849 24915 11883
rect 24857 11843 24915 11849
rect 21542 11772 21548 11824
rect 21600 11812 21606 11824
rect 22005 11815 22063 11821
rect 22005 11812 22017 11815
rect 21600 11784 22017 11812
rect 21600 11772 21606 11784
rect 22005 11781 22017 11784
rect 22051 11781 22063 11815
rect 22005 11775 22063 11781
rect 23014 11772 23020 11824
rect 23072 11812 23078 11824
rect 23477 11815 23535 11821
rect 23477 11812 23489 11815
rect 23072 11784 23489 11812
rect 23072 11772 23078 11784
rect 23477 11781 23489 11784
rect 23523 11812 23535 11815
rect 24872 11812 24900 11843
rect 25038 11840 25044 11892
rect 25096 11880 25102 11892
rect 25225 11883 25283 11889
rect 25225 11880 25237 11883
rect 25096 11852 25237 11880
rect 25096 11840 25102 11852
rect 25225 11849 25237 11852
rect 25271 11849 25283 11883
rect 25225 11843 25283 11849
rect 26510 11812 26516 11824
rect 23523 11784 24532 11812
rect 24872 11784 26516 11812
rect 23523 11781 23535 11784
rect 23477 11775 23535 11781
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11713 18107 11747
rect 18598 11744 18604 11756
rect 18511 11716 18604 11744
rect 18049 11707 18107 11713
rect 18598 11704 18604 11716
rect 18656 11744 18662 11756
rect 19334 11744 19340 11756
rect 18656 11716 19340 11744
rect 18656 11704 18662 11716
rect 19334 11704 19340 11716
rect 19392 11744 19398 11756
rect 19429 11747 19487 11753
rect 19429 11744 19441 11747
rect 19392 11716 19441 11744
rect 19392 11704 19398 11716
rect 19429 11713 19441 11716
rect 19475 11713 19487 11747
rect 24302 11744 24308 11756
rect 24263 11716 24308 11744
rect 19429 11707 19487 11713
rect 24302 11704 24308 11716
rect 24360 11704 24366 11756
rect 24504 11753 24532 11784
rect 26510 11772 26516 11784
rect 26568 11772 26574 11824
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11744 24547 11747
rect 24946 11744 24952 11756
rect 24535 11716 24952 11744
rect 24535 11713 24547 11716
rect 24489 11707 24547 11713
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 25866 11704 25872 11756
rect 25924 11744 25930 11756
rect 26237 11747 26295 11753
rect 26237 11744 26249 11747
rect 25924 11716 26249 11744
rect 25924 11704 25930 11716
rect 26237 11713 26249 11716
rect 26283 11713 26295 11747
rect 26237 11707 26295 11713
rect 26329 11747 26387 11753
rect 26329 11713 26341 11747
rect 26375 11713 26387 11747
rect 26329 11707 26387 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1443 11648 1961 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1949 11645 1961 11648
rect 1995 11676 2007 11679
rect 7650 11676 7656 11688
rect 1995 11648 7656 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 7984 11648 8217 11676
rect 7984 11636 7990 11648
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 9674 11676 9680 11688
rect 8343 11648 9680 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 3666 11611 3724 11617
rect 3666 11608 3678 11611
rect 3344 11580 3678 11608
rect 3344 11552 3372 11580
rect 3666 11577 3678 11580
rect 3712 11577 3724 11611
rect 3666 11571 3724 11577
rect 8018 11568 8024 11620
rect 8076 11608 8082 11620
rect 8312 11608 8340 11639
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 16390 11676 16396 11688
rect 12636 11648 16396 11676
rect 8076 11580 8340 11608
rect 8076 11568 8082 11580
rect 8386 11568 8392 11620
rect 8444 11608 8450 11620
rect 9309 11611 9367 11617
rect 9309 11608 9321 11611
rect 8444 11580 9321 11608
rect 8444 11568 8450 11580
rect 9309 11577 9321 11580
rect 9355 11608 9367 11611
rect 9861 11611 9919 11617
rect 9861 11608 9873 11611
rect 9355 11580 9873 11608
rect 9355 11577 9367 11580
rect 9309 11571 9367 11577
rect 9861 11577 9873 11580
rect 9907 11608 9919 11611
rect 12636 11608 12664 11648
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 16853 11679 16911 11685
rect 16853 11676 16865 11679
rect 16540 11648 16865 11676
rect 16540 11636 16546 11648
rect 16853 11645 16865 11648
rect 16899 11645 16911 11679
rect 16853 11639 16911 11645
rect 24118 11636 24124 11688
rect 24176 11676 24182 11688
rect 24213 11679 24271 11685
rect 24213 11676 24225 11679
rect 24176 11648 24225 11676
rect 24176 11636 24182 11648
rect 24213 11645 24225 11648
rect 24259 11645 24271 11679
rect 24213 11639 24271 11645
rect 25958 11636 25964 11688
rect 26016 11676 26022 11688
rect 26344 11676 26372 11707
rect 26016 11648 26372 11676
rect 26016 11636 26022 11648
rect 9907 11580 12664 11608
rect 12713 11611 12771 11617
rect 9907 11577 9919 11580
rect 9861 11571 9919 11577
rect 12713 11577 12725 11611
rect 12759 11608 12771 11611
rect 13072 11611 13130 11617
rect 13072 11608 13084 11611
rect 12759 11580 13084 11608
rect 12759 11577 12771 11580
rect 12713 11571 12771 11577
rect 13072 11577 13084 11580
rect 13118 11608 13130 11611
rect 13722 11608 13728 11620
rect 13118 11580 13728 11608
rect 13118 11577 13130 11580
rect 13072 11571 13130 11577
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 16298 11608 16304 11620
rect 16211 11580 16304 11608
rect 16298 11568 16304 11580
rect 16356 11608 16362 11620
rect 19702 11617 19708 11620
rect 19337 11611 19395 11617
rect 16356 11580 16804 11608
rect 16356 11568 16362 11580
rect 16776 11552 16804 11580
rect 19337 11577 19349 11611
rect 19383 11608 19395 11611
rect 19696 11608 19708 11617
rect 19383 11580 19708 11608
rect 19383 11577 19395 11580
rect 19337 11571 19395 11577
rect 19696 11571 19708 11580
rect 19702 11568 19708 11571
rect 19760 11568 19766 11620
rect 26145 11611 26203 11617
rect 26145 11608 26157 11611
rect 25608 11580 26157 11608
rect 25608 11552 25636 11580
rect 26145 11577 26157 11580
rect 26191 11577 26203 11611
rect 26145 11571 26203 11577
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 2498 11540 2504 11552
rect 2459 11512 2504 11540
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 3326 11540 3332 11552
rect 3287 11512 3332 11540
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 7834 11540 7840 11552
rect 7795 11512 7840 11540
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9548 11512 9781 11540
rect 9548 11500 9554 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 9769 11503 9827 11509
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 10594 11540 10600 11552
rect 10551 11512 10600 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 10965 11543 11023 11549
rect 10965 11540 10977 11543
rect 10928 11512 10977 11540
rect 10928 11500 10934 11512
rect 10965 11509 10977 11512
rect 11011 11509 11023 11543
rect 10965 11503 11023 11509
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 14090 11540 14096 11552
rect 12952 11512 14096 11540
rect 12952 11500 12958 11512
rect 14090 11500 14096 11512
rect 14148 11540 14154 11552
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 14148 11512 14197 11540
rect 14148 11500 14154 11512
rect 14185 11509 14197 11512
rect 14231 11509 14243 11543
rect 16390 11540 16396 11552
rect 16351 11512 16396 11540
rect 14185 11503 14243 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 16758 11540 16764 11552
rect 16719 11512 16764 11540
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 18874 11540 18880 11552
rect 18835 11512 18880 11540
rect 18874 11500 18880 11512
rect 18932 11500 18938 11552
rect 20806 11540 20812 11552
rect 20767 11512 20812 11540
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 23842 11540 23848 11552
rect 23803 11512 23848 11540
rect 23842 11500 23848 11512
rect 23900 11500 23906 11552
rect 25590 11540 25596 11552
rect 25551 11512 25596 11540
rect 25590 11500 25596 11512
rect 25648 11500 25654 11552
rect 25774 11540 25780 11552
rect 25735 11512 25780 11540
rect 25774 11500 25780 11512
rect 25832 11500 25838 11552
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 2556 11308 2789 11336
rect 2556 11296 2562 11308
rect 2777 11305 2789 11308
rect 2823 11305 2835 11339
rect 2777 11299 2835 11305
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 4709 11339 4767 11345
rect 4709 11336 4721 11339
rect 2915 11308 4721 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 4709 11305 4721 11308
rect 4755 11305 4767 11339
rect 4709 11299 4767 11305
rect 7929 11339 7987 11345
rect 7929 11305 7941 11339
rect 7975 11336 7987 11339
rect 8018 11336 8024 11348
rect 7975 11308 8024 11336
rect 7975 11305 7987 11308
rect 7929 11299 7987 11305
rect 2317 11271 2375 11277
rect 2317 11237 2329 11271
rect 2363 11268 2375 11271
rect 2884 11268 2912 11299
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 8297 11339 8355 11345
rect 8297 11305 8309 11339
rect 8343 11336 8355 11339
rect 9490 11336 9496 11348
rect 8343 11308 9496 11336
rect 8343 11305 8355 11308
rect 8297 11299 8355 11305
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 10505 11339 10563 11345
rect 10505 11305 10517 11339
rect 10551 11336 10563 11339
rect 10870 11336 10876 11348
rect 10551 11308 10876 11336
rect 10551 11305 10563 11308
rect 10505 11299 10563 11305
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 19242 11296 19248 11348
rect 19300 11336 19306 11348
rect 19981 11339 20039 11345
rect 19981 11336 19993 11339
rect 19300 11308 19993 11336
rect 19300 11296 19306 11308
rect 19981 11305 19993 11308
rect 20027 11305 20039 11339
rect 22278 11336 22284 11348
rect 19981 11299 20039 11305
rect 22112 11308 22284 11336
rect 3418 11268 3424 11280
rect 2363 11240 2912 11268
rect 3379 11240 3424 11268
rect 2363 11237 2375 11240
rect 2317 11231 2375 11237
rect 3418 11228 3424 11240
rect 3476 11228 3482 11280
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 8757 11271 8815 11277
rect 8757 11268 8769 11271
rect 7892 11240 8769 11268
rect 7892 11228 7898 11240
rect 8757 11237 8769 11240
rect 8803 11237 8815 11271
rect 8757 11231 8815 11237
rect 15838 11228 15844 11280
rect 15896 11268 15902 11280
rect 16270 11271 16328 11277
rect 16270 11268 16282 11271
rect 15896 11240 16282 11268
rect 15896 11228 15902 11240
rect 16270 11237 16282 11240
rect 16316 11237 16328 11271
rect 16270 11231 16328 11237
rect 18690 11228 18696 11280
rect 18748 11268 18754 11280
rect 18868 11271 18926 11277
rect 18868 11268 18880 11271
rect 18748 11240 18880 11268
rect 18748 11228 18754 11240
rect 18868 11237 18880 11240
rect 18914 11268 18926 11271
rect 20806 11268 20812 11280
rect 18914 11240 20812 11268
rect 18914 11237 18926 11240
rect 18868 11231 18926 11237
rect 20806 11228 20812 11240
rect 20864 11228 20870 11280
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 5074 11200 5080 11212
rect 4663 11172 5080 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13061 11203 13119 11209
rect 13061 11200 13073 11203
rect 12952 11172 13073 11200
rect 12952 11160 12958 11172
rect 13061 11169 13073 11172
rect 13107 11169 13119 11203
rect 18598 11200 18604 11212
rect 18559 11172 18604 11200
rect 13061 11163 13119 11169
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 21542 11160 21548 11212
rect 21600 11200 21606 11212
rect 21913 11203 21971 11209
rect 21913 11200 21925 11203
rect 21600 11172 21925 11200
rect 21600 11160 21606 11172
rect 21913 11169 21925 11172
rect 21959 11200 21971 11203
rect 22112 11200 22140 11308
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 23290 11336 23296 11348
rect 23251 11308 23296 11336
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 23937 11339 23995 11345
rect 23937 11305 23949 11339
rect 23983 11336 23995 11339
rect 24302 11336 24308 11348
rect 23983 11308 24308 11336
rect 23983 11305 23995 11308
rect 23937 11299 23995 11305
rect 24302 11296 24308 11308
rect 24360 11296 24366 11348
rect 24394 11296 24400 11348
rect 24452 11336 24458 11348
rect 25314 11336 25320 11348
rect 24452 11308 24497 11336
rect 25227 11308 25320 11336
rect 24452 11296 24458 11308
rect 25314 11296 25320 11308
rect 25372 11336 25378 11348
rect 25774 11336 25780 11348
rect 25372 11308 25780 11336
rect 25372 11296 25378 11308
rect 25774 11296 25780 11308
rect 25832 11296 25838 11348
rect 26513 11339 26571 11345
rect 26513 11305 26525 11339
rect 26559 11305 26571 11339
rect 26970 11336 26976 11348
rect 26931 11308 26976 11336
rect 26513 11299 26571 11305
rect 22186 11277 22192 11280
rect 22180 11231 22192 11277
rect 22244 11268 22250 11280
rect 23014 11268 23020 11280
rect 22244 11240 23020 11268
rect 22186 11228 22192 11231
rect 22244 11228 22250 11240
rect 23014 11228 23020 11240
rect 23072 11228 23078 11280
rect 21959 11172 22140 11200
rect 24412 11200 24440 11296
rect 24854 11228 24860 11280
rect 24912 11268 24918 11280
rect 25038 11268 25044 11280
rect 24912 11240 25044 11268
rect 24912 11228 24918 11240
rect 25038 11228 25044 11240
rect 25096 11228 25102 11280
rect 25225 11271 25283 11277
rect 25225 11237 25237 11271
rect 25271 11268 25283 11271
rect 25498 11268 25504 11280
rect 25271 11240 25504 11268
rect 25271 11237 25283 11240
rect 25225 11231 25283 11237
rect 25498 11228 25504 11240
rect 25556 11268 25562 11280
rect 26528 11268 26556 11299
rect 26970 11296 26976 11308
rect 27028 11296 27034 11348
rect 26878 11268 26884 11280
rect 25556 11240 26556 11268
rect 26839 11240 26884 11268
rect 25556 11228 25562 11240
rect 26878 11228 26884 11240
rect 26936 11228 26942 11280
rect 25866 11200 25872 11212
rect 24412 11172 25872 11200
rect 21959 11169 21971 11172
rect 21913 11163 21971 11169
rect 25866 11160 25872 11172
rect 25924 11200 25930 11212
rect 27154 11200 27160 11212
rect 25924 11172 27160 11200
rect 25924 11160 25930 11172
rect 2590 11092 2596 11144
rect 2648 11132 2654 11144
rect 2774 11132 2780 11144
rect 2648 11104 2780 11132
rect 2648 11092 2654 11104
rect 2774 11092 2780 11104
rect 2832 11132 2838 11144
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2832 11104 2973 11132
rect 2832 11092 2838 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 5166 11132 5172 11144
rect 5127 11104 5172 11132
rect 2961 11095 3019 11101
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 10597 11135 10655 11141
rect 5316 11104 5361 11132
rect 5316 11092 5322 11104
rect 10597 11101 10609 11135
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 10962 11132 10968 11144
rect 10827 11104 10968 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 2314 11024 2320 11076
rect 2372 11064 2378 11076
rect 2409 11067 2467 11073
rect 2409 11064 2421 11067
rect 2372 11036 2421 11064
rect 2372 11024 2378 11036
rect 2409 11033 2421 11036
rect 2455 11033 2467 11067
rect 9950 11064 9956 11076
rect 9911 11036 9956 11064
rect 2409 11027 2467 11033
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 10612 11064 10640 11095
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12492 11104 12817 11132
rect 12492 11092 12498 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 16025 11135 16083 11141
rect 16025 11101 16037 11135
rect 16071 11101 16083 11135
rect 16025 11095 16083 11101
rect 10612 11036 11100 11064
rect 5718 10996 5724 11008
rect 5679 10968 5724 10996
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 10137 10999 10195 11005
rect 10137 10965 10149 10999
rect 10183 10996 10195 10999
rect 10318 10996 10324 11008
rect 10183 10968 10324 10996
rect 10183 10965 10195 10968
rect 10137 10959 10195 10965
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 11072 10996 11100 11036
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 14185 11067 14243 11073
rect 14185 11064 14197 11067
rect 13872 11036 14197 11064
rect 13872 11024 13878 11036
rect 14185 11033 14197 11036
rect 14231 11033 14243 11067
rect 14185 11027 14243 11033
rect 11330 10996 11336 11008
rect 11072 10968 11336 10996
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 16040 10996 16068 11095
rect 24946 11092 24952 11144
rect 25004 11132 25010 11144
rect 27080 11141 27108 11172
rect 27154 11160 27160 11172
rect 27212 11160 27218 11212
rect 25409 11135 25467 11141
rect 25409 11132 25421 11135
rect 25004 11104 25421 11132
rect 25004 11092 25010 11104
rect 25409 11101 25421 11104
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 27065 11135 27123 11141
rect 27065 11101 27077 11135
rect 27111 11101 27123 11135
rect 27065 11095 27123 11101
rect 17773 11067 17831 11073
rect 17773 11033 17785 11067
rect 17819 11064 17831 11067
rect 24854 11064 24860 11076
rect 17819 11036 17908 11064
rect 24815 11036 24860 11064
rect 17819 11033 17831 11036
rect 17773 11027 17831 11033
rect 17880 11008 17908 11036
rect 24854 11024 24860 11036
rect 24912 11024 24918 11076
rect 16942 10996 16948 11008
rect 16040 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 17405 10999 17463 11005
rect 17405 10996 17417 10999
rect 17092 10968 17417 10996
rect 17092 10956 17098 10968
rect 17405 10965 17417 10968
rect 17451 10965 17463 10999
rect 17862 10996 17868 11008
rect 17775 10968 17868 10996
rect 17405 10959 17463 10965
rect 17862 10956 17868 10968
rect 17920 10996 17926 11008
rect 19242 10996 19248 11008
rect 17920 10968 19248 10996
rect 17920 10956 17926 10968
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 1857 10795 1915 10801
rect 1857 10792 1869 10795
rect 1728 10764 1869 10792
rect 1728 10752 1734 10764
rect 1857 10761 1869 10764
rect 1903 10761 1915 10795
rect 1857 10755 1915 10761
rect 2409 10795 2467 10801
rect 2409 10761 2421 10795
rect 2455 10792 2467 10795
rect 2498 10792 2504 10804
rect 2455 10764 2504 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 1872 10656 1900 10755
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 4154 10792 4160 10804
rect 4115 10764 4160 10792
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4985 10795 5043 10801
rect 4985 10792 4997 10795
rect 4488 10764 4997 10792
rect 4488 10752 4494 10764
rect 4985 10761 4997 10764
rect 5031 10761 5043 10795
rect 4985 10755 5043 10761
rect 2317 10727 2375 10733
rect 2317 10693 2329 10727
rect 2363 10724 2375 10727
rect 2590 10724 2596 10736
rect 2363 10696 2596 10724
rect 2363 10693 2375 10696
rect 2317 10687 2375 10693
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 5000 10724 5028 10755
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 5132 10764 5181 10792
rect 5132 10752 5138 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 5169 10755 5227 10761
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11425 10795 11483 10801
rect 11425 10792 11437 10795
rect 11112 10764 11437 10792
rect 11112 10752 11118 10764
rect 11425 10761 11437 10764
rect 11471 10761 11483 10795
rect 11425 10755 11483 10761
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12342 10792 12348 10804
rect 12299 10764 12348 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12894 10792 12900 10804
rect 12855 10764 12900 10792
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15896 10764 16037 10792
rect 15896 10752 15902 10764
rect 16025 10761 16037 10764
rect 16071 10761 16083 10795
rect 16025 10755 16083 10761
rect 18598 10752 18604 10804
rect 18656 10792 18662 10804
rect 18969 10795 19027 10801
rect 18969 10792 18981 10795
rect 18656 10764 18981 10792
rect 18656 10752 18662 10764
rect 18969 10761 18981 10764
rect 19015 10761 19027 10795
rect 22002 10792 22008 10804
rect 21963 10764 22008 10792
rect 18969 10755 19027 10761
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 22278 10792 22284 10804
rect 22239 10764 22284 10792
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 23474 10792 23480 10804
rect 23435 10764 23480 10792
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 24946 10792 24952 10804
rect 24907 10764 24952 10792
rect 24946 10752 24952 10764
rect 25004 10752 25010 10804
rect 25314 10792 25320 10804
rect 25275 10764 25320 10792
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 25866 10792 25872 10804
rect 25827 10764 25872 10792
rect 25866 10752 25872 10764
rect 25924 10752 25930 10804
rect 26329 10795 26387 10801
rect 26329 10761 26341 10795
rect 26375 10792 26387 10795
rect 26878 10792 26884 10804
rect 26375 10764 26884 10792
rect 26375 10761 26387 10764
rect 26329 10755 26387 10761
rect 26878 10752 26884 10764
rect 26936 10752 26942 10804
rect 26970 10752 26976 10804
rect 27028 10792 27034 10804
rect 27341 10795 27399 10801
rect 27341 10792 27353 10795
rect 27028 10764 27353 10792
rect 27028 10752 27034 10764
rect 27341 10761 27353 10764
rect 27387 10761 27399 10795
rect 27341 10755 27399 10761
rect 5000 10696 5396 10724
rect 3053 10659 3111 10665
rect 3053 10656 3065 10659
rect 1872 10628 3065 10656
rect 3053 10625 3065 10628
rect 3099 10656 3111 10659
rect 5258 10656 5264 10668
rect 3099 10628 5264 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4614 10588 4620 10600
rect 4019 10560 4620 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 2869 10523 2927 10529
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 3050 10520 3056 10532
rect 2915 10492 3056 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 3050 10480 3056 10492
rect 3108 10520 3114 10532
rect 3421 10523 3479 10529
rect 3421 10520 3433 10523
rect 3108 10492 3433 10520
rect 3108 10480 3114 10492
rect 3421 10489 3433 10492
rect 3467 10489 3479 10523
rect 3421 10483 3479 10489
rect 3881 10523 3939 10529
rect 3881 10489 3893 10523
rect 3927 10520 3939 10523
rect 5166 10520 5172 10532
rect 3927 10492 5172 10520
rect 3927 10489 3939 10492
rect 3881 10483 3939 10489
rect 5166 10480 5172 10492
rect 5224 10480 5230 10532
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 5368 10452 5396 10696
rect 14366 10684 14372 10736
rect 14424 10724 14430 10736
rect 14921 10727 14979 10733
rect 14921 10724 14933 10727
rect 14424 10696 14933 10724
rect 14424 10684 14430 10696
rect 14921 10693 14933 10696
rect 14967 10693 14979 10727
rect 17494 10724 17500 10736
rect 14921 10687 14979 10693
rect 15028 10696 17500 10724
rect 5718 10656 5724 10668
rect 5679 10628 5724 10656
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10656 9275 10659
rect 9582 10656 9588 10668
rect 9263 10628 9588 10656
rect 9263 10625 9275 10628
rect 9217 10619 9275 10625
rect 9582 10616 9588 10628
rect 9640 10656 9646 10668
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 9640 10628 10701 10656
rect 9640 10616 9646 10628
rect 10689 10625 10701 10628
rect 10735 10656 10747 10659
rect 10778 10656 10784 10668
rect 10735 10628 10784 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 10778 10616 10784 10628
rect 10836 10656 10842 10668
rect 10962 10656 10968 10668
rect 10836 10628 10968 10656
rect 10836 10616 10842 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11241 10659 11299 10665
rect 11241 10625 11253 10659
rect 11287 10656 11299 10659
rect 15028 10656 15056 10696
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 18690 10724 18696 10736
rect 18651 10696 18696 10724
rect 18690 10684 18696 10696
rect 18748 10684 18754 10736
rect 23492 10724 23520 10752
rect 26602 10724 26608 10736
rect 23492 10696 24256 10724
rect 26563 10696 26608 10724
rect 11287 10628 15056 10656
rect 15749 10659 15807 10665
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 16390 10656 16396 10668
rect 15795 10628 16396 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 16390 10616 16396 10628
rect 16448 10656 16454 10668
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16448 10628 16865 10656
rect 16448 10616 16454 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 17034 10656 17040 10668
rect 16995 10628 17040 10656
rect 16853 10619 16911 10625
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 18598 10616 18604 10668
rect 18656 10656 18662 10668
rect 18782 10656 18788 10668
rect 18656 10628 18788 10656
rect 18656 10616 18662 10628
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 23842 10616 23848 10668
rect 23900 10656 23906 10668
rect 24228 10665 24256 10696
rect 26602 10684 26608 10696
rect 26660 10684 26666 10736
rect 24121 10659 24179 10665
rect 24121 10656 24133 10659
rect 23900 10628 24133 10656
rect 23900 10616 23906 10628
rect 24121 10625 24133 10628
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 24213 10659 24271 10665
rect 24213 10625 24225 10659
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5592 10560 5641 10588
rect 5592 10548 5598 10560
rect 5629 10557 5641 10560
rect 5675 10588 5687 10591
rect 5810 10588 5816 10600
rect 5675 10560 5816 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 5810 10548 5816 10560
rect 5868 10588 5874 10600
rect 6181 10591 6239 10597
rect 6181 10588 6193 10591
rect 5868 10560 6193 10588
rect 5868 10548 5874 10560
rect 6181 10557 6193 10560
rect 6227 10557 6239 10591
rect 6181 10551 6239 10557
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10588 10011 10591
rect 10410 10588 10416 10600
rect 9999 10560 10416 10588
rect 9999 10557 10011 10560
rect 9953 10551 10011 10557
rect 10410 10548 10416 10560
rect 10468 10548 10474 10600
rect 16574 10588 16580 10600
rect 10520 10560 16580 10588
rect 10520 10529 10548 10560
rect 16574 10548 16580 10560
rect 16632 10548 16638 10600
rect 16761 10591 16819 10597
rect 16761 10557 16773 10591
rect 16807 10588 16819 10591
rect 17126 10588 17132 10600
rect 16807 10560 17132 10588
rect 16807 10557 16819 10560
rect 16761 10551 16819 10557
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 23109 10591 23167 10597
rect 23109 10557 23121 10591
rect 23155 10588 23167 10591
rect 24029 10591 24087 10597
rect 24029 10588 24041 10591
rect 23155 10560 24041 10588
rect 23155 10557 23167 10560
rect 23109 10551 23167 10557
rect 24029 10557 24041 10560
rect 24075 10588 24087 10591
rect 24762 10588 24768 10600
rect 24075 10560 24768 10588
rect 24075 10557 24087 10560
rect 24029 10551 24087 10557
rect 24762 10548 24768 10560
rect 24820 10548 24826 10600
rect 26418 10588 26424 10600
rect 26379 10560 26424 10588
rect 26418 10548 26424 10560
rect 26476 10588 26482 10600
rect 26973 10591 27031 10597
rect 26973 10588 26985 10591
rect 26476 10560 26985 10588
rect 26476 10548 26482 10560
rect 26973 10557 26985 10560
rect 27019 10557 27031 10591
rect 26973 10551 27031 10557
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 9508 10492 10517 10520
rect 9508 10464 9536 10492
rect 10505 10489 10517 10492
rect 10551 10489 10563 10523
rect 11241 10523 11299 10529
rect 11241 10520 11253 10523
rect 10505 10483 10563 10489
rect 11072 10492 11253 10520
rect 5534 10452 5540 10464
rect 2832 10424 2877 10452
rect 5368 10424 5540 10452
rect 2832 10412 2838 10424
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 9490 10452 9496 10464
rect 9451 10424 9496 10452
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10410 10452 10416 10464
rect 10323 10424 10416 10452
rect 10410 10412 10416 10424
rect 10468 10452 10474 10464
rect 11072 10452 11100 10492
rect 11241 10489 11253 10492
rect 11287 10489 11299 10523
rect 11241 10483 11299 10489
rect 13633 10523 13691 10529
rect 13633 10489 13645 10523
rect 13679 10489 13691 10523
rect 13633 10483 13691 10489
rect 10468 10424 11100 10452
rect 11149 10455 11207 10461
rect 10468 10412 10474 10424
rect 11149 10421 11161 10455
rect 11195 10452 11207 10455
rect 11330 10452 11336 10464
rect 11195 10424 11336 10452
rect 11195 10421 11207 10424
rect 11149 10415 11207 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 13446 10452 13452 10464
rect 13407 10424 13452 10452
rect 13446 10412 13452 10424
rect 13504 10452 13510 10464
rect 13648 10452 13676 10483
rect 16390 10452 16396 10464
rect 13504 10424 13676 10452
rect 16351 10424 16396 10452
rect 13504 10412 13510 10424
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 17402 10452 17408 10464
rect 17000 10424 17408 10452
rect 17000 10412 17006 10424
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 23658 10452 23664 10464
rect 23619 10424 23664 10452
rect 23658 10412 23664 10424
rect 23716 10412 23722 10464
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2774 10248 2780 10260
rect 2363 10220 2780 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 4985 10251 5043 10257
rect 4985 10217 4997 10251
rect 5031 10248 5043 10251
rect 5166 10248 5172 10260
rect 5031 10220 5172 10248
rect 5031 10217 5043 10220
rect 4985 10211 5043 10217
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 5353 10251 5411 10257
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 6638 10248 6644 10260
rect 5399 10220 6644 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 4801 10183 4859 10189
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 5258 10180 5264 10192
rect 4847 10152 5264 10180
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 5258 10140 5264 10152
rect 5316 10140 5322 10192
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 3234 10112 3240 10124
rect 2823 10084 3240 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5368 10112 5396 10211
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 6880 10220 6929 10248
rect 6880 10208 6886 10220
rect 6917 10217 6929 10220
rect 6963 10248 6975 10251
rect 7190 10248 7196 10260
rect 6963 10220 7196 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10413 10251 10471 10257
rect 10413 10248 10425 10251
rect 10100 10220 10425 10248
rect 10100 10208 10106 10220
rect 10413 10217 10425 10220
rect 10459 10217 10471 10251
rect 10413 10211 10471 10217
rect 12621 10251 12679 10257
rect 12621 10217 12633 10251
rect 12667 10248 12679 10251
rect 13081 10251 13139 10257
rect 13081 10248 13093 10251
rect 12667 10220 13093 10248
rect 12667 10217 12679 10220
rect 12621 10211 12679 10217
rect 13081 10217 13093 10220
rect 13127 10248 13139 10251
rect 15289 10251 15347 10257
rect 15289 10248 15301 10251
rect 13127 10220 15301 10248
rect 13127 10217 13139 10220
rect 13081 10211 13139 10217
rect 15289 10217 15301 10220
rect 15335 10217 15347 10251
rect 15289 10211 15347 10217
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 15749 10251 15807 10257
rect 15749 10248 15761 10251
rect 15436 10220 15761 10248
rect 15436 10208 15442 10220
rect 15749 10217 15761 10220
rect 15795 10217 15807 10251
rect 15749 10211 15807 10217
rect 16853 10251 16911 10257
rect 16853 10217 16865 10251
rect 16899 10248 16911 10251
rect 17126 10248 17132 10260
rect 16899 10220 17132 10248
rect 16899 10217 16911 10220
rect 16853 10211 16911 10217
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 19337 10251 19395 10257
rect 19337 10217 19349 10251
rect 19383 10248 19395 10251
rect 19518 10248 19524 10260
rect 19383 10220 19524 10248
rect 19383 10217 19395 10220
rect 19337 10211 19395 10217
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 23017 10251 23075 10257
rect 23017 10248 23029 10251
rect 21876 10220 23029 10248
rect 21876 10208 21882 10220
rect 23017 10217 23029 10220
rect 23063 10217 23075 10251
rect 23017 10211 23075 10217
rect 23753 10251 23811 10257
rect 23753 10217 23765 10251
rect 23799 10248 23811 10251
rect 23842 10248 23848 10260
rect 23799 10220 23848 10248
rect 23799 10217 23811 10220
rect 23753 10211 23811 10217
rect 23842 10208 23848 10220
rect 23900 10208 23906 10260
rect 25498 10248 25504 10260
rect 25459 10220 25504 10248
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 26694 10248 26700 10260
rect 26655 10220 26700 10248
rect 26694 10208 26700 10220
rect 26752 10208 26758 10260
rect 10318 10180 10324 10192
rect 10279 10152 10324 10180
rect 10318 10140 10324 10152
rect 10376 10140 10382 10192
rect 13906 10180 13912 10192
rect 13867 10152 13912 10180
rect 13906 10140 13912 10152
rect 13964 10180 13970 10192
rect 14274 10180 14280 10192
rect 13964 10152 14280 10180
rect 13964 10140 13970 10152
rect 14274 10140 14280 10152
rect 14332 10140 14338 10192
rect 16485 10183 16543 10189
rect 16485 10149 16497 10183
rect 16531 10180 16543 10183
rect 17034 10180 17040 10192
rect 16531 10152 17040 10180
rect 16531 10149 16543 10152
rect 16485 10143 16543 10149
rect 5132 10084 5396 10112
rect 5132 10072 5138 10084
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 11057 10115 11115 10121
rect 11057 10112 11069 10115
rect 10836 10084 11069 10112
rect 10836 10072 10842 10084
rect 11057 10081 11069 10084
rect 11103 10112 11115 10115
rect 12710 10112 12716 10124
rect 11103 10084 12716 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 12710 10072 12716 10084
rect 12768 10112 12774 10124
rect 15654 10112 15660 10124
rect 12768 10084 13400 10112
rect 15615 10084 15660 10112
rect 12768 10072 12774 10084
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3326 10044 3332 10056
rect 3007 10016 3332 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3326 10004 3332 10016
rect 3384 10044 3390 10056
rect 5445 10047 5503 10053
rect 3384 10016 3464 10044
rect 3384 10004 3390 10016
rect 2409 9979 2467 9985
rect 2409 9945 2421 9979
rect 2455 9976 2467 9979
rect 3050 9976 3056 9988
rect 2455 9948 3056 9976
rect 2455 9945 2467 9948
rect 2409 9939 2467 9945
rect 3050 9936 3056 9948
rect 3108 9936 3114 9988
rect 3436 9920 3464 10016
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5626 10044 5632 10056
rect 5587 10016 5632 10044
rect 5445 10007 5503 10013
rect 1670 9908 1676 9920
rect 1631 9880 1676 9908
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 3418 9908 3424 9920
rect 3379 9880 3424 9908
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 5460 9908 5488 10007
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 7006 10044 7012 10056
rect 6967 10016 7012 10044
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7098 10004 7104 10056
rect 7156 10044 7162 10056
rect 10594 10044 10600 10056
rect 7156 10016 7201 10044
rect 10555 10016 10600 10044
rect 7156 10004 7162 10016
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 13170 10044 13176 10056
rect 13131 10016 13176 10044
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13372 10053 13400 10084
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 15746 10072 15752 10124
rect 15804 10112 15810 10124
rect 16500 10112 16528 10143
rect 17034 10140 17040 10152
rect 17092 10140 17098 10192
rect 24765 10183 24823 10189
rect 24765 10149 24777 10183
rect 24811 10180 24823 10183
rect 24946 10180 24952 10192
rect 24811 10152 24952 10180
rect 24811 10149 24823 10152
rect 24765 10143 24823 10149
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 15804 10084 16528 10112
rect 15804 10072 15810 10084
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18322 10112 18328 10124
rect 18104 10084 18328 10112
rect 18104 10072 18110 10084
rect 18322 10072 18328 10084
rect 18380 10112 18386 10124
rect 21910 10121 21916 10124
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 18380 10084 18613 10112
rect 18380 10072 18386 10084
rect 18601 10081 18613 10084
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 21904 10075 21916 10121
rect 21968 10112 21974 10124
rect 21968 10084 22004 10112
rect 21910 10072 21916 10075
rect 21968 10072 21974 10084
rect 25590 10072 25596 10124
rect 25648 10112 25654 10124
rect 26513 10115 26571 10121
rect 26513 10112 26525 10115
rect 25648 10084 26525 10112
rect 25648 10072 25654 10084
rect 26513 10081 26525 10084
rect 26559 10112 26571 10115
rect 27338 10112 27344 10124
rect 26559 10084 27344 10112
rect 26559 10081 26571 10084
rect 26513 10075 26571 10081
rect 27338 10072 27344 10084
rect 27396 10072 27402 10124
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10044 13415 10047
rect 13722 10044 13728 10056
rect 13403 10016 13728 10044
rect 13403 10013 13415 10016
rect 13357 10007 13415 10013
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 13998 10044 14004 10056
rect 13959 10016 14004 10044
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 14090 10004 14096 10056
rect 14148 10044 14154 10056
rect 15838 10044 15844 10056
rect 14148 10016 14193 10044
rect 15799 10016 15844 10044
rect 14148 10004 14154 10016
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 18690 10044 18696 10056
rect 18651 10016 18696 10044
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 18877 10047 18935 10053
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 19242 10044 19248 10056
rect 18923 10016 19248 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 21634 10044 21640 10056
rect 21595 10016 21640 10044
rect 21634 10004 21640 10016
rect 21692 10004 21698 10056
rect 24854 10044 24860 10056
rect 24815 10016 24860 10044
rect 24854 10004 24860 10016
rect 24912 10004 24918 10056
rect 25038 10044 25044 10056
rect 24999 10016 25044 10044
rect 25038 10004 25044 10016
rect 25096 10004 25102 10056
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 11330 9976 11336 9988
rect 9999 9948 11336 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 11330 9936 11336 9948
rect 11388 9936 11394 9988
rect 13188 9976 13216 10004
rect 13541 9979 13599 9985
rect 13541 9976 13553 9979
rect 13188 9948 13553 9976
rect 13541 9945 13553 9948
rect 13587 9945 13599 9979
rect 14642 9976 14648 9988
rect 14603 9948 14648 9976
rect 13541 9939 13599 9945
rect 14642 9936 14648 9948
rect 14700 9936 14706 9988
rect 5810 9908 5816 9920
rect 5460 9880 5816 9908
rect 5810 9868 5816 9880
rect 5868 9908 5874 9920
rect 6549 9911 6607 9917
rect 6549 9908 6561 9911
rect 5868 9880 6561 9908
rect 5868 9868 5874 9880
rect 6549 9877 6561 9880
rect 6595 9877 6607 9911
rect 9306 9908 9312 9920
rect 9267 9880 9312 9908
rect 6549 9871 6607 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 12253 9911 12311 9917
rect 12253 9877 12265 9911
rect 12299 9908 12311 9911
rect 12342 9908 12348 9920
rect 12299 9880 12348 9908
rect 12299 9877 12311 9880
rect 12253 9871 12311 9877
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 12713 9911 12771 9917
rect 12713 9877 12725 9911
rect 12759 9908 12771 9911
rect 12894 9908 12900 9920
rect 12759 9880 12900 9908
rect 12759 9877 12771 9880
rect 12713 9871 12771 9877
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18233 9911 18291 9917
rect 18233 9908 18245 9911
rect 18012 9880 18245 9908
rect 18012 9868 18018 9880
rect 18233 9877 18245 9880
rect 18279 9877 18291 9911
rect 18233 9871 18291 9877
rect 23474 9868 23480 9920
rect 23532 9908 23538 9920
rect 24397 9911 24455 9917
rect 24397 9908 24409 9911
rect 23532 9880 24409 9908
rect 23532 9868 23538 9880
rect 24397 9877 24409 9880
rect 24443 9877 24455 9911
rect 24397 9871 24455 9877
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 3234 9704 3240 9716
rect 2832 9676 2877 9704
rect 2976 9676 3240 9704
rect 2832 9664 2838 9676
rect 2501 9639 2559 9645
rect 2501 9605 2513 9639
rect 2547 9636 2559 9639
rect 2976 9636 3004 9676
rect 3234 9664 3240 9676
rect 3292 9664 3298 9716
rect 5074 9704 5080 9716
rect 4816 9676 5080 9704
rect 2547 9608 3004 9636
rect 2547 9605 2559 9608
rect 2501 9599 2559 9605
rect 2130 9568 2136 9580
rect 2043 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9568 2194 9580
rect 3234 9568 3240 9580
rect 2188 9540 3240 9568
rect 2188 9528 2194 9540
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3418 9568 3424 9580
rect 3331 9540 3424 9568
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 4816 9568 4844 9676
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 5810 9704 5816 9716
rect 5771 9676 5816 9704
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 10318 9664 10324 9716
rect 10376 9704 10382 9716
rect 10965 9707 11023 9713
rect 10965 9704 10977 9707
rect 10376 9676 10977 9704
rect 10376 9664 10382 9676
rect 10965 9673 10977 9676
rect 11011 9673 11023 9707
rect 10965 9667 11023 9673
rect 11885 9707 11943 9713
rect 11885 9673 11897 9707
rect 11931 9704 11943 9707
rect 13170 9704 13176 9716
rect 11931 9676 13176 9704
rect 11931 9673 11943 9676
rect 11885 9667 11943 9673
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 13998 9704 14004 9716
rect 13832 9676 14004 9704
rect 5718 9596 5724 9648
rect 5776 9636 5782 9648
rect 6273 9639 6331 9645
rect 6273 9636 6285 9639
rect 5776 9608 6285 9636
rect 5776 9596 5782 9608
rect 6273 9605 6285 9608
rect 6319 9636 6331 9639
rect 6822 9636 6828 9648
rect 6319 9608 6828 9636
rect 6319 9605 6331 9608
rect 6273 9599 6331 9605
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 5166 9568 5172 9580
rect 4816 9540 5172 9568
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12544 9540 13001 9568
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1670 9500 1676 9512
rect 1443 9472 1676 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 3436 9500 3464 9528
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 3436 9472 4261 9500
rect 4249 9469 4261 9472
rect 4295 9500 4307 9503
rect 4295 9472 5488 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 5460 9441 5488 9472
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6696 9472 6837 9500
rect 6696 9460 6702 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 9214 9500 9220 9512
rect 9175 9472 9220 9500
rect 6825 9463 6883 9469
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9306 9460 9312 9512
rect 9364 9500 9370 9512
rect 9582 9509 9588 9512
rect 9576 9500 9588 9509
rect 9364 9472 9409 9500
rect 9508 9472 9588 9500
rect 9364 9460 9370 9472
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3881 9435 3939 9441
rect 3881 9432 3893 9435
rect 3191 9404 3893 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 3881 9401 3893 9404
rect 3927 9432 3939 9435
rect 4341 9435 4399 9441
rect 4341 9432 4353 9435
rect 3927 9404 4353 9432
rect 3927 9401 3939 9404
rect 3881 9395 3939 9401
rect 4341 9401 4353 9404
rect 4387 9401 4399 9435
rect 4341 9395 4399 9401
rect 5445 9435 5503 9441
rect 5445 9401 5457 9435
rect 5491 9432 5503 9435
rect 5626 9432 5632 9444
rect 5491 9404 5632 9432
rect 5491 9401 5503 9404
rect 5445 9395 5503 9401
rect 5626 9392 5632 9404
rect 5684 9432 5690 9444
rect 5684 9404 6960 9432
rect 5684 9392 5690 9404
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5166 9364 5172 9376
rect 5123 9336 5172 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6420 9336 6561 9364
rect 6420 9324 6426 9336
rect 6549 9333 6561 9336
rect 6595 9364 6607 9367
rect 6822 9364 6828 9376
rect 6595 9336 6828 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 6932 9364 6960 9404
rect 7006 9392 7012 9444
rect 7064 9441 7070 9444
rect 7064 9435 7128 9441
rect 7064 9401 7082 9435
rect 7116 9401 7128 9435
rect 7064 9395 7128 9401
rect 8941 9435 8999 9441
rect 8941 9401 8953 9435
rect 8987 9432 8999 9435
rect 9508 9432 9536 9472
rect 9576 9463 9588 9472
rect 9582 9460 9588 9463
rect 9640 9460 9646 9512
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 11514 9500 11520 9512
rect 10744 9472 11520 9500
rect 10744 9460 10750 9472
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12544 9500 12572 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 12894 9500 12900 9512
rect 12299 9472 12572 9500
rect 12855 9472 12900 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 8987 9404 9536 9432
rect 8987 9401 8999 9404
rect 8941 9395 8999 9401
rect 7064 9392 7070 9395
rect 10594 9392 10600 9444
rect 10652 9432 10658 9444
rect 12268 9432 12296 9463
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 13832 9500 13860 9676
rect 13998 9664 14004 9676
rect 14056 9704 14062 9716
rect 18598 9704 18604 9716
rect 14056 9676 18604 9704
rect 14056 9664 14062 9676
rect 18598 9664 18604 9676
rect 18656 9664 18662 9716
rect 21634 9704 21640 9716
rect 20640 9676 21640 9704
rect 15378 9636 15384 9648
rect 15339 9608 15384 9636
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 17862 9636 17868 9648
rect 17823 9608 17868 9636
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 18322 9636 18328 9648
rect 18283 9608 18328 9636
rect 18322 9596 18328 9608
rect 18380 9596 18386 9648
rect 18782 9596 18788 9648
rect 18840 9636 18846 9648
rect 19702 9636 19708 9648
rect 18840 9608 19708 9636
rect 18840 9596 18846 9608
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 14553 9571 14611 9577
rect 14553 9568 14565 9571
rect 14148 9540 14565 9568
rect 14148 9528 14154 9540
rect 14553 9537 14565 9540
rect 14599 9568 14611 9571
rect 14734 9568 14740 9580
rect 14599 9540 14740 9568
rect 14599 9537 14611 9540
rect 14553 9531 14611 9537
rect 14734 9528 14740 9540
rect 14792 9568 14798 9580
rect 15838 9568 15844 9580
rect 14792 9540 15844 9568
rect 14792 9528 14798 9540
rect 15838 9528 15844 9540
rect 15896 9568 15902 9580
rect 19628 9577 19656 9608
rect 19702 9596 19708 9608
rect 19760 9636 19766 9648
rect 20073 9639 20131 9645
rect 20073 9636 20085 9639
rect 19760 9608 20085 9636
rect 19760 9596 19766 9608
rect 20073 9605 20085 9608
rect 20119 9605 20131 9639
rect 20073 9599 20131 9605
rect 20530 9596 20536 9648
rect 20588 9636 20594 9648
rect 20640 9636 20668 9676
rect 21634 9664 21640 9676
rect 21692 9664 21698 9716
rect 21729 9707 21787 9713
rect 21729 9673 21741 9707
rect 21775 9704 21787 9707
rect 21910 9704 21916 9716
rect 21775 9676 21916 9704
rect 21775 9673 21787 9676
rect 21729 9667 21787 9673
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 22005 9707 22063 9713
rect 22005 9673 22017 9707
rect 22051 9704 22063 9707
rect 22051 9676 22085 9704
rect 22051 9673 22063 9676
rect 22005 9667 22063 9673
rect 20588 9608 20668 9636
rect 20588 9596 20594 9608
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15896 9540 16037 9568
rect 15896 9528 15902 9540
rect 16025 9537 16037 9540
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9568 19671 9571
rect 19659 9540 19693 9568
rect 19659 9537 19671 9540
rect 19613 9531 19671 9537
rect 21358 9528 21364 9580
rect 21416 9568 21422 9580
rect 21450 9568 21456 9580
rect 21416 9540 21456 9568
rect 21416 9528 21422 9540
rect 21450 9528 21456 9540
rect 21508 9528 21514 9580
rect 21652 9568 21680 9664
rect 22020 9568 22048 9667
rect 23198 9664 23204 9716
rect 23256 9704 23262 9716
rect 25406 9704 25412 9716
rect 23256 9676 25412 9704
rect 23256 9664 23262 9676
rect 25406 9664 25412 9676
rect 25464 9664 25470 9716
rect 27338 9704 27344 9716
rect 27299 9676 27344 9704
rect 27338 9664 27344 9676
rect 27396 9664 27402 9716
rect 24854 9596 24860 9648
rect 24912 9636 24918 9648
rect 25317 9639 25375 9645
rect 25317 9636 25329 9639
rect 24912 9608 25329 9636
rect 24912 9596 24918 9608
rect 25317 9605 25329 9608
rect 25363 9605 25375 9639
rect 26602 9636 26608 9648
rect 26563 9608 26608 9636
rect 25317 9599 25375 9605
rect 26602 9596 26608 9608
rect 26660 9596 26666 9648
rect 21652 9540 23704 9568
rect 13556 9472 13860 9500
rect 14369 9503 14427 9509
rect 10652 9404 12296 9432
rect 10652 9392 10658 9404
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 6932 9336 8217 9364
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 8205 9327 8263 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 10704 9373 10732 9404
rect 10689 9367 10747 9373
rect 10689 9333 10701 9367
rect 10735 9333 10747 9367
rect 10689 9327 10747 9333
rect 12250 9324 12256 9376
rect 12308 9364 12314 9376
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 12308 9336 12449 9364
rect 12308 9324 12314 9336
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12802 9364 12808 9376
rect 12763 9336 12808 9364
rect 12437 9327 12495 9333
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 13556 9373 13584 9472
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 14642 9500 14648 9512
rect 14415 9472 14648 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 18874 9460 18880 9512
rect 18932 9500 18938 9512
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 18932 9472 18981 9500
rect 18932 9460 18938 9472
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 19518 9500 19524 9512
rect 19475 9472 19524 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 23676 9509 23704 9540
rect 24946 9528 24952 9580
rect 25004 9568 25010 9580
rect 25406 9568 25412 9580
rect 25004 9540 25412 9568
rect 25004 9528 25010 9540
rect 25406 9528 25412 9540
rect 25464 9568 25470 9580
rect 25685 9571 25743 9577
rect 25685 9568 25697 9571
rect 25464 9540 25697 9568
rect 25464 9528 25470 9540
rect 25685 9537 25697 9540
rect 25731 9537 25743 9571
rect 25685 9531 25743 9537
rect 23477 9503 23535 9509
rect 23477 9469 23489 9503
rect 23523 9500 23535 9503
rect 23661 9503 23719 9509
rect 23523 9472 23612 9500
rect 23523 9469 23535 9472
rect 23477 9463 23535 9469
rect 23584 9444 23612 9472
rect 23661 9469 23673 9503
rect 23707 9500 23719 9503
rect 23750 9500 23756 9512
rect 23707 9472 23756 9500
rect 23707 9469 23719 9472
rect 23661 9463 23719 9469
rect 23750 9460 23756 9472
rect 23808 9460 23814 9512
rect 26326 9460 26332 9512
rect 26384 9500 26390 9512
rect 26421 9503 26479 9509
rect 26421 9500 26433 9503
rect 26384 9472 26433 9500
rect 26384 9460 26390 9472
rect 26421 9469 26433 9472
rect 26467 9500 26479 9503
rect 26973 9503 27031 9509
rect 26973 9500 26985 9503
rect 26467 9472 26985 9500
rect 26467 9469 26479 9472
rect 26421 9463 26479 9469
rect 26973 9469 26985 9472
rect 27019 9469 27031 9503
rect 26973 9463 27031 9469
rect 18693 9435 18751 9441
rect 18693 9401 18705 9435
rect 18739 9432 18751 9435
rect 19150 9432 19156 9444
rect 18739 9404 19156 9432
rect 18739 9401 18751 9404
rect 18693 9395 18751 9401
rect 19150 9392 19156 9404
rect 19208 9432 19214 9444
rect 19208 9404 19564 9432
rect 19208 9392 19214 9404
rect 19536 9376 19564 9404
rect 21910 9392 21916 9444
rect 21968 9432 21974 9444
rect 22094 9432 22100 9444
rect 21968 9404 22100 9432
rect 21968 9392 21974 9404
rect 22094 9392 22100 9404
rect 22152 9432 22158 9444
rect 22152 9404 23520 9432
rect 22152 9392 22158 9404
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 13044 9336 13553 9364
rect 13044 9324 13050 9336
rect 13541 9333 13553 9336
rect 13587 9333 13599 9367
rect 13998 9364 14004 9376
rect 13959 9336 14004 9364
rect 13541 9327 13599 9333
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14240 9336 14473 9364
rect 14240 9324 14246 9336
rect 14461 9333 14473 9336
rect 14507 9333 14519 9367
rect 15654 9364 15660 9376
rect 15615 9336 15660 9364
rect 14461 9327 14519 9333
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 18782 9364 18788 9376
rect 18743 9336 18788 9364
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 19058 9364 19064 9376
rect 19019 9336 19064 9364
rect 19058 9324 19064 9336
rect 19116 9324 19122 9376
rect 19518 9364 19524 9376
rect 19479 9336 19524 9364
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 23492 9364 23520 9404
rect 23566 9392 23572 9444
rect 23624 9432 23630 9444
rect 23928 9435 23986 9441
rect 23928 9432 23940 9435
rect 23624 9404 23940 9432
rect 23624 9392 23630 9404
rect 23928 9401 23940 9404
rect 23974 9432 23986 9435
rect 25498 9432 25504 9444
rect 23974 9404 25504 9432
rect 23974 9401 23986 9404
rect 23928 9395 23986 9401
rect 25498 9392 25504 9404
rect 25556 9392 25562 9444
rect 25038 9364 25044 9376
rect 23492 9336 25044 9364
rect 25038 9324 25044 9336
rect 25096 9324 25102 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 2682 9160 2688 9172
rect 2643 9132 2688 9160
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9214 9160 9220 9172
rect 9171 9132 9220 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10321 9163 10379 9169
rect 10321 9160 10333 9163
rect 10100 9132 10333 9160
rect 10100 9120 10106 9132
rect 10321 9129 10333 9132
rect 10367 9129 10379 9163
rect 10321 9123 10379 9129
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 11698 9160 11704 9172
rect 11388 9132 11704 9160
rect 11388 9120 11394 9132
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 12437 9163 12495 9169
rect 12437 9129 12449 9163
rect 12483 9160 12495 9163
rect 12894 9160 12900 9172
rect 12483 9132 12900 9160
rect 12483 9129 12495 9132
rect 12437 9123 12495 9129
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 13354 9160 13360 9172
rect 13267 9132 13360 9160
rect 13354 9120 13360 9132
rect 13412 9160 13418 9172
rect 13998 9160 14004 9172
rect 13412 9132 14004 9160
rect 13412 9120 13418 9132
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14734 9160 14740 9172
rect 14695 9132 14740 9160
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 15746 9160 15752 9172
rect 15707 9132 15752 9160
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 16301 9163 16359 9169
rect 16301 9129 16313 9163
rect 16347 9160 16359 9163
rect 16390 9160 16396 9172
rect 16347 9132 16396 9160
rect 16347 9129 16359 9132
rect 16301 9123 16359 9129
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 18601 9163 18659 9169
rect 18601 9129 18613 9163
rect 18647 9160 18659 9163
rect 18690 9160 18696 9172
rect 18647 9132 18696 9160
rect 18647 9129 18659 9132
rect 18601 9123 18659 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 18874 9160 18880 9172
rect 18835 9132 18880 9160
rect 18874 9120 18880 9132
rect 18932 9120 18938 9172
rect 24854 9160 24860 9172
rect 24815 9132 24860 9160
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 25222 9160 25228 9172
rect 25183 9132 25228 9160
rect 25222 9120 25228 9132
rect 25280 9120 25286 9172
rect 25314 9120 25320 9172
rect 25372 9160 25378 9172
rect 26694 9160 26700 9172
rect 25372 9132 25417 9160
rect 26655 9132 26700 9160
rect 25372 9120 25378 9132
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 12710 9092 12716 9104
rect 10744 9064 12572 9092
rect 12671 9064 12716 9092
rect 10744 9052 10750 9064
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1670 9024 1676 9036
rect 1443 8996 1676 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1670 8984 1676 8996
rect 1728 9024 1734 9036
rect 2130 9024 2136 9036
rect 1728 8996 2136 9024
rect 1728 8984 1734 8996
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 2498 9024 2504 9036
rect 2459 8996 2504 9024
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10594 9024 10600 9036
rect 10091 8996 10600 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 12250 9024 12256 9036
rect 11808 8996 12256 9024
rect 4062 8956 4068 8968
rect 4023 8928 4068 8956
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 6696 8928 7297 8956
rect 6696 8916 6702 8928
rect 7285 8925 7297 8928
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 11422 8916 11428 8968
rect 11480 8956 11486 8968
rect 11808 8965 11836 8996
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12544 9024 12572 9064
rect 12710 9052 12716 9064
rect 12768 9092 12774 9104
rect 17405 9095 17463 9101
rect 12768 9064 13492 9092
rect 12768 9052 12774 9064
rect 12986 9024 12992 9036
rect 12544 8996 12992 9024
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 13170 8984 13176 9036
rect 13228 9024 13234 9036
rect 13265 9027 13323 9033
rect 13265 9024 13277 9027
rect 13228 8996 13277 9024
rect 13228 8984 13234 8996
rect 13265 8993 13277 8996
rect 13311 8993 13323 9027
rect 13265 8987 13323 8993
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11480 8928 11805 8956
rect 11480 8916 11486 8928
rect 11793 8925 11805 8928
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 13464 8965 13492 9064
rect 17405 9061 17417 9095
rect 17451 9092 17463 9095
rect 17865 9095 17923 9101
rect 17865 9092 17877 9095
rect 17451 9064 17877 9092
rect 17451 9061 17463 9064
rect 17405 9055 17463 9061
rect 17865 9061 17877 9064
rect 17911 9092 17923 9095
rect 19058 9092 19064 9104
rect 17911 9064 19064 9092
rect 17911 9061 17923 9064
rect 17865 9055 17923 9061
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 24489 9095 24547 9101
rect 24489 9061 24501 9095
rect 24535 9092 24547 9095
rect 25038 9092 25044 9104
rect 24535 9064 25044 9092
rect 24535 9061 24547 9064
rect 24489 9055 24547 9061
rect 25038 9052 25044 9064
rect 25096 9052 25102 9104
rect 17880 8996 18092 9024
rect 17880 8968 17908 8996
rect 13449 8959 13507 8965
rect 11940 8928 11985 8956
rect 11940 8916 11946 8928
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 16390 8956 16396 8968
rect 16351 8928 16396 8956
rect 13449 8919 13507 8925
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 16482 8916 16488 8968
rect 16540 8956 16546 8968
rect 16540 8928 16585 8956
rect 16540 8916 16546 8928
rect 17862 8916 17868 8968
rect 17920 8916 17926 8968
rect 18064 8965 18092 8996
rect 18138 8984 18144 9036
rect 18196 9024 18202 9036
rect 19429 9027 19487 9033
rect 19429 9024 19441 9027
rect 18196 8996 19441 9024
rect 18196 8984 18202 8996
rect 19429 8993 19441 8996
rect 19475 9024 19487 9027
rect 19794 9024 19800 9036
rect 19475 8996 19800 9024
rect 19475 8993 19487 8996
rect 19429 8987 19487 8993
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 21913 9027 21971 9033
rect 21913 8993 21925 9027
rect 21959 9024 21971 9027
rect 23382 9024 23388 9036
rect 21959 8996 23388 9024
rect 21959 8993 21971 8996
rect 21913 8987 21971 8993
rect 23382 8984 23388 8996
rect 23440 8984 23446 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 18049 8959 18107 8965
rect 18049 8925 18061 8959
rect 18095 8925 18107 8959
rect 18049 8919 18107 8925
rect 12802 8848 12808 8900
rect 12860 8888 12866 8900
rect 12897 8891 12955 8897
rect 12897 8888 12909 8891
rect 12860 8860 12909 8888
rect 12860 8848 12866 8860
rect 12897 8857 12909 8860
rect 12943 8857 12955 8891
rect 17972 8888 18000 8919
rect 18874 8916 18880 8968
rect 18932 8956 18938 8968
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 18932 8928 19533 8956
rect 18932 8916 18938 8928
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 19702 8956 19708 8968
rect 19663 8928 19708 8956
rect 19521 8919 19579 8925
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 22002 8956 22008 8968
rect 21963 8928 22008 8956
rect 22002 8916 22008 8928
rect 22060 8916 22066 8968
rect 22097 8959 22155 8965
rect 22097 8925 22109 8959
rect 22143 8925 22155 8959
rect 23842 8956 23848 8968
rect 23803 8928 23848 8956
rect 22097 8919 22155 8925
rect 18322 8888 18328 8900
rect 17972 8860 18328 8888
rect 12897 8851 12955 8857
rect 18322 8848 18328 8860
rect 18380 8888 18386 8900
rect 19061 8891 19119 8897
rect 19061 8888 19073 8891
rect 18380 8860 19073 8888
rect 18380 8848 18386 8860
rect 19061 8857 19073 8860
rect 19107 8857 19119 8891
rect 19061 8851 19119 8857
rect 21818 8848 21824 8900
rect 21876 8888 21882 8900
rect 22112 8888 22140 8919
rect 23842 8916 23848 8928
rect 23900 8916 23906 8968
rect 25498 8956 25504 8968
rect 25411 8928 25504 8956
rect 25498 8916 25504 8928
rect 25556 8956 25562 8968
rect 25556 8928 25912 8956
rect 25556 8916 25562 8928
rect 21876 8860 22140 8888
rect 21876 8848 21882 8860
rect 25884 8832 25912 8928
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 3053 8823 3111 8829
rect 3053 8820 3065 8823
rect 2924 8792 3065 8820
rect 2924 8780 2930 8792
rect 3053 8789 3065 8792
rect 3099 8789 3111 8823
rect 3694 8820 3700 8832
rect 3655 8792 3700 8820
rect 3053 8783 3111 8789
rect 3694 8780 3700 8792
rect 3752 8780 3758 8832
rect 6641 8823 6699 8829
rect 6641 8789 6653 8823
rect 6687 8820 6699 8823
rect 7006 8820 7012 8832
rect 6687 8792 7012 8820
rect 6687 8789 6699 8792
rect 6641 8783 6699 8789
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 11333 8823 11391 8829
rect 11333 8789 11345 8823
rect 11379 8820 11391 8823
rect 12342 8820 12348 8832
rect 11379 8792 12348 8820
rect 11379 8789 11391 8792
rect 11333 8783 11391 8789
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 14093 8823 14151 8829
rect 14093 8789 14105 8823
rect 14139 8820 14151 8823
rect 14182 8820 14188 8832
rect 14139 8792 14188 8820
rect 14139 8789 14151 8792
rect 14093 8783 14151 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 14274 8780 14280 8832
rect 14332 8820 14338 8832
rect 14461 8823 14519 8829
rect 14461 8820 14473 8823
rect 14332 8792 14473 8820
rect 14332 8780 14338 8792
rect 14461 8789 14473 8792
rect 14507 8820 14519 8823
rect 14642 8820 14648 8832
rect 14507 8792 14648 8820
rect 14507 8789 14519 8792
rect 14461 8783 14519 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15838 8780 15844 8832
rect 15896 8820 15902 8832
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 15896 8792 15945 8820
rect 15896 8780 15902 8792
rect 15933 8789 15945 8792
rect 15979 8789 15991 8823
rect 17494 8820 17500 8832
rect 17455 8792 17500 8820
rect 15933 8783 15991 8789
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 21542 8820 21548 8832
rect 21503 8792 21548 8820
rect 21542 8780 21548 8792
rect 21600 8780 21606 8832
rect 23750 8820 23756 8832
rect 23663 8792 23756 8820
rect 23750 8780 23756 8792
rect 23808 8820 23814 8832
rect 24670 8820 24676 8832
rect 23808 8792 24676 8820
rect 23808 8780 23814 8792
rect 24670 8780 24676 8792
rect 24728 8780 24734 8832
rect 25866 8820 25872 8832
rect 25827 8792 25872 8820
rect 25866 8780 25872 8792
rect 25924 8780 25930 8832
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 7064 8588 8217 8616
rect 7064 8576 7070 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 8205 8579 8263 8585
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 13354 8616 13360 8628
rect 12299 8588 13360 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13633 8619 13691 8625
rect 13633 8585 13645 8619
rect 13679 8616 13691 8619
rect 14090 8616 14096 8628
rect 13679 8588 14096 8616
rect 13679 8585 13691 8588
rect 13633 8579 13691 8585
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 16298 8616 16304 8628
rect 15243 8588 16304 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 17589 8619 17647 8625
rect 17589 8585 17601 8619
rect 17635 8616 17647 8619
rect 17862 8616 17868 8628
rect 17635 8588 17868 8616
rect 17635 8585 17647 8588
rect 17589 8579 17647 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18046 8576 18052 8628
rect 18104 8616 18110 8628
rect 18417 8619 18475 8625
rect 18417 8616 18429 8619
rect 18104 8588 18429 8616
rect 18104 8576 18110 8588
rect 18417 8585 18429 8588
rect 18463 8585 18475 8619
rect 18417 8579 18475 8585
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 18969 8619 19027 8625
rect 18969 8616 18981 8619
rect 18748 8588 18981 8616
rect 18748 8576 18754 8588
rect 18969 8585 18981 8588
rect 19015 8585 19027 8619
rect 19702 8616 19708 8628
rect 18969 8579 19027 8585
rect 19536 8588 19708 8616
rect 1578 8548 1584 8560
rect 1539 8520 1584 8548
rect 1578 8508 1584 8520
rect 1636 8508 1642 8560
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 9861 8551 9919 8557
rect 9861 8548 9873 8551
rect 9364 8520 9873 8548
rect 9364 8508 9370 8520
rect 9861 8517 9873 8520
rect 9907 8548 9919 8551
rect 12989 8551 13047 8557
rect 9907 8520 10180 8548
rect 9907 8517 9919 8520
rect 9861 8511 9919 8517
rect 3694 8440 3700 8492
rect 3752 8480 3758 8492
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 3752 8452 4261 8480
rect 3752 8440 3758 8452
rect 4249 8449 4261 8452
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2038 8412 2044 8424
rect 1443 8384 2044 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4062 8412 4068 8424
rect 4019 8384 4068 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 2498 8304 2504 8356
rect 2556 8344 2562 8356
rect 2593 8347 2651 8353
rect 2593 8344 2605 8347
rect 2556 8316 2605 8344
rect 2556 8304 2562 8316
rect 2593 8313 2605 8316
rect 2639 8344 2651 8347
rect 3513 8347 3571 8353
rect 3513 8344 3525 8347
rect 2639 8316 3525 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 3513 8313 3525 8316
rect 3559 8344 3571 8347
rect 3878 8344 3884 8356
rect 3559 8316 3884 8344
rect 3559 8313 3571 8316
rect 3513 8307 3571 8313
rect 3878 8304 3884 8316
rect 3936 8344 3942 8356
rect 3936 8316 4108 8344
rect 3936 8304 3942 8316
rect 3602 8276 3608 8288
rect 3563 8248 3608 8276
rect 3602 8236 3608 8248
rect 3660 8236 3666 8288
rect 4080 8285 4108 8316
rect 4065 8279 4123 8285
rect 4065 8245 4077 8279
rect 4111 8245 4123 8279
rect 4264 8276 4292 8443
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6546 8480 6552 8492
rect 6328 8452 6552 8480
rect 6328 8440 6334 8452
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6696 8384 6837 8412
rect 6696 8372 6702 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 10042 8412 10048 8424
rect 10003 8384 10048 8412
rect 6825 8375 6883 8381
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10152 8421 10180 8520
rect 12989 8517 13001 8551
rect 13035 8548 13047 8551
rect 13170 8548 13176 8560
rect 13035 8520 13176 8548
rect 13035 8517 13047 8520
rect 12989 8511 13047 8517
rect 13170 8508 13176 8520
rect 13228 8508 13234 8560
rect 17037 8551 17095 8557
rect 17037 8517 17049 8551
rect 17083 8517 17095 8551
rect 17037 8511 17095 8517
rect 10137 8415 10195 8421
rect 10137 8381 10149 8415
rect 10183 8412 10195 8415
rect 10226 8412 10232 8424
rect 10183 8384 10232 8412
rect 10183 8381 10195 8384
rect 10137 8375 10195 8381
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 15657 8415 15715 8421
rect 15657 8412 15669 8415
rect 15304 8384 15669 8412
rect 15304 8356 15332 8384
rect 15657 8381 15669 8384
rect 15703 8381 15715 8415
rect 16482 8412 16488 8424
rect 15657 8375 15715 8381
rect 15764 8384 16488 8412
rect 6546 8344 6552 8356
rect 6507 8316 6552 8344
rect 6546 8304 6552 8316
rect 6604 8344 6610 8356
rect 7070 8347 7128 8353
rect 7070 8344 7082 8347
rect 6604 8316 7082 8344
rect 6604 8304 6610 8316
rect 7070 8313 7082 8316
rect 7116 8313 7128 8347
rect 7070 8307 7128 8313
rect 9769 8347 9827 8353
rect 9769 8313 9781 8347
rect 9815 8344 9827 8347
rect 10404 8347 10462 8353
rect 10404 8344 10416 8347
rect 9815 8316 10416 8344
rect 9815 8313 9827 8316
rect 9769 8307 9827 8313
rect 10404 8313 10416 8316
rect 10450 8344 10462 8347
rect 10594 8344 10600 8356
rect 10450 8316 10600 8344
rect 10450 8313 10462 8316
rect 10404 8307 10462 8313
rect 10594 8304 10600 8316
rect 10652 8304 10658 8356
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8344 14887 8347
rect 15286 8344 15292 8356
rect 14875 8316 15292 8344
rect 14875 8313 14887 8316
rect 14829 8307 14887 8313
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 15470 8344 15476 8356
rect 15431 8316 15476 8344
rect 15470 8304 15476 8316
rect 15528 8344 15534 8356
rect 15764 8344 15792 8384
rect 16482 8372 16488 8384
rect 16540 8412 16546 8424
rect 17052 8412 17080 8511
rect 19426 8480 19432 8492
rect 19387 8452 19432 8480
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 19536 8489 19564 8588
rect 19702 8576 19708 8588
rect 19760 8616 19766 8628
rect 19981 8619 20039 8625
rect 19981 8616 19993 8619
rect 19760 8588 19993 8616
rect 19760 8576 19766 8588
rect 19981 8585 19993 8588
rect 20027 8585 20039 8619
rect 20530 8616 20536 8628
rect 20491 8588 20536 8616
rect 19981 8579 20039 8585
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 21637 8619 21695 8625
rect 21637 8585 21649 8619
rect 21683 8616 21695 8619
rect 21818 8616 21824 8628
rect 21683 8588 21824 8616
rect 21683 8585 21695 8588
rect 21637 8579 21695 8585
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 21913 8619 21971 8625
rect 21913 8585 21925 8619
rect 21959 8616 21971 8619
rect 22002 8616 22008 8628
rect 21959 8588 22008 8616
rect 21959 8585 21971 8588
rect 21913 8579 21971 8585
rect 22002 8576 22008 8588
rect 22060 8576 22066 8628
rect 23382 8616 23388 8628
rect 23343 8588 23388 8616
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 24486 8616 24492 8628
rect 24447 8588 24492 8616
rect 24486 8576 24492 8588
rect 24544 8576 24550 8628
rect 24949 8619 25007 8625
rect 24949 8585 24961 8619
rect 24995 8616 25007 8619
rect 25222 8616 25228 8628
rect 24995 8588 25228 8616
rect 24995 8585 25007 8588
rect 24949 8579 25007 8585
rect 25222 8576 25228 8588
rect 25280 8576 25286 8628
rect 25406 8616 25412 8628
rect 25367 8588 25412 8616
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 26510 8616 26516 8628
rect 26471 8588 26516 8616
rect 26510 8576 26516 8588
rect 26568 8576 26574 8628
rect 27154 8616 27160 8628
rect 27115 8588 27160 8616
rect 27154 8576 27160 8588
rect 27212 8576 27218 8628
rect 25240 8548 25268 8576
rect 27525 8551 27583 8557
rect 27525 8548 27537 8551
rect 25240 8520 27537 8548
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 21910 8440 21916 8492
rect 21968 8480 21974 8492
rect 22094 8480 22100 8492
rect 21968 8452 22100 8480
rect 21968 8440 21974 8452
rect 22094 8440 22100 8452
rect 22152 8480 22158 8492
rect 22465 8483 22523 8489
rect 22465 8480 22477 8483
rect 22152 8452 22477 8480
rect 22152 8440 22158 8452
rect 22465 8449 22477 8452
rect 22511 8449 22523 8483
rect 25314 8480 25320 8492
rect 25275 8452 25320 8480
rect 22465 8443 22523 8449
rect 25314 8440 25320 8452
rect 25372 8440 25378 8492
rect 25958 8440 25964 8492
rect 26016 8480 26022 8492
rect 26053 8483 26111 8489
rect 26053 8480 26065 8483
rect 26016 8452 26065 8480
rect 26016 8440 26022 8452
rect 26053 8449 26065 8452
rect 26099 8480 26111 8483
rect 26142 8480 26148 8492
rect 26099 8452 26148 8480
rect 26099 8449 26111 8452
rect 26053 8443 26111 8449
rect 26142 8440 26148 8452
rect 26200 8440 26206 8492
rect 16540 8384 17080 8412
rect 16540 8372 16546 8384
rect 18782 8372 18788 8424
rect 18840 8372 18846 8424
rect 18874 8372 18880 8424
rect 18932 8412 18938 8424
rect 19337 8415 19395 8421
rect 18932 8384 18977 8412
rect 18932 8372 18938 8384
rect 19337 8381 19349 8415
rect 19383 8412 19395 8415
rect 19610 8412 19616 8424
rect 19383 8384 19616 8412
rect 19383 8381 19395 8384
rect 19337 8375 19395 8381
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 20717 8415 20775 8421
rect 20717 8381 20729 8415
rect 20763 8381 20775 8415
rect 20717 8375 20775 8381
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 21818 8412 21824 8424
rect 21315 8384 21824 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 15930 8353 15936 8356
rect 15528 8316 15792 8344
rect 15528 8304 15534 8316
rect 15924 8307 15936 8353
rect 15988 8344 15994 8356
rect 17218 8344 17224 8356
rect 15988 8316 17224 8344
rect 15930 8304 15936 8307
rect 15988 8304 15994 8316
rect 17218 8304 17224 8316
rect 17276 8304 17282 8356
rect 18800 8344 18828 8372
rect 20349 8347 20407 8353
rect 20349 8344 20361 8347
rect 18800 8316 20361 8344
rect 20349 8313 20361 8316
rect 20395 8344 20407 8347
rect 20732 8344 20760 8375
rect 21818 8372 21824 8384
rect 21876 8412 21882 8424
rect 22373 8415 22431 8421
rect 22373 8412 22385 8415
rect 21876 8384 22385 8412
rect 21876 8372 21882 8384
rect 22373 8381 22385 8384
rect 22419 8381 22431 8415
rect 22373 8375 22431 8381
rect 23842 8372 23848 8424
rect 23900 8412 23906 8424
rect 25777 8415 25835 8421
rect 25777 8412 25789 8415
rect 23900 8384 25789 8412
rect 23900 8372 23906 8384
rect 25777 8381 25789 8384
rect 25823 8412 25835 8415
rect 25866 8412 25872 8424
rect 25823 8384 25872 8412
rect 25823 8381 25835 8384
rect 25777 8375 25835 8381
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 26988 8421 27016 8520
rect 27525 8517 27537 8520
rect 27571 8517 27583 8551
rect 27525 8511 27583 8517
rect 26973 8415 27031 8421
rect 26973 8381 26985 8415
rect 27019 8381 27031 8415
rect 26973 8375 27031 8381
rect 20395 8316 20760 8344
rect 20395 8313 20407 8316
rect 20349 8307 20407 8313
rect 24486 8304 24492 8356
rect 24544 8344 24550 8356
rect 24544 8316 25912 8344
rect 24544 8304 24550 8316
rect 4706 8276 4712 8288
rect 4264 8248 4712 8276
rect 4065 8239 4123 8245
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 6273 8279 6331 8285
rect 6273 8245 6285 8279
rect 6319 8276 6331 8279
rect 6638 8276 6644 8288
rect 6319 8248 6644 8276
rect 6319 8245 6331 8248
rect 6273 8239 6331 8245
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 11517 8279 11575 8285
rect 11517 8245 11529 8279
rect 11563 8276 11575 8279
rect 11882 8276 11888 8288
rect 11563 8248 11888 8276
rect 11563 8245 11575 8248
rect 11517 8239 11575 8245
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 22281 8279 22339 8285
rect 22281 8245 22293 8279
rect 22327 8276 22339 8279
rect 22370 8276 22376 8288
rect 22327 8248 22376 8276
rect 22327 8245 22339 8248
rect 22281 8239 22339 8245
rect 22370 8236 22376 8248
rect 22428 8276 22434 8288
rect 25884 8285 25912 8316
rect 22925 8279 22983 8285
rect 22925 8276 22937 8279
rect 22428 8248 22937 8276
rect 22428 8236 22434 8248
rect 22925 8245 22937 8248
rect 22971 8245 22983 8279
rect 22925 8239 22983 8245
rect 25869 8279 25927 8285
rect 25869 8245 25881 8279
rect 25915 8245 25927 8279
rect 25869 8239 25927 8245
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 1670 8072 1676 8084
rect 1631 8044 1676 8072
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 2317 8075 2375 8081
rect 2317 8041 2329 8075
rect 2363 8072 2375 8075
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2363 8044 2789 8072
rect 2363 8041 2375 8044
rect 2317 8035 2375 8041
rect 2777 8041 2789 8044
rect 2823 8072 2835 8075
rect 3602 8072 3608 8084
rect 2823 8044 3608 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 3697 8075 3755 8081
rect 3697 8041 3709 8075
rect 3743 8072 3755 8075
rect 4062 8072 4068 8084
rect 3743 8044 4068 8072
rect 3743 8041 3755 8044
rect 3697 8035 3755 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4396 8044 4445 8072
rect 4396 8032 4402 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 11422 8072 11428 8084
rect 11383 8044 11428 8072
rect 4433 8035 4491 8041
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 11698 8072 11704 8084
rect 11659 8044 11704 8072
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12526 8072 12532 8084
rect 12487 8044 12532 8072
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12710 8032 12716 8084
rect 12768 8072 12774 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12768 8044 12909 8072
rect 12768 8032 12774 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 12897 8035 12955 8041
rect 16117 8075 16175 8081
rect 16117 8041 16129 8075
rect 16163 8072 16175 8075
rect 16390 8072 16396 8084
rect 16163 8044 16396 8072
rect 16163 8041 16175 8044
rect 16117 8035 16175 8041
rect 16390 8032 16396 8044
rect 16448 8072 16454 8084
rect 17221 8075 17279 8081
rect 17221 8072 17233 8075
rect 16448 8044 17233 8072
rect 16448 8032 16454 8044
rect 17221 8041 17233 8044
rect 17267 8041 17279 8075
rect 17221 8035 17279 8041
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 17552 8044 17693 8072
rect 17552 8032 17558 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 18322 8072 18328 8084
rect 18283 8044 18328 8072
rect 17681 8035 17739 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 19061 8075 19119 8081
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 19242 8072 19248 8084
rect 19107 8044 19248 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 19429 8075 19487 8081
rect 19429 8041 19441 8075
rect 19475 8072 19487 8075
rect 19610 8072 19616 8084
rect 19475 8044 19616 8072
rect 19475 8041 19487 8044
rect 19429 8035 19487 8041
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 19702 8032 19708 8084
rect 19760 8072 19766 8084
rect 21637 8075 21695 8081
rect 19760 8044 19805 8072
rect 19760 8032 19766 8044
rect 21637 8041 21649 8075
rect 21683 8072 21695 8075
rect 22002 8072 22008 8084
rect 21683 8044 22008 8072
rect 21683 8041 21695 8044
rect 21637 8035 21695 8041
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 22370 8072 22376 8084
rect 22331 8044 22376 8072
rect 22370 8032 22376 8044
rect 22428 8032 22434 8084
rect 23753 8075 23811 8081
rect 23753 8041 23765 8075
rect 23799 8072 23811 8075
rect 23934 8072 23940 8084
rect 23799 8044 23940 8072
rect 23799 8041 23811 8044
rect 23753 8035 23811 8041
rect 23934 8032 23940 8044
rect 23992 8072 23998 8084
rect 25130 8072 25136 8084
rect 23992 8044 25136 8072
rect 23992 8032 23998 8044
rect 25130 8032 25136 8044
rect 25188 8032 25194 8084
rect 25866 8072 25872 8084
rect 25827 8044 25872 8072
rect 25866 8032 25872 8044
rect 25924 8032 25930 8084
rect 26694 8072 26700 8084
rect 26655 8044 26700 8072
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 4525 8007 4583 8013
rect 4525 7973 4537 8007
rect 4571 8004 4583 8007
rect 4614 8004 4620 8016
rect 4571 7976 4620 8004
rect 4571 7973 4583 7976
rect 4525 7967 4583 7973
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 10318 8004 10324 8016
rect 10279 7976 10324 8004
rect 10318 7964 10324 7976
rect 10376 7964 10382 8016
rect 17589 8007 17647 8013
rect 17589 7973 17601 8007
rect 17635 8004 17647 8007
rect 17862 8004 17868 8016
rect 17635 7976 17868 8004
rect 17635 7973 17647 7976
rect 17589 7967 17647 7973
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 21910 8004 21916 8016
rect 21871 7976 21916 8004
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 24949 8007 25007 8013
rect 22664 7976 24808 8004
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 7101 7939 7159 7945
rect 7101 7936 7113 7939
rect 6328 7908 7113 7936
rect 6328 7896 6334 7908
rect 7101 7905 7113 7908
rect 7147 7936 7159 7939
rect 9030 7936 9036 7948
rect 7147 7908 9036 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 9030 7896 9036 7908
rect 9088 7936 9094 7948
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 9088 7908 9873 7936
rect 9088 7896 9094 7908
rect 9861 7905 9873 7908
rect 9907 7936 9919 7939
rect 10042 7936 10048 7948
rect 9907 7908 10048 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 17126 7936 17132 7948
rect 17087 7908 17132 7936
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 21358 7896 21364 7948
rect 21416 7936 21422 7948
rect 22664 7936 22692 7976
rect 21416 7908 22692 7936
rect 22741 7939 22799 7945
rect 21416 7896 21422 7908
rect 22741 7905 22753 7939
rect 22787 7936 22799 7939
rect 23106 7936 23112 7948
rect 22787 7908 23112 7936
rect 22787 7905 22799 7908
rect 22741 7899 22799 7905
rect 23106 7896 23112 7908
rect 23164 7896 23170 7948
rect 24780 7936 24808 7976
rect 24949 7973 24961 8007
rect 24995 8004 25007 8007
rect 26326 8004 26332 8016
rect 24995 7976 26332 8004
rect 24995 7973 25007 7976
rect 24949 7967 25007 7973
rect 26326 7964 26332 7976
rect 26384 7964 26390 8016
rect 25038 7936 25044 7948
rect 24780 7908 25044 7936
rect 25038 7896 25044 7908
rect 25096 7936 25102 7948
rect 25317 7939 25375 7945
rect 25317 7936 25329 7939
rect 25096 7908 25329 7936
rect 25096 7896 25102 7908
rect 25317 7905 25329 7908
rect 25363 7905 25375 7939
rect 26510 7936 26516 7948
rect 26471 7908 26516 7936
rect 25317 7899 25375 7905
rect 26510 7896 26516 7908
rect 26568 7896 26574 7948
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3878 7868 3884 7880
rect 3099 7840 3884 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 2682 7760 2688 7812
rect 2740 7800 2746 7812
rect 2884 7800 2912 7831
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 17034 7868 17040 7880
rect 10560 7840 17040 7868
rect 10560 7828 10566 7840
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 17276 7840 17785 7868
rect 17276 7828 17282 7840
rect 17773 7837 17785 7840
rect 17819 7837 17831 7871
rect 22830 7868 22836 7880
rect 22791 7840 22836 7868
rect 17773 7831 17831 7837
rect 22830 7828 22836 7840
rect 22888 7828 22894 7880
rect 22922 7828 22928 7880
rect 22980 7868 22986 7880
rect 23017 7871 23075 7877
rect 23017 7868 23029 7871
rect 22980 7840 23029 7868
rect 22980 7828 22986 7840
rect 23017 7837 23029 7840
rect 23063 7868 23075 7871
rect 23382 7868 23388 7880
rect 23063 7840 23388 7868
rect 23063 7837 23075 7840
rect 23017 7831 23075 7837
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 4065 7803 4123 7809
rect 4065 7800 4077 7803
rect 2740 7772 4077 7800
rect 2740 7760 2746 7772
rect 4065 7769 4077 7772
rect 4111 7769 4123 7803
rect 4065 7763 4123 7769
rect 2406 7732 2412 7744
rect 2367 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 6638 7692 6644 7744
rect 6696 7732 6702 7744
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 6696 7704 6929 7732
rect 6696 7692 6702 7704
rect 6917 7701 6929 7704
rect 6963 7732 6975 7735
rect 7377 7735 7435 7741
rect 7377 7732 7389 7735
rect 6963 7704 7389 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7377 7701 7389 7704
rect 7423 7701 7435 7735
rect 7377 7695 7435 7701
rect 15749 7735 15807 7741
rect 15749 7701 15761 7735
rect 15795 7732 15807 7735
rect 16390 7732 16396 7744
rect 15795 7704 16396 7732
rect 15795 7701 15807 7704
rect 15749 7695 15807 7701
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 16482 7692 16488 7744
rect 16540 7732 16546 7744
rect 16945 7735 17003 7741
rect 16945 7732 16957 7735
rect 16540 7704 16957 7732
rect 16540 7692 16546 7704
rect 16945 7701 16957 7704
rect 16991 7732 17003 7735
rect 17402 7732 17408 7744
rect 16991 7704 17408 7732
rect 16991 7701 17003 7704
rect 16945 7695 17003 7701
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 24118 7732 24124 7744
rect 24079 7704 24124 7732
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 25498 7732 25504 7744
rect 25459 7704 25504 7732
rect 25498 7692 25504 7704
rect 25556 7692 25562 7744
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 4249 7531 4307 7537
rect 4249 7497 4261 7531
rect 4295 7528 4307 7531
rect 4338 7528 4344 7540
rect 4295 7500 4344 7528
rect 4295 7497 4307 7500
rect 4249 7491 4307 7497
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 6270 7528 6276 7540
rect 6231 7500 6276 7528
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 6604 7500 8217 7528
rect 6604 7488 6610 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 8205 7491 8263 7497
rect 16945 7531 17003 7537
rect 16945 7497 16957 7531
rect 16991 7528 17003 7531
rect 17494 7528 17500 7540
rect 16991 7500 17500 7528
rect 16991 7497 17003 7500
rect 16945 7491 17003 7497
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 18509 7531 18567 7537
rect 18509 7528 18521 7531
rect 18472 7500 18521 7528
rect 18472 7488 18478 7500
rect 18509 7497 18521 7500
rect 18555 7497 18567 7531
rect 18509 7491 18567 7497
rect 17218 7460 17224 7472
rect 17179 7432 17224 7460
rect 17218 7420 17224 7432
rect 17276 7420 17282 7472
rect 4614 7392 4620 7404
rect 4575 7364 4620 7392
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 6696 7364 6837 7392
rect 6696 7352 6702 7364
rect 6825 7361 6837 7364
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 12250 7352 12256 7404
rect 12308 7392 12314 7404
rect 12434 7392 12440 7404
rect 12308 7364 12440 7392
rect 12308 7352 12314 7364
rect 12434 7352 12440 7364
rect 12492 7392 12498 7404
rect 12492 7364 12585 7392
rect 12492 7352 12498 7364
rect 15194 7352 15200 7404
rect 15252 7392 15258 7404
rect 16209 7395 16267 7401
rect 16209 7392 16221 7395
rect 15252 7364 16221 7392
rect 15252 7352 15258 7364
rect 16209 7361 16221 7364
rect 16255 7361 16267 7395
rect 18524 7392 18552 7491
rect 21818 7488 21824 7540
rect 21876 7528 21882 7540
rect 22005 7531 22063 7537
rect 22005 7528 22017 7531
rect 21876 7500 22017 7528
rect 21876 7488 21882 7500
rect 22005 7497 22017 7500
rect 22051 7497 22063 7531
rect 25038 7528 25044 7540
rect 24999 7500 25044 7528
rect 22005 7491 22063 7497
rect 25038 7488 25044 7500
rect 25096 7488 25102 7540
rect 26510 7488 26516 7540
rect 26568 7528 26574 7540
rect 26881 7531 26939 7537
rect 26881 7528 26893 7531
rect 26568 7500 26893 7528
rect 26568 7488 26574 7500
rect 26881 7497 26893 7500
rect 26927 7497 26939 7531
rect 27614 7528 27620 7540
rect 27575 7500 27620 7528
rect 26881 7491 26939 7497
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 22830 7420 22836 7472
rect 22888 7460 22894 7472
rect 23661 7463 23719 7469
rect 23661 7460 23673 7463
rect 22888 7432 23673 7460
rect 22888 7420 22894 7432
rect 23661 7429 23673 7432
rect 23707 7429 23719 7463
rect 23661 7423 23719 7429
rect 26326 7420 26332 7472
rect 26384 7460 26390 7472
rect 26605 7463 26663 7469
rect 26605 7460 26617 7463
rect 26384 7432 26617 7460
rect 26384 7420 26390 7432
rect 26605 7429 26617 7432
rect 26651 7429 26663 7463
rect 26605 7423 26663 7429
rect 19153 7395 19211 7401
rect 19153 7392 19165 7395
rect 18524 7364 19165 7392
rect 16209 7355 16267 7361
rect 19153 7361 19165 7364
rect 19199 7361 19211 7395
rect 19153 7355 19211 7361
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7392 19395 7395
rect 19426 7392 19432 7404
rect 19383 7364 19432 7392
rect 19383 7361 19395 7364
rect 19337 7355 19395 7361
rect 19426 7352 19432 7364
rect 19484 7392 19490 7404
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 19484 7364 19717 7392
rect 19484 7352 19490 7364
rect 19705 7361 19717 7364
rect 19751 7361 19763 7395
rect 19705 7355 19763 7361
rect 21913 7395 21971 7401
rect 21913 7361 21925 7395
rect 21959 7392 21971 7395
rect 22278 7392 22284 7404
rect 21959 7364 22284 7392
rect 21959 7361 21971 7364
rect 21913 7355 21971 7361
rect 22278 7352 22284 7364
rect 22336 7392 22342 7404
rect 22649 7395 22707 7401
rect 22649 7392 22661 7395
rect 22336 7364 22661 7392
rect 22336 7352 22342 7364
rect 22649 7361 22661 7364
rect 22695 7392 22707 7395
rect 22922 7392 22928 7404
rect 22695 7364 22928 7392
rect 22695 7361 22707 7364
rect 22649 7355 22707 7361
rect 22922 7352 22928 7364
rect 22980 7352 22986 7404
rect 24118 7352 24124 7404
rect 24176 7392 24182 7404
rect 24213 7395 24271 7401
rect 24213 7392 24225 7395
rect 24176 7364 24225 7392
rect 24176 7352 24182 7364
rect 24213 7361 24225 7364
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7293 1455 7327
rect 1397 7287 1455 7293
rect 1412 7256 1440 7287
rect 1946 7284 1952 7336
rect 2004 7324 2010 7336
rect 2501 7327 2559 7333
rect 2501 7324 2513 7327
rect 2004 7296 2513 7324
rect 2004 7284 2010 7296
rect 2501 7293 2513 7296
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9122 7324 9128 7336
rect 9079 7296 9128 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9122 7284 9128 7296
rect 9180 7324 9186 7336
rect 10318 7324 10324 7336
rect 9180 7296 10324 7324
rect 9180 7284 9186 7296
rect 10318 7284 10324 7296
rect 10376 7284 10382 7336
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7324 15623 7327
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15611 7296 16037 7324
rect 15611 7293 15623 7296
rect 15565 7287 15623 7293
rect 16025 7293 16037 7296
rect 16071 7324 16083 7327
rect 16298 7324 16304 7336
rect 16071 7296 16304 7324
rect 16071 7293 16083 7296
rect 16025 7287 16083 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 23934 7284 23940 7336
rect 23992 7324 23998 7336
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23992 7296 24041 7324
rect 23992 7284 23998 7296
rect 24029 7293 24041 7296
rect 24075 7293 24087 7327
rect 25225 7327 25283 7333
rect 25225 7324 25237 7327
rect 24029 7287 24087 7293
rect 24688 7296 25237 7324
rect 2038 7256 2044 7268
rect 1412 7228 2044 7256
rect 2038 7216 2044 7228
rect 2096 7216 2102 7268
rect 2409 7259 2467 7265
rect 2409 7225 2421 7259
rect 2455 7256 2467 7259
rect 2768 7259 2826 7265
rect 2768 7256 2780 7259
rect 2455 7228 2780 7256
rect 2455 7225 2467 7228
rect 2409 7219 2467 7225
rect 2768 7225 2780 7228
rect 2814 7256 2826 7259
rect 6641 7259 6699 7265
rect 2814 7228 4016 7256
rect 2814 7225 2826 7228
rect 2768 7219 2826 7225
rect 3988 7200 4016 7228
rect 6641 7225 6653 7259
rect 6687 7256 6699 7259
rect 7006 7256 7012 7268
rect 6687 7228 7012 7256
rect 6687 7225 6699 7228
rect 6641 7219 6699 7225
rect 7006 7216 7012 7228
rect 7064 7265 7070 7268
rect 7064 7259 7128 7265
rect 7064 7225 7082 7259
rect 7116 7225 7128 7259
rect 7064 7219 7128 7225
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 9300 7259 9358 7265
rect 9300 7256 9312 7259
rect 8987 7228 9312 7256
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 9300 7225 9312 7228
rect 9346 7256 9358 7259
rect 9582 7256 9588 7268
rect 9346 7228 9588 7256
rect 9346 7225 9358 7228
rect 9300 7219 9358 7225
rect 7064 7216 7070 7219
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 11882 7216 11888 7268
rect 11940 7256 11946 7268
rect 12253 7259 12311 7265
rect 12253 7256 12265 7259
rect 11940 7228 12265 7256
rect 11940 7216 11946 7228
rect 12253 7225 12265 7228
rect 12299 7256 12311 7259
rect 12682 7259 12740 7265
rect 12682 7256 12694 7259
rect 12299 7228 12694 7256
rect 12299 7225 12311 7228
rect 12253 7219 12311 7225
rect 12682 7225 12694 7228
rect 12728 7225 12740 7259
rect 12682 7219 12740 7225
rect 16117 7259 16175 7265
rect 16117 7225 16129 7259
rect 16163 7256 16175 7259
rect 16390 7256 16396 7268
rect 16163 7228 16396 7256
rect 16163 7225 16175 7228
rect 16117 7219 16175 7225
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 17770 7216 17776 7268
rect 17828 7256 17834 7268
rect 17865 7259 17923 7265
rect 17865 7256 17877 7259
rect 17828 7228 17877 7256
rect 17828 7216 17834 7228
rect 17865 7225 17877 7228
rect 17911 7256 17923 7259
rect 19061 7259 19119 7265
rect 19061 7256 19073 7259
rect 17911 7228 19073 7256
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 19061 7225 19073 7228
rect 19107 7225 19119 7259
rect 19061 7219 19119 7225
rect 21545 7259 21603 7265
rect 21545 7225 21557 7259
rect 21591 7256 21603 7259
rect 22373 7259 22431 7265
rect 22373 7256 22385 7259
rect 21591 7228 22385 7256
rect 21591 7225 21603 7228
rect 21545 7219 21603 7225
rect 22373 7225 22385 7228
rect 22419 7256 22431 7259
rect 23382 7256 23388 7268
rect 22419 7228 23388 7256
rect 22419 7225 22431 7228
rect 22373 7219 22431 7225
rect 23382 7216 23388 7228
rect 23440 7216 23446 7268
rect 23477 7259 23535 7265
rect 23477 7225 23489 7259
rect 23523 7256 23535 7259
rect 23523 7228 24164 7256
rect 23523 7225 23535 7228
rect 23477 7219 23535 7225
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 3878 7188 3884 7200
rect 3839 7160 3884 7188
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 4706 7188 4712 7200
rect 4028 7160 4712 7188
rect 4028 7148 4034 7160
rect 4706 7148 4712 7160
rect 4764 7188 4770 7200
rect 4893 7191 4951 7197
rect 4893 7188 4905 7191
rect 4764 7160 4905 7188
rect 4764 7148 4770 7160
rect 4893 7157 4905 7160
rect 4939 7157 4951 7191
rect 10410 7188 10416 7200
rect 10371 7160 10416 7188
rect 4893 7151 4951 7157
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7188 13875 7191
rect 13906 7188 13912 7200
rect 13863 7160 13912 7188
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 15194 7188 15200 7200
rect 15155 7160 15200 7188
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 15654 7188 15660 7200
rect 15615 7160 15660 7188
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 18690 7188 18696 7200
rect 18651 7160 18696 7188
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 22462 7188 22468 7200
rect 22423 7160 22468 7188
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 23106 7188 23112 7200
rect 23067 7160 23112 7188
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 24136 7197 24164 7228
rect 24688 7200 24716 7296
rect 25225 7293 25237 7296
rect 25271 7293 25283 7327
rect 27430 7324 27436 7336
rect 27391 7296 27436 7324
rect 25225 7287 25283 7293
rect 27430 7284 27436 7296
rect 27488 7324 27494 7336
rect 27985 7327 28043 7333
rect 27985 7324 27997 7327
rect 27488 7296 27997 7324
rect 27488 7284 27494 7296
rect 27985 7293 27997 7296
rect 28031 7293 28043 7327
rect 27985 7287 28043 7293
rect 25470 7259 25528 7265
rect 25470 7256 25482 7259
rect 25240 7228 25482 7256
rect 25240 7200 25268 7228
rect 25470 7225 25482 7228
rect 25516 7225 25528 7259
rect 25470 7219 25528 7225
rect 24121 7191 24179 7197
rect 24121 7157 24133 7191
rect 24167 7188 24179 7191
rect 24302 7188 24308 7200
rect 24167 7160 24308 7188
rect 24167 7157 24179 7160
rect 24121 7151 24179 7157
rect 24302 7148 24308 7160
rect 24360 7148 24366 7200
rect 24670 7188 24676 7200
rect 24631 7160 24676 7188
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 25222 7148 25228 7200
rect 25280 7148 25286 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 9122 6984 9128 6996
rect 9083 6956 9128 6984
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10045 6987 10103 6993
rect 10045 6984 10057 6987
rect 9732 6956 10057 6984
rect 9732 6944 9738 6956
rect 10045 6953 10057 6956
rect 10091 6984 10103 6987
rect 11241 6987 11299 6993
rect 11241 6984 11253 6987
rect 10091 6956 11253 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 11241 6953 11253 6956
rect 11287 6953 11299 6987
rect 11241 6947 11299 6953
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17589 6987 17647 6993
rect 17589 6984 17601 6987
rect 17184 6956 17601 6984
rect 17184 6944 17190 6956
rect 17589 6953 17601 6956
rect 17635 6953 17647 6987
rect 17770 6984 17776 6996
rect 17731 6956 17776 6984
rect 17589 6947 17647 6953
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 19150 6984 19156 6996
rect 19111 6956 19156 6984
rect 19150 6944 19156 6956
rect 19208 6944 19214 6996
rect 19610 6944 19616 6996
rect 19668 6984 19674 6996
rect 19889 6987 19947 6993
rect 19889 6984 19901 6987
rect 19668 6956 19901 6984
rect 19668 6944 19674 6956
rect 19889 6953 19901 6956
rect 19935 6984 19947 6987
rect 20530 6984 20536 6996
rect 19935 6956 20536 6984
rect 19935 6953 19947 6956
rect 19889 6947 19947 6953
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 22097 6987 22155 6993
rect 22097 6953 22109 6987
rect 22143 6984 22155 6987
rect 22462 6984 22468 6996
rect 22143 6956 22468 6984
rect 22143 6953 22155 6956
rect 22097 6947 22155 6953
rect 22462 6944 22468 6956
rect 22520 6984 22526 6996
rect 23017 6987 23075 6993
rect 23017 6984 23029 6987
rect 22520 6956 23029 6984
rect 22520 6944 22526 6956
rect 23017 6953 23029 6956
rect 23063 6953 23075 6987
rect 23017 6947 23075 6953
rect 23290 6944 23296 6996
rect 23348 6984 23354 6996
rect 23385 6987 23443 6993
rect 23385 6984 23397 6987
rect 23348 6956 23397 6984
rect 23348 6944 23354 6956
rect 23385 6953 23397 6956
rect 23431 6953 23443 6987
rect 23385 6947 23443 6953
rect 17313 6919 17371 6925
rect 17313 6885 17325 6919
rect 17359 6916 17371 6919
rect 17862 6916 17868 6928
rect 17359 6888 17868 6916
rect 17359 6885 17371 6888
rect 17313 6879 17371 6885
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 22278 6876 22284 6928
rect 22336 6916 22342 6928
rect 22373 6919 22431 6925
rect 22373 6916 22385 6919
rect 22336 6888 22385 6916
rect 22336 6876 22342 6888
rect 22373 6885 22385 6888
rect 22419 6885 22431 6919
rect 22830 6916 22836 6928
rect 22791 6888 22836 6916
rect 22373 6879 22431 6885
rect 22830 6876 22836 6888
rect 22888 6876 22894 6928
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2130 6848 2136 6860
rect 1443 6820 2136 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 2498 6848 2504 6860
rect 2459 6820 2504 6848
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2682 6808 2688 6860
rect 2740 6808 2746 6860
rect 6822 6848 6828 6860
rect 6783 6820 6828 6848
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 11606 6848 11612 6860
rect 11567 6820 11612 6848
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 11701 6851 11759 6857
rect 11701 6817 11713 6851
rect 11747 6848 11759 6851
rect 11790 6848 11796 6860
rect 11747 6820 11796 6848
rect 11747 6817 11759 6820
rect 11701 6811 11759 6817
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 13446 6848 13452 6860
rect 12676 6820 13452 6848
rect 12676 6808 12682 6820
rect 13446 6808 13452 6820
rect 13504 6848 13510 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13504 6820 13737 6848
rect 13504 6808 13510 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 15545 6851 15603 6857
rect 15545 6848 15557 6851
rect 13725 6811 13783 6817
rect 13924 6820 15557 6848
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2700 6780 2728 6808
rect 13924 6792 13952 6820
rect 15545 6817 15557 6820
rect 15591 6817 15603 6851
rect 15545 6811 15603 6817
rect 19242 6808 19248 6860
rect 19300 6848 19306 6860
rect 19300 6820 19345 6848
rect 19300 6808 19306 6820
rect 23198 6808 23204 6860
rect 23256 6848 23262 6860
rect 23477 6851 23535 6857
rect 23477 6848 23489 6851
rect 23256 6820 23489 6848
rect 23256 6808 23262 6820
rect 23477 6817 23489 6820
rect 23523 6817 23535 6851
rect 23477 6811 23535 6817
rect 24121 6851 24179 6857
rect 24121 6817 24133 6851
rect 24167 6848 24179 6851
rect 24210 6848 24216 6860
rect 24167 6820 24216 6848
rect 24167 6817 24179 6820
rect 24121 6811 24179 6817
rect 24210 6808 24216 6820
rect 24268 6808 24274 6860
rect 26510 6848 26516 6860
rect 26423 6820 26516 6848
rect 26510 6808 26516 6820
rect 26568 6848 26574 6860
rect 27338 6848 27344 6860
rect 26568 6820 27344 6848
rect 26568 6808 26574 6820
rect 27338 6808 27344 6820
rect 27396 6808 27402 6860
rect 6914 6780 6920 6792
rect 2455 6752 2728 6780
rect 6875 6752 6920 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6749 7067 6783
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 7009 6743 7067 6749
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2648 6684 2697 6712
rect 2648 6672 2654 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 6546 6672 6552 6724
rect 6604 6712 6610 6724
rect 7024 6712 7052 6743
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6780 10379 6783
rect 10410 6780 10416 6792
rect 10367 6752 10416 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 11882 6780 11888 6792
rect 11843 6752 11888 6780
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 13814 6780 13820 6792
rect 13775 6752 13820 6780
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 13964 6752 14009 6780
rect 13964 6740 13970 6752
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 15286 6780 15292 6792
rect 15068 6752 15292 6780
rect 15068 6740 15074 6752
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 19426 6780 19432 6792
rect 19387 6752 19432 6780
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 23566 6780 23572 6792
rect 23527 6752 23572 6780
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 6604 6684 7052 6712
rect 9677 6715 9735 6721
rect 6604 6672 6610 6684
rect 9677 6681 9689 6715
rect 9723 6712 9735 6715
rect 9766 6712 9772 6724
rect 9723 6684 9772 6712
rect 9723 6681 9735 6684
rect 9677 6675 9735 6681
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 12621 6715 12679 6721
rect 12621 6681 12633 6715
rect 12667 6712 12679 6715
rect 13354 6712 13360 6724
rect 12667 6684 13360 6712
rect 12667 6681 12679 6684
rect 12621 6675 12679 6681
rect 13354 6672 13360 6684
rect 13412 6672 13418 6724
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 1946 6644 1952 6656
rect 1907 6616 1952 6644
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 3878 6644 3884 6656
rect 3191 6616 3884 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 6457 6647 6515 6653
rect 6457 6613 6469 6647
rect 6503 6644 6515 6647
rect 6730 6644 6736 6656
rect 6503 6616 6736 6644
rect 6503 6613 6515 6616
rect 6457 6607 6515 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 7469 6647 7527 6653
rect 7469 6644 7481 6647
rect 7432 6616 7481 6644
rect 7432 6604 7438 6616
rect 7469 6613 7481 6616
rect 7515 6613 7527 6647
rect 7469 6607 7527 6613
rect 12989 6647 13047 6653
rect 12989 6613 13001 6647
rect 13035 6644 13047 6647
rect 13078 6644 13084 6656
rect 13035 6616 13084 6644
rect 13035 6613 13047 6616
rect 12989 6607 13047 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 15304 6644 15332 6740
rect 26694 6712 26700 6724
rect 26655 6684 26700 6712
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 16482 6644 16488 6656
rect 15304 6616 16488 6644
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 16666 6644 16672 6656
rect 16627 6616 16672 6644
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 18785 6647 18843 6653
rect 18785 6644 18797 6647
rect 18564 6616 18797 6644
rect 18564 6604 18570 6616
rect 18785 6613 18797 6616
rect 18831 6613 18843 6647
rect 25222 6644 25228 6656
rect 25183 6616 25228 6644
rect 18785 6607 18843 6613
rect 25222 6604 25228 6616
rect 25280 6604 25286 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2130 6440 2136 6452
rect 2087 6412 2136 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 2130 6400 2136 6412
rect 2188 6400 2194 6452
rect 2409 6443 2467 6449
rect 2409 6409 2421 6443
rect 2455 6440 2467 6443
rect 2866 6440 2872 6452
rect 2455 6412 2872 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 2516 6245 2544 6412
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 5813 6443 5871 6449
rect 5813 6409 5825 6443
rect 5859 6440 5871 6443
rect 6822 6440 6828 6452
rect 5859 6412 6828 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6972 6412 7021 6440
rect 6972 6400 6978 6412
rect 7009 6409 7021 6412
rect 7055 6409 7067 6443
rect 7009 6403 7067 6409
rect 8849 6443 8907 6449
rect 8849 6409 8861 6443
rect 8895 6440 8907 6443
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 8895 6412 10057 6440
rect 8895 6409 8907 6412
rect 8849 6403 8907 6409
rect 10045 6409 10057 6412
rect 10091 6440 10103 6443
rect 10134 6440 10140 6452
rect 10091 6412 10140 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11790 6440 11796 6452
rect 11379 6412 11796 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 11977 6443 12035 6449
rect 11977 6440 11989 6443
rect 11940 6412 11989 6440
rect 11940 6400 11946 6412
rect 11977 6409 11989 6412
rect 12023 6409 12035 6443
rect 11977 6403 12035 6409
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 13964 6412 14289 6440
rect 13964 6400 13970 6412
rect 14277 6409 14289 6412
rect 14323 6440 14335 6443
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 14323 6412 14841 6440
rect 14323 6409 14335 6412
rect 14277 6403 14335 6409
rect 14829 6409 14841 6412
rect 14875 6409 14887 6443
rect 14829 6403 14887 6409
rect 15746 6400 15752 6452
rect 15804 6440 15810 6452
rect 16482 6440 16488 6452
rect 15804 6412 16488 6440
rect 15804 6400 15810 6412
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 19150 6440 19156 6452
rect 19111 6412 19156 6440
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 19300 6412 19441 6440
rect 19300 6400 19306 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 22741 6443 22799 6449
rect 22741 6409 22753 6443
rect 22787 6440 22799 6443
rect 23290 6440 23296 6452
rect 22787 6412 23296 6440
rect 22787 6409 22799 6412
rect 22741 6403 22799 6409
rect 23290 6400 23296 6412
rect 23348 6400 23354 6452
rect 23474 6400 23480 6452
rect 23532 6440 23538 6452
rect 23661 6443 23719 6449
rect 23661 6440 23673 6443
rect 23532 6412 23673 6440
rect 23532 6400 23538 6412
rect 23661 6409 23673 6412
rect 23707 6409 23719 6443
rect 27338 6440 27344 6452
rect 27299 6412 27344 6440
rect 23661 6403 23719 6409
rect 27338 6400 27344 6412
rect 27396 6400 27402 6452
rect 6546 6372 6552 6384
rect 6507 6344 6552 6372
rect 6546 6332 6552 6344
rect 6604 6332 6610 6384
rect 10410 6372 10416 6384
rect 9140 6344 10416 6372
rect 7006 6264 7012 6316
rect 7064 6304 7070 6316
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7064 6276 7573 6304
rect 7064 6264 7070 6276
rect 7561 6273 7573 6276
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6205 2559 6239
rect 2501 6199 2559 6205
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3234 6236 3240 6248
rect 3191 6208 3240 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 3973 6239 4031 6245
rect 3973 6236 3985 6239
rect 3712 6208 3985 6236
rect 1946 6128 1952 6180
rect 2004 6168 2010 6180
rect 3421 6171 3479 6177
rect 3421 6168 3433 6171
rect 2004 6140 3433 6168
rect 2004 6128 2010 6140
rect 3421 6137 3433 6140
rect 3467 6168 3479 6171
rect 3712 6168 3740 6208
rect 3973 6205 3985 6208
rect 4019 6205 4031 6239
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 3973 6199 4031 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7576 6236 7604 6267
rect 9140 6245 9168 6344
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 9582 6304 9588 6316
rect 9495 6276 9588 6304
rect 9582 6264 9588 6276
rect 9640 6304 9646 6316
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 9640 6276 10701 6304
rect 9640 6264 9646 6276
rect 10689 6273 10701 6276
rect 10735 6304 10747 6307
rect 11330 6304 11336 6316
rect 10735 6276 11336 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 11330 6264 11336 6276
rect 11388 6304 11394 6316
rect 11900 6304 11928 6400
rect 17865 6375 17923 6381
rect 17865 6341 17877 6375
rect 17911 6372 17923 6375
rect 22373 6375 22431 6381
rect 17911 6344 18644 6372
rect 17911 6341 17923 6344
rect 17865 6335 17923 6341
rect 18616 6316 18644 6344
rect 22373 6341 22385 6375
rect 22419 6372 22431 6375
rect 23566 6372 23572 6384
rect 22419 6344 23572 6372
rect 22419 6341 22431 6344
rect 22373 6335 22431 6341
rect 23566 6332 23572 6344
rect 23624 6372 23630 6384
rect 24118 6372 24124 6384
rect 23624 6344 24124 6372
rect 23624 6332 23630 6344
rect 24118 6332 24124 6344
rect 24176 6372 24182 6384
rect 24673 6375 24731 6381
rect 24673 6372 24685 6375
rect 24176 6344 24685 6372
rect 24176 6332 24182 6344
rect 13354 6304 13360 6316
rect 11388 6276 11928 6304
rect 13315 6276 13360 6304
rect 11388 6264 11394 6276
rect 13354 6264 13360 6276
rect 13412 6264 13418 6316
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 7576 6208 9137 6236
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9858 6236 9864 6248
rect 9819 6208 9864 6236
rect 9125 6199 9183 6205
rect 9858 6196 9864 6208
rect 9916 6236 9922 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 9916 6208 10425 6236
rect 9916 6196 9922 6208
rect 10413 6205 10425 6208
rect 10459 6205 10471 6239
rect 10413 6199 10471 6205
rect 13078 6196 13084 6248
rect 13136 6236 13142 6248
rect 13464 6236 13492 6267
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 13909 6307 13967 6313
rect 13909 6304 13921 6307
rect 13872 6276 13921 6304
rect 13872 6264 13878 6276
rect 13909 6273 13921 6276
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 15194 6264 15200 6316
rect 15252 6304 15258 6316
rect 16301 6307 16359 6313
rect 16301 6304 16313 6307
rect 15252 6276 16313 6304
rect 15252 6264 15258 6276
rect 16301 6273 16313 6276
rect 16347 6304 16359 6307
rect 16666 6304 16672 6316
rect 16347 6276 16672 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 16666 6264 16672 6276
rect 16724 6304 16730 6316
rect 16761 6307 16819 6313
rect 16761 6304 16773 6307
rect 16724 6276 16773 6304
rect 16724 6264 16730 6276
rect 16761 6273 16773 6276
rect 16807 6273 16819 6307
rect 18506 6304 18512 6316
rect 18467 6276 18512 6304
rect 16761 6267 16819 6273
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 19610 6304 19616 6316
rect 18656 6276 18749 6304
rect 19571 6276 19616 6304
rect 18656 6264 18662 6276
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 23109 6307 23167 6313
rect 23109 6273 23121 6307
rect 23155 6304 23167 6307
rect 23198 6304 23204 6316
rect 23155 6276 23204 6304
rect 23155 6273 23167 6276
rect 23109 6267 23167 6273
rect 23198 6264 23204 6276
rect 23256 6264 23262 6316
rect 24228 6313 24256 6344
rect 24673 6341 24685 6344
rect 24719 6372 24731 6375
rect 25222 6372 25228 6384
rect 24719 6344 25228 6372
rect 24719 6341 24731 6344
rect 24673 6335 24731 6341
rect 25222 6332 25228 6344
rect 25280 6332 25286 6384
rect 26602 6372 26608 6384
rect 26563 6344 26608 6372
rect 26602 6332 26608 6344
rect 26660 6332 26666 6384
rect 24213 6307 24271 6313
rect 24213 6273 24225 6307
rect 24259 6273 24271 6307
rect 24213 6267 24271 6273
rect 15562 6236 15568 6248
rect 13136 6208 13492 6236
rect 15523 6208 15568 6236
rect 13136 6196 13142 6208
rect 15562 6196 15568 6208
rect 15620 6236 15626 6248
rect 16209 6239 16267 6245
rect 16209 6236 16221 6239
rect 15620 6208 16221 6236
rect 15620 6196 15626 6208
rect 16209 6205 16221 6208
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 17497 6239 17555 6245
rect 17497 6205 17509 6239
rect 17543 6236 17555 6239
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 17543 6208 18429 6236
rect 17543 6205 17555 6208
rect 17497 6199 17555 6205
rect 18417 6205 18429 6208
rect 18463 6236 18475 6239
rect 18690 6236 18696 6248
rect 18463 6208 18696 6236
rect 18463 6205 18475 6208
rect 18417 6199 18475 6205
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 19426 6196 19432 6248
rect 19484 6196 19490 6248
rect 23474 6236 23480 6248
rect 23387 6208 23480 6236
rect 23474 6196 23480 6208
rect 23532 6236 23538 6248
rect 24121 6239 24179 6245
rect 24121 6236 24133 6239
rect 23532 6208 24133 6236
rect 23532 6196 23538 6208
rect 24121 6205 24133 6208
rect 24167 6236 24179 6239
rect 24762 6236 24768 6248
rect 24167 6208 24768 6236
rect 24167 6205 24179 6208
rect 24121 6199 24179 6205
rect 24762 6196 24768 6208
rect 24820 6196 24826 6248
rect 26418 6236 26424 6248
rect 26379 6208 26424 6236
rect 26418 6196 26424 6208
rect 26476 6236 26482 6248
rect 26973 6239 27031 6245
rect 26973 6236 26985 6239
rect 26476 6208 26985 6236
rect 26476 6196 26482 6208
rect 26973 6205 26985 6208
rect 27019 6205 27031 6239
rect 26973 6199 27031 6205
rect 3878 6168 3884 6180
rect 3467 6140 3740 6168
rect 3791 6140 3884 6168
rect 3467 6137 3479 6140
rect 3421 6131 3479 6137
rect 3878 6128 3884 6140
rect 3936 6168 3942 6180
rect 4240 6171 4298 6177
rect 4240 6168 4252 6171
rect 3936 6140 4252 6168
rect 3936 6128 3942 6140
rect 4240 6137 4252 6140
rect 4286 6168 4298 6171
rect 4982 6168 4988 6180
rect 4286 6140 4988 6168
rect 4286 6137 4298 6140
rect 4240 6131 4298 6137
rect 4982 6128 4988 6140
rect 5040 6128 5046 6180
rect 6181 6171 6239 6177
rect 6181 6137 6193 6171
rect 6227 6168 6239 6171
rect 7469 6171 7527 6177
rect 7469 6168 7481 6171
rect 6227 6140 7481 6168
rect 6227 6137 6239 6140
rect 6181 6131 6239 6137
rect 7469 6137 7481 6140
rect 7515 6168 7527 6171
rect 7558 6168 7564 6180
rect 7515 6140 7564 6168
rect 7515 6137 7527 6140
rect 7469 6131 7527 6137
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 10042 6128 10048 6180
rect 10100 6168 10106 6180
rect 10502 6168 10508 6180
rect 10100 6140 10508 6168
rect 10100 6128 10106 6140
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 12802 6168 12808 6180
rect 12715 6140 12808 6168
rect 12802 6128 12808 6140
rect 12860 6168 12866 6180
rect 15289 6171 15347 6177
rect 12860 6140 13308 6168
rect 12860 6128 12866 6140
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2498 6060 2504 6112
rect 2556 6100 2562 6112
rect 2685 6103 2743 6109
rect 2685 6100 2697 6103
rect 2556 6072 2697 6100
rect 2556 6060 2562 6072
rect 2685 6069 2697 6072
rect 2731 6069 2743 6103
rect 5350 6100 5356 6112
rect 5311 6072 5356 6100
rect 2685 6063 2743 6069
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 11606 6100 11612 6112
rect 11567 6072 11612 6100
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 12894 6100 12900 6112
rect 12855 6072 12900 6100
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13280 6109 13308 6140
rect 15289 6137 15301 6171
rect 15335 6168 15347 6171
rect 15838 6168 15844 6180
rect 15335 6140 15844 6168
rect 15335 6137 15347 6140
rect 15289 6131 15347 6137
rect 15838 6128 15844 6140
rect 15896 6168 15902 6180
rect 16117 6171 16175 6177
rect 16117 6168 16129 6171
rect 15896 6140 16129 6168
rect 15896 6128 15902 6140
rect 16117 6137 16129 6140
rect 16163 6137 16175 6171
rect 19444 6168 19472 6196
rect 19858 6171 19916 6177
rect 19858 6168 19870 6171
rect 19444 6140 19870 6168
rect 16117 6131 16175 6137
rect 19858 6137 19870 6140
rect 19904 6137 19916 6171
rect 19858 6131 19916 6137
rect 24029 6171 24087 6177
rect 24029 6137 24041 6171
rect 24075 6168 24087 6171
rect 24210 6168 24216 6180
rect 24075 6140 24216 6168
rect 24075 6137 24087 6140
rect 24029 6131 24087 6137
rect 24210 6128 24216 6140
rect 24268 6128 24274 6180
rect 13265 6103 13323 6109
rect 13265 6069 13277 6103
rect 13311 6100 13323 6103
rect 13354 6100 13360 6112
rect 13311 6072 13360 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 15746 6100 15752 6112
rect 15707 6072 15752 6100
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 17954 6060 17960 6112
rect 18012 6100 18018 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 18012 6072 18061 6100
rect 18012 6060 18018 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 20806 6060 20812 6112
rect 20864 6100 20870 6112
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 20864 6072 21005 6100
rect 20864 6060 20870 6072
rect 20993 6069 21005 6072
rect 21039 6069 21051 6103
rect 20993 6063 21051 6069
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1452 5868 1593 5896
rect 1452 5856 1458 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 2317 5899 2375 5905
rect 2317 5865 2329 5899
rect 2363 5896 2375 5899
rect 2406 5896 2412 5908
rect 2363 5868 2412 5896
rect 2363 5865 2375 5868
rect 2317 5859 2375 5865
rect 2406 5856 2412 5868
rect 2464 5896 2470 5908
rect 2777 5899 2835 5905
rect 2777 5896 2789 5899
rect 2464 5868 2789 5896
rect 2464 5856 2470 5868
rect 2777 5865 2789 5868
rect 2823 5865 2835 5899
rect 2777 5859 2835 5865
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 2915 5868 4077 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 6914 5896 6920 5908
rect 6595 5868 6920 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 2884 5828 2912 5859
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7006 5856 7012 5908
rect 7064 5896 7070 5908
rect 7064 5868 7109 5896
rect 7064 5856 7070 5868
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7745 5899 7803 5905
rect 7745 5896 7757 5899
rect 7432 5868 7757 5896
rect 7432 5856 7438 5868
rect 7745 5865 7757 5868
rect 7791 5865 7803 5899
rect 7745 5859 7803 5865
rect 8018 5856 8024 5908
rect 8076 5896 8082 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 8076 5868 8125 5896
rect 8076 5856 8082 5868
rect 8113 5865 8125 5868
rect 8159 5865 8171 5899
rect 8113 5859 8171 5865
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 9582 5896 9588 5908
rect 9539 5868 9588 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 10229 5899 10287 5905
rect 10229 5865 10241 5899
rect 10275 5896 10287 5899
rect 11606 5896 11612 5908
rect 10275 5868 11612 5896
rect 10275 5865 10287 5868
rect 10229 5859 10287 5865
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 12250 5896 12256 5908
rect 12211 5868 12256 5896
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12897 5899 12955 5905
rect 12897 5865 12909 5899
rect 12943 5896 12955 5899
rect 13170 5896 13176 5908
rect 12943 5868 13176 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 13170 5856 13176 5868
rect 13228 5856 13234 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15712 5868 15761 5896
rect 15712 5856 15718 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 15749 5859 15807 5865
rect 18141 5899 18199 5905
rect 18141 5865 18153 5899
rect 18187 5896 18199 5899
rect 18506 5896 18512 5908
rect 18187 5868 18512 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 19426 5896 19432 5908
rect 19387 5868 19432 5896
rect 19426 5856 19432 5868
rect 19484 5896 19490 5908
rect 19797 5899 19855 5905
rect 19797 5896 19809 5899
rect 19484 5868 19809 5896
rect 19484 5856 19490 5868
rect 19797 5865 19809 5868
rect 19843 5865 19855 5899
rect 24118 5896 24124 5908
rect 24079 5868 24124 5896
rect 19797 5859 19855 5865
rect 24118 5856 24124 5868
rect 24176 5856 24182 5908
rect 2740 5800 2912 5828
rect 2740 5788 2746 5800
rect 17954 5788 17960 5840
rect 18012 5828 18018 5840
rect 18785 5831 18843 5837
rect 18785 5828 18797 5831
rect 18012 5800 18797 5828
rect 18012 5788 18018 5800
rect 18785 5797 18797 5800
rect 18831 5797 18843 5831
rect 18785 5791 18843 5797
rect 22738 5788 22744 5840
rect 22796 5828 22802 5840
rect 22986 5831 23044 5837
rect 22986 5828 22998 5831
rect 22796 5800 22998 5828
rect 22796 5788 22802 5800
rect 22986 5797 22998 5800
rect 23032 5797 23044 5831
rect 22986 5791 23044 5797
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4212 5732 4445 5760
rect 4212 5720 4218 5732
rect 4433 5729 4445 5732
rect 4479 5760 4491 5763
rect 5442 5760 5448 5772
rect 4479 5732 5448 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 12802 5760 12808 5772
rect 12763 5732 12808 5760
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 15252 5732 15669 5760
rect 15252 5720 15258 5732
rect 15657 5729 15669 5732
rect 15703 5760 15715 5763
rect 15746 5760 15752 5772
rect 15703 5732 15752 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 21358 5720 21364 5772
rect 21416 5760 21422 5772
rect 23382 5760 23388 5772
rect 21416 5732 23388 5760
rect 21416 5720 21422 5732
rect 2406 5652 2412 5704
rect 2464 5692 2470 5704
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2464 5664 3065 5692
rect 2464 5652 2470 5664
rect 3053 5661 3065 5664
rect 3099 5692 3111 5695
rect 4522 5692 4528 5704
rect 3099 5664 4384 5692
rect 4483 5664 4528 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 4356 5624 4384 5664
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4982 5692 4988 5704
rect 4755 5664 4988 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7926 5692 7932 5704
rect 7064 5664 7932 5692
rect 7064 5652 7070 5664
rect 7926 5652 7932 5664
rect 7984 5692 7990 5704
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 7984 5664 8217 5692
rect 7984 5652 7990 5664
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 9490 5692 9496 5704
rect 8435 5664 9496 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 5350 5624 5356 5636
rect 4356 5596 5356 5624
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 7653 5627 7711 5633
rect 7653 5593 7665 5627
rect 7699 5624 7711 5627
rect 8404 5624 8432 5655
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 13078 5692 13084 5704
rect 13039 5664 13084 5692
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 15378 5652 15384 5704
rect 15436 5692 15442 5704
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 15436 5664 15853 5692
rect 15436 5652 15442 5664
rect 15841 5661 15853 5664
rect 15887 5661 15899 5695
rect 18874 5692 18880 5704
rect 18835 5664 18880 5692
rect 15841 5655 15899 5661
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 19058 5692 19064 5704
rect 19019 5664 19064 5692
rect 19058 5652 19064 5664
rect 19116 5652 19122 5704
rect 22756 5701 22784 5732
rect 23382 5720 23388 5732
rect 23440 5760 23446 5772
rect 24670 5760 24676 5772
rect 23440 5732 24676 5760
rect 23440 5720 23446 5732
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 26513 5763 26571 5769
rect 26513 5729 26525 5763
rect 26559 5760 26571 5763
rect 27062 5760 27068 5772
rect 26559 5732 27068 5760
rect 26559 5729 26571 5732
rect 26513 5723 26571 5729
rect 27062 5720 27068 5732
rect 27120 5720 27126 5772
rect 22741 5695 22799 5701
rect 22741 5661 22753 5695
rect 22787 5661 22799 5695
rect 22741 5655 22799 5661
rect 26694 5624 26700 5636
rect 7699 5596 8432 5624
rect 26655 5596 26700 5624
rect 7699 5593 7711 5596
rect 7653 5587 7711 5593
rect 26694 5584 26700 5596
rect 26752 5584 26758 5636
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 2590 5556 2596 5568
rect 2455 5528 2596 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 12437 5559 12495 5565
rect 12437 5525 12449 5559
rect 12483 5556 12495 5559
rect 12986 5556 12992 5568
rect 12483 5528 12992 5556
rect 12483 5525 12495 5528
rect 12437 5519 12495 5525
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 13446 5556 13452 5568
rect 13407 5528 13452 5556
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 15010 5556 15016 5568
rect 14608 5528 15016 5556
rect 14608 5516 14614 5528
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 18417 5559 18475 5565
rect 18417 5525 18429 5559
rect 18463 5556 18475 5559
rect 19150 5556 19156 5568
rect 18463 5528 19156 5556
rect 18463 5525 18475 5528
rect 18417 5519 18475 5525
rect 19150 5516 19156 5528
rect 19208 5516 19214 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 2406 5352 2412 5364
rect 2367 5324 2412 5352
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 4062 5352 4068 5364
rect 4019 5324 4068 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4982 5352 4988 5364
rect 4943 5324 4988 5352
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 5721 5355 5779 5361
rect 5721 5352 5733 5355
rect 5500 5324 5733 5352
rect 5500 5312 5506 5324
rect 5721 5321 5733 5324
rect 5767 5321 5779 5355
rect 7558 5352 7564 5364
rect 7519 5324 7564 5352
rect 5721 5315 5779 5321
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 8570 5352 8576 5364
rect 8076 5324 8576 5352
rect 8076 5312 8082 5324
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 9033 5355 9091 5361
rect 9033 5321 9045 5355
rect 9079 5352 9091 5355
rect 9490 5352 9496 5364
rect 9079 5324 9496 5352
rect 9079 5321 9091 5324
rect 9033 5315 9091 5321
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3513 5219 3571 5225
rect 3513 5216 3525 5219
rect 3108 5188 3525 5216
rect 3108 5176 3114 5188
rect 3513 5185 3525 5188
rect 3559 5216 3571 5219
rect 3970 5216 3976 5228
rect 3559 5188 3976 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3970 5176 3976 5188
rect 4028 5216 4034 5228
rect 4614 5216 4620 5228
rect 4028 5188 4620 5216
rect 4028 5176 4034 5188
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5216 8263 5219
rect 9048 5216 9076 5315
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 12158 5352 12164 5364
rect 12119 5324 12164 5352
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 15013 5355 15071 5361
rect 15013 5321 15025 5355
rect 15059 5352 15071 5355
rect 15194 5352 15200 5364
rect 15059 5324 15200 5352
rect 15059 5321 15071 5324
rect 15013 5315 15071 5321
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 15378 5352 15384 5364
rect 15339 5324 15384 5352
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 15654 5352 15660 5364
rect 15615 5324 15660 5352
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 17862 5352 17868 5364
rect 17823 5324 17868 5352
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 18874 5352 18880 5364
rect 18835 5324 18880 5352
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 22738 5352 22744 5364
rect 22699 5324 22744 5352
rect 22738 5312 22744 5324
rect 22796 5352 22802 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22796 5324 23029 5352
rect 22796 5312 22802 5324
rect 23017 5321 23029 5324
rect 23063 5321 23075 5355
rect 23382 5352 23388 5364
rect 23343 5324 23388 5352
rect 23017 5315 23075 5321
rect 23382 5312 23388 5324
rect 23440 5312 23446 5364
rect 27062 5312 27068 5364
rect 27120 5352 27126 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 27120 5324 27353 5352
rect 27120 5312 27126 5324
rect 27341 5321 27353 5324
rect 27387 5321 27399 5355
rect 27341 5315 27399 5321
rect 13817 5287 13875 5293
rect 13817 5253 13829 5287
rect 13863 5284 13875 5287
rect 14366 5284 14372 5296
rect 13863 5256 14372 5284
rect 13863 5253 13875 5256
rect 13817 5247 13875 5253
rect 14366 5244 14372 5256
rect 14424 5284 14430 5296
rect 15396 5284 15424 5312
rect 14424 5256 15424 5284
rect 18509 5287 18567 5293
rect 14424 5244 14430 5256
rect 18509 5253 18521 5287
rect 18555 5284 18567 5287
rect 19058 5284 19064 5296
rect 18555 5256 19064 5284
rect 18555 5253 18567 5256
rect 18509 5247 18567 5253
rect 19058 5244 19064 5256
rect 19116 5244 19122 5296
rect 8251 5188 9076 5216
rect 8251 5185 8263 5188
rect 8205 5179 8263 5185
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 12308 5188 12449 5216
rect 12308 5176 12314 5188
rect 12437 5185 12449 5188
rect 12483 5185 12495 5219
rect 12437 5179 12495 5185
rect 15838 5176 15844 5228
rect 15896 5216 15902 5228
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 15896 5188 15945 5216
rect 15896 5176 15902 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 18598 5176 18604 5228
rect 18656 5216 18662 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 18656 5188 19441 5216
rect 18656 5176 18662 5188
rect 19429 5185 19441 5188
rect 19475 5216 19487 5219
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 19475 5188 19901 5216
rect 19475 5185 19487 5188
rect 19429 5179 19487 5185
rect 19889 5185 19901 5188
rect 19935 5216 19947 5219
rect 20806 5216 20812 5228
rect 19935 5188 20812 5216
rect 19935 5185 19947 5188
rect 19889 5179 19947 5185
rect 20806 5176 20812 5188
rect 20864 5216 20870 5228
rect 21177 5219 21235 5225
rect 21177 5216 21189 5219
rect 20864 5188 21189 5216
rect 20864 5176 20870 5188
rect 21177 5185 21189 5188
rect 21223 5185 21235 5219
rect 21177 5179 21235 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 3881 5151 3939 5157
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 3927 5120 4353 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 4341 5117 4353 5120
rect 4387 5148 4399 5151
rect 5074 5148 5080 5160
rect 4387 5120 5080 5148
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 1412 5080 1440 5111
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 19058 5108 19064 5160
rect 19116 5148 19122 5160
rect 19337 5151 19395 5157
rect 19337 5148 19349 5151
rect 19116 5120 19349 5148
rect 19116 5108 19122 5120
rect 19337 5117 19349 5120
rect 19383 5148 19395 5151
rect 20257 5151 20315 5157
rect 20257 5148 20269 5151
rect 19383 5120 20269 5148
rect 19383 5117 19395 5120
rect 19337 5111 19395 5117
rect 20257 5117 20269 5120
rect 20303 5117 20315 5151
rect 20257 5111 20315 5117
rect 2038 5080 2044 5092
rect 1412 5052 2044 5080
rect 2038 5040 2044 5052
rect 2096 5040 2102 5092
rect 3145 5083 3203 5089
rect 3145 5049 3157 5083
rect 3191 5080 3203 5083
rect 4430 5080 4436 5092
rect 3191 5052 4436 5080
rect 3191 5049 3203 5052
rect 3145 5043 3203 5049
rect 4430 5040 4436 5052
rect 4488 5040 4494 5092
rect 4522 5040 4528 5092
rect 4580 5080 4586 5092
rect 5353 5083 5411 5089
rect 5353 5080 5365 5083
rect 4580 5052 5365 5080
rect 4580 5040 4586 5052
rect 5353 5049 5365 5052
rect 5399 5049 5411 5083
rect 8018 5080 8024 5092
rect 7931 5052 8024 5080
rect 5353 5043 5411 5049
rect 8018 5040 8024 5052
rect 8076 5080 8082 5092
rect 9309 5083 9367 5089
rect 9309 5080 9321 5083
rect 8076 5052 9321 5080
rect 8076 5040 8082 5052
rect 9309 5049 9321 5052
rect 9355 5049 9367 5083
rect 9309 5043 9367 5049
rect 11885 5083 11943 5089
rect 11885 5049 11897 5083
rect 11931 5080 11943 5083
rect 12682 5083 12740 5089
rect 12682 5080 12694 5083
rect 11931 5052 12694 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 12682 5049 12694 5052
rect 12728 5080 12740 5083
rect 13078 5080 13084 5092
rect 12728 5052 13084 5080
rect 12728 5049 12740 5052
rect 12682 5043 12740 5049
rect 13078 5040 13084 5052
rect 13136 5080 13142 5092
rect 14093 5083 14151 5089
rect 14093 5080 14105 5083
rect 13136 5052 14105 5080
rect 13136 5040 13142 5052
rect 14093 5049 14105 5052
rect 14139 5080 14151 5083
rect 15102 5080 15108 5092
rect 14139 5052 15108 5080
rect 14139 5049 14151 5052
rect 14093 5043 14151 5049
rect 15102 5040 15108 5052
rect 15160 5040 15166 5092
rect 19242 5080 19248 5092
rect 19155 5052 19248 5080
rect 19242 5040 19248 5052
rect 19300 5080 19306 5092
rect 20717 5083 20775 5089
rect 20717 5080 20729 5083
rect 19300 5052 20729 5080
rect 19300 5040 19306 5052
rect 20717 5049 20729 5052
rect 20763 5049 20775 5083
rect 21192 5080 21220 5179
rect 21358 5148 21364 5160
rect 21319 5120 21364 5148
rect 21358 5108 21364 5120
rect 21416 5108 21422 5160
rect 26418 5148 26424 5160
rect 26379 5120 26424 5148
rect 26418 5108 26424 5120
rect 26476 5148 26482 5160
rect 26973 5151 27031 5157
rect 26973 5148 26985 5151
rect 26476 5120 26985 5148
rect 26476 5108 26482 5120
rect 26973 5117 26985 5120
rect 27019 5117 27031 5151
rect 26973 5111 27031 5117
rect 21606 5083 21664 5089
rect 21606 5080 21618 5083
rect 21192 5052 21618 5080
rect 20717 5043 20775 5049
rect 21606 5049 21618 5052
rect 21652 5049 21664 5083
rect 21606 5043 21664 5049
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 7006 5012 7012 5024
rect 6967 4984 7012 5012
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7469 5015 7527 5021
rect 7469 4981 7481 5015
rect 7515 5012 7527 5015
rect 7929 5015 7987 5021
rect 7929 5012 7941 5015
rect 7515 4984 7941 5012
rect 7515 4981 7527 4984
rect 7469 4975 7527 4981
rect 7929 4981 7941 4984
rect 7975 5012 7987 5015
rect 8202 5012 8208 5024
rect 7975 4984 8208 5012
rect 7975 4981 7987 4984
rect 7929 4975 7987 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 26602 5012 26608 5024
rect 26563 4984 26608 5012
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 2501 4811 2559 4817
rect 2501 4777 2513 4811
rect 2547 4808 2559 4811
rect 2682 4808 2688 4820
rect 2547 4780 2688 4808
rect 2547 4777 2559 4780
rect 2501 4771 2559 4777
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 4065 4811 4123 4817
rect 4065 4777 4077 4811
rect 4111 4808 4123 4811
rect 4522 4808 4528 4820
rect 4111 4780 4528 4808
rect 4111 4777 4123 4780
rect 4065 4771 4123 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 11057 4811 11115 4817
rect 11057 4777 11069 4811
rect 11103 4808 11115 4811
rect 11330 4808 11336 4820
rect 11103 4780 11336 4808
rect 11103 4777 11115 4780
rect 11057 4771 11115 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 12526 4808 12532 4820
rect 12487 4780 12532 4808
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 12621 4811 12679 4817
rect 12621 4777 12633 4811
rect 12667 4777 12679 4811
rect 12621 4771 12679 4777
rect 2041 4743 2099 4749
rect 2041 4740 2053 4743
rect 1412 4712 2053 4740
rect 1412 4681 1440 4712
rect 2041 4709 2053 4712
rect 2087 4740 2099 4743
rect 2866 4740 2872 4752
rect 2087 4712 2872 4740
rect 2087 4709 2099 4712
rect 2041 4703 2099 4709
rect 2866 4700 2872 4712
rect 2924 4700 2930 4752
rect 10134 4740 10140 4752
rect 9692 4712 10140 4740
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4641 1455 4675
rect 1397 4635 1455 4641
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4672 2835 4675
rect 3234 4672 3240 4684
rect 2823 4644 3240 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 3878 4632 3884 4684
rect 3936 4672 3942 4684
rect 7098 4681 7104 4684
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 3936 4644 4445 4672
rect 3936 4632 3942 4644
rect 4433 4641 4445 4644
rect 4479 4641 4491 4675
rect 7092 4672 7104 4681
rect 7059 4644 7104 4672
rect 4433 4635 4491 4641
rect 7092 4635 7104 4644
rect 7098 4632 7104 4635
rect 7156 4632 7162 4684
rect 9692 4681 9720 4712
rect 10134 4700 10140 4712
rect 10192 4700 10198 4752
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 9933 4675 9991 4681
rect 9933 4672 9945 4675
rect 9824 4644 9945 4672
rect 9824 4632 9830 4644
rect 9933 4641 9945 4644
rect 9979 4641 9991 4675
rect 12636 4672 12664 4771
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 12952 4780 13093 4808
rect 12952 4768 12958 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15344 4780 15669 4808
rect 15344 4768 15350 4780
rect 15657 4777 15669 4780
rect 15703 4808 15715 4811
rect 15838 4808 15844 4820
rect 15703 4780 15844 4808
rect 15703 4777 15715 4780
rect 15657 4771 15715 4777
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 18509 4811 18567 4817
rect 18509 4777 18521 4811
rect 18555 4808 18567 4811
rect 18874 4808 18880 4820
rect 18555 4780 18880 4808
rect 18555 4777 18567 4780
rect 18509 4771 18567 4777
rect 18874 4768 18880 4780
rect 18932 4768 18938 4820
rect 19242 4808 19248 4820
rect 19203 4780 19248 4808
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 19613 4811 19671 4817
rect 19613 4777 19625 4811
rect 19659 4808 19671 4811
rect 19886 4808 19892 4820
rect 19659 4780 19892 4808
rect 19659 4777 19671 4780
rect 19613 4771 19671 4777
rect 19886 4768 19892 4780
rect 19944 4768 19950 4820
rect 21358 4808 21364 4820
rect 21319 4780 21364 4808
rect 21358 4768 21364 4780
rect 21416 4768 21422 4820
rect 12986 4740 12992 4752
rect 12947 4712 12992 4740
rect 12986 4700 12992 4712
rect 13044 4700 13050 4752
rect 19153 4743 19211 4749
rect 19153 4709 19165 4743
rect 19199 4740 19211 4743
rect 19426 4740 19432 4752
rect 19199 4712 19432 4740
rect 19199 4709 19211 4712
rect 19153 4703 19211 4709
rect 19426 4700 19432 4712
rect 19484 4740 19490 4752
rect 19484 4712 19748 4740
rect 19484 4700 19490 4712
rect 15746 4672 15752 4684
rect 12636 4644 15752 4672
rect 9933 4635 9991 4641
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 19720 4672 19748 4712
rect 26510 4672 26516 4684
rect 19720 4644 19840 4672
rect 26423 4644 26516 4672
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 4120 4576 4537 4604
rect 4120 4564 4126 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4614 4564 4620 4616
rect 4672 4604 4678 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4672 4576 4721 4604
rect 4672 4564 4678 4576
rect 4709 4573 4721 4576
rect 4755 4604 4767 4607
rect 5442 4604 5448 4616
rect 4755 4576 5448 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6604 4576 6837 4604
rect 6604 4564 6610 4576
rect 6825 4573 6837 4576
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 13265 4607 13323 4613
rect 13265 4604 13277 4607
rect 12768 4576 13277 4604
rect 12768 4564 12774 4576
rect 13265 4573 13277 4576
rect 13311 4604 13323 4607
rect 14366 4604 14372 4616
rect 13311 4576 14372 4604
rect 13311 4573 13323 4576
rect 13265 4567 13323 4573
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16298 4604 16304 4616
rect 15979 4576 16304 4604
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16298 4564 16304 4576
rect 16356 4564 16362 4616
rect 19242 4564 19248 4616
rect 19300 4604 19306 4616
rect 19812 4613 19840 4644
rect 26510 4632 26516 4644
rect 26568 4672 26574 4684
rect 27338 4672 27344 4684
rect 26568 4644 27344 4672
rect 26568 4632 26574 4644
rect 27338 4632 27344 4644
rect 27396 4632 27402 4684
rect 19705 4607 19763 4613
rect 19705 4604 19717 4607
rect 19300 4576 19717 4604
rect 19300 4564 19306 4576
rect 19705 4573 19717 4576
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 1486 4496 1492 4548
rect 1544 4536 1550 4548
rect 1946 4536 1952 4548
rect 1544 4508 1952 4536
rect 1544 4496 1550 4508
rect 1946 4496 1952 4508
rect 2004 4536 2010 4548
rect 3329 4539 3387 4545
rect 3329 4536 3341 4539
rect 2004 4508 3341 4536
rect 2004 4496 2010 4508
rect 3329 4505 3341 4508
rect 3375 4505 3387 4539
rect 3329 4499 3387 4505
rect 1394 4428 1400 4480
rect 1452 4468 1458 4480
rect 1581 4471 1639 4477
rect 1581 4468 1593 4471
rect 1452 4440 1593 4468
rect 1452 4428 1458 4440
rect 1581 4437 1593 4440
rect 1627 4437 1639 4471
rect 2958 4468 2964 4480
rect 2919 4440 2964 4468
rect 1581 4431 1639 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3878 4468 3884 4480
rect 3839 4440 3884 4468
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 8202 4468 8208 4480
rect 8163 4440 8208 4468
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 26694 4468 26700 4480
rect 26655 4440 26700 4468
rect 26694 4428 26700 4440
rect 26752 4428 26758 4480
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 2869 4267 2927 4273
rect 2869 4233 2881 4267
rect 2915 4264 2927 4267
rect 3050 4264 3056 4276
rect 2915 4236 3056 4264
rect 2915 4233 2927 4236
rect 2869 4227 2927 4233
rect 3050 4224 3056 4236
rect 3108 4224 3114 4276
rect 4157 4267 4215 4273
rect 4157 4233 4169 4267
rect 4203 4264 4215 4267
rect 4246 4264 4252 4276
rect 4203 4236 4252 4264
rect 4203 4233 4215 4236
rect 4157 4227 4215 4233
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 4617 4267 4675 4273
rect 4617 4264 4629 4267
rect 4488 4236 4629 4264
rect 4488 4224 4494 4236
rect 4617 4233 4629 4236
rect 4663 4233 4675 4267
rect 7098 4264 7104 4276
rect 7059 4236 7104 4264
rect 4617 4227 4675 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 8018 4264 8024 4276
rect 7979 4236 8024 4264
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 9766 4264 9772 4276
rect 9727 4236 9772 4264
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 10134 4264 10140 4276
rect 10095 4236 10140 4264
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 12710 4264 12716 4276
rect 12671 4236 12716 4264
rect 12710 4224 12716 4236
rect 12768 4224 12774 4276
rect 12894 4224 12900 4276
rect 12952 4264 12958 4276
rect 12989 4267 13047 4273
rect 12989 4264 13001 4267
rect 12952 4236 13001 4264
rect 12952 4224 12958 4236
rect 12989 4233 13001 4236
rect 13035 4233 13047 4267
rect 14366 4264 14372 4276
rect 14327 4236 14372 4264
rect 12989 4227 13047 4233
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 16209 4267 16267 4273
rect 16209 4264 16221 4267
rect 15804 4236 16221 4264
rect 15804 4224 15810 4236
rect 16209 4233 16221 4236
rect 16255 4233 16267 4267
rect 19058 4264 19064 4276
rect 19019 4236 19064 4264
rect 16209 4227 16267 4233
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 19886 4224 19892 4276
rect 19944 4264 19950 4276
rect 20073 4267 20131 4273
rect 20073 4264 20085 4267
rect 19944 4236 20085 4264
rect 19944 4224 19950 4236
rect 20073 4233 20085 4236
rect 20119 4233 20131 4267
rect 27338 4264 27344 4276
rect 27299 4236 27344 4264
rect 20073 4227 20131 4233
rect 27338 4224 27344 4236
rect 27396 4224 27402 4276
rect 7561 4199 7619 4205
rect 7561 4165 7573 4199
rect 7607 4196 7619 4199
rect 8202 4196 8208 4208
rect 7607 4168 8208 4196
rect 7607 4165 7619 4168
rect 7561 4159 7619 4165
rect 8202 4156 8208 4168
rect 8260 4196 8266 4208
rect 9784 4196 9812 4224
rect 8260 4168 9812 4196
rect 8260 4156 8266 4168
rect 4614 4088 4620 4140
rect 4672 4128 4678 4140
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4672 4100 5181 4128
rect 4672 4088 4678 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 8680 4137 8708 4168
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5500 4100 5641 4128
rect 5500 4088 5506 4100
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13357 4131 13415 4137
rect 13357 4128 13369 4131
rect 13044 4100 13369 4128
rect 13044 4088 13050 4100
rect 13357 4097 13369 4100
rect 13403 4097 13415 4131
rect 14384 4128 14412 4224
rect 15933 4199 15991 4205
rect 15933 4165 15945 4199
rect 15979 4196 15991 4199
rect 16298 4196 16304 4208
rect 15979 4168 16304 4196
rect 15979 4165 15991 4168
rect 15933 4159 15991 4165
rect 16298 4156 16304 4168
rect 16356 4156 16362 4208
rect 18601 4131 18659 4137
rect 14384 4100 14688 4128
rect 13357 4091 13415 4097
rect 1486 4060 1492 4072
rect 1447 4032 1492 4060
rect 1486 4020 1492 4032
rect 1544 4020 1550 4072
rect 3234 4060 3240 4072
rect 3195 4032 3240 4060
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 4246 4020 4252 4072
rect 4304 4060 4310 4072
rect 4985 4063 5043 4069
rect 4985 4060 4997 4063
rect 4304 4032 4997 4060
rect 4304 4020 4310 4032
rect 4985 4029 4997 4032
rect 5031 4029 5043 4063
rect 4985 4023 5043 4029
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4060 7987 4063
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 7975 4032 8493 4060
rect 7975 4029 7987 4032
rect 7929 4023 7987 4029
rect 8481 4029 8493 4032
rect 8527 4060 8539 4063
rect 9582 4060 9588 4072
rect 8527 4032 9588 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 14660 4060 14688 4100
rect 18601 4097 18613 4131
rect 18647 4128 18659 4131
rect 19242 4128 19248 4140
rect 18647 4100 19248 4128
rect 18647 4097 18659 4100
rect 18601 4091 18659 4097
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 19484 4100 19625 4128
rect 19484 4088 19490 4100
rect 19613 4097 19625 4100
rect 19659 4128 19671 4131
rect 20441 4131 20499 4137
rect 20441 4128 20453 4131
rect 19659 4100 20453 4128
rect 19659 4097 19671 4100
rect 19613 4091 19671 4097
rect 20441 4097 20453 4100
rect 20487 4097 20499 4131
rect 20441 4091 20499 4097
rect 14809 4063 14867 4069
rect 14809 4060 14821 4063
rect 14660 4032 14821 4060
rect 14809 4029 14821 4032
rect 14855 4029 14867 4063
rect 26418 4060 26424 4072
rect 26379 4032 26424 4060
rect 14809 4023 14867 4029
rect 26418 4020 26424 4032
rect 26476 4060 26482 4072
rect 26973 4063 27031 4069
rect 26973 4060 26985 4063
rect 26476 4032 26985 4060
rect 26476 4020 26482 4032
rect 26973 4029 26985 4032
rect 27019 4029 27031 4063
rect 27522 4060 27528 4072
rect 27483 4032 27528 4060
rect 26973 4023 27031 4029
rect 27522 4020 27528 4032
rect 27580 4060 27586 4072
rect 28077 4063 28135 4069
rect 28077 4060 28089 4063
rect 27580 4032 28089 4060
rect 27580 4020 27586 4032
rect 28077 4029 28089 4032
rect 28123 4029 28135 4063
rect 28077 4023 28135 4029
rect 1756 3995 1814 4001
rect 1756 3961 1768 3995
rect 1802 3992 1814 3995
rect 2314 3992 2320 4004
rect 1802 3964 2320 3992
rect 1802 3961 1814 3964
rect 1756 3955 1814 3961
rect 2314 3952 2320 3964
rect 2372 3992 2378 4004
rect 2774 3992 2780 4004
rect 2372 3964 2780 3992
rect 2372 3952 2378 3964
rect 2774 3952 2780 3964
rect 2832 3992 2838 4004
rect 3697 3995 3755 4001
rect 3697 3992 3709 3995
rect 2832 3964 3709 3992
rect 2832 3952 2838 3964
rect 3697 3961 3709 3964
rect 3743 3961 3755 3995
rect 8386 3992 8392 4004
rect 8347 3964 8392 3992
rect 3697 3955 3755 3961
rect 8386 3952 8392 3964
rect 8444 3952 8450 4004
rect 18966 3952 18972 4004
rect 19024 3992 19030 4004
rect 19521 3995 19579 4001
rect 19521 3992 19533 3995
rect 19024 3964 19533 3992
rect 19024 3952 19030 3964
rect 19521 3961 19533 3964
rect 19567 3992 19579 3995
rect 20809 3995 20867 4001
rect 20809 3992 20821 3995
rect 19567 3964 20821 3992
rect 19567 3961 19579 3964
rect 19521 3955 19579 3961
rect 20809 3961 20821 3964
rect 20855 3961 20867 3995
rect 20809 3955 20867 3961
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 5074 3924 5080 3936
rect 4571 3896 5080 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 6546 3924 6552 3936
rect 6507 3896 6552 3924
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 18874 3924 18880 3936
rect 18787 3896 18880 3924
rect 18874 3884 18880 3896
rect 18932 3924 18938 3936
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 18932 3896 19441 3924
rect 18932 3884 18938 3896
rect 19429 3893 19441 3896
rect 19475 3924 19487 3927
rect 19610 3924 19616 3936
rect 19475 3896 19616 3924
rect 19475 3893 19487 3896
rect 19429 3887 19487 3893
rect 19610 3884 19616 3896
rect 19668 3884 19674 3936
rect 26602 3924 26608 3936
rect 26563 3896 26608 3924
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 27706 3924 27712 3936
rect 27667 3896 27712 3924
rect 27706 3884 27712 3896
rect 27764 3884 27770 3936
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 2314 3720 2320 3732
rect 2275 3692 2320 3720
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 3142 3720 3148 3732
rect 3103 3692 3148 3720
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4062 3720 4068 3732
rect 3927 3692 4068 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 8113 3723 8171 3729
rect 8113 3689 8125 3723
rect 8159 3720 8171 3723
rect 8386 3720 8392 3732
rect 8159 3692 8392 3720
rect 8159 3689 8171 3692
rect 8113 3683 8171 3689
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 15838 3720 15844 3732
rect 15799 3692 15844 3720
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19889 3723 19947 3729
rect 19889 3720 19901 3723
rect 19484 3692 19901 3720
rect 19484 3680 19490 3692
rect 19889 3689 19901 3692
rect 19935 3689 19947 3723
rect 19889 3683 19947 3689
rect 2041 3655 2099 3661
rect 2041 3652 2053 3655
rect 1412 3624 2053 3652
rect 1412 3593 1440 3624
rect 2041 3621 2053 3624
rect 2087 3652 2099 3655
rect 4246 3652 4252 3664
rect 2087 3624 4252 3652
rect 2087 3621 2099 3624
rect 2041 3615 2099 3621
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 2498 3584 2504 3596
rect 2411 3556 2504 3584
rect 1397 3547 1455 3553
rect 2498 3544 2504 3556
rect 2556 3584 2562 3596
rect 4430 3584 4436 3596
rect 2556 3556 4436 3584
rect 2556 3544 2562 3556
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 5626 3584 5632 3596
rect 5587 3556 5632 3584
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 16298 3593 16304 3596
rect 15565 3587 15623 3593
rect 15565 3553 15577 3587
rect 15611 3584 15623 3587
rect 16292 3584 16304 3593
rect 15611 3556 16304 3584
rect 15611 3553 15623 3556
rect 15565 3547 15623 3553
rect 16292 3547 16304 3556
rect 16298 3544 16304 3547
rect 16356 3544 16362 3596
rect 17770 3544 17776 3596
rect 17828 3584 17834 3596
rect 18765 3587 18823 3593
rect 18765 3584 18777 3587
rect 17828 3556 18777 3584
rect 17828 3544 17834 3556
rect 18765 3553 18777 3556
rect 18811 3584 18823 3587
rect 19058 3584 19064 3596
rect 18811 3556 19064 3584
rect 18811 3553 18823 3556
rect 18765 3547 18823 3553
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 26510 3584 26516 3596
rect 26471 3556 26516 3584
rect 26510 3544 26516 3556
rect 26568 3544 26574 3596
rect 3694 3476 3700 3528
rect 3752 3516 3758 3528
rect 4338 3516 4344 3528
rect 3752 3488 4344 3516
rect 3752 3476 3758 3488
rect 4338 3476 4344 3488
rect 4396 3516 4402 3528
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 4396 3488 4537 3516
rect 4396 3476 4402 3488
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 5905 3519 5963 3525
rect 4672 3488 4717 3516
rect 4672 3476 4678 3488
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 7742 3516 7748 3528
rect 5951 3488 7748 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 14608 3488 14657 3516
rect 14608 3476 14614 3488
rect 14645 3485 14657 3488
rect 14691 3516 14703 3519
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 14691 3488 16037 3516
rect 14691 3485 14703 3488
rect 14645 3479 14703 3485
rect 16025 3485 16037 3488
rect 16071 3485 16083 3519
rect 18506 3516 18512 3528
rect 18467 3488 18512 3516
rect 16025 3479 16083 3485
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 16040 3380 16068 3479
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 16390 3380 16396 3392
rect 16040 3352 16396 3380
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 17405 3383 17463 3389
rect 17405 3349 17417 3383
rect 17451 3380 17463 3383
rect 17770 3380 17776 3392
rect 17451 3352 17776 3380
rect 17451 3349 17463 3352
rect 17405 3343 17463 3349
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 26697 3383 26755 3389
rect 26697 3349 26709 3383
rect 26743 3380 26755 3383
rect 26786 3380 26792 3392
rect 26743 3352 26792 3380
rect 26743 3349 26755 3352
rect 26697 3343 26755 3349
rect 26786 3340 26792 3352
rect 26844 3340 26850 3392
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 3936 3148 4077 3176
rect 3936 3136 3942 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 4065 3139 4123 3145
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5684 3148 6193 3176
rect 5684 3136 5690 3148
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 13262 3176 13268 3188
rect 13223 3148 13268 3176
rect 6181 3139 6239 3145
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 14458 3176 14464 3188
rect 14419 3148 14464 3176
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 16117 3179 16175 3185
rect 16117 3145 16129 3179
rect 16163 3176 16175 3179
rect 16298 3176 16304 3188
rect 16163 3148 16304 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 17770 3176 17776 3188
rect 17731 3148 17776 3176
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18782 3176 18788 3188
rect 18743 3148 18788 3176
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 18966 3176 18972 3188
rect 18927 3148 18972 3176
rect 18966 3136 18972 3148
rect 19024 3136 19030 3188
rect 21361 3179 21419 3185
rect 21361 3145 21373 3179
rect 21407 3176 21419 3179
rect 21542 3176 21548 3188
rect 21407 3148 21548 3176
rect 21407 3145 21419 3148
rect 21361 3139 21419 3145
rect 3973 3111 4031 3117
rect 3973 3077 3985 3111
rect 4019 3108 4031 3111
rect 4338 3108 4344 3120
rect 4019 3080 4344 3108
rect 4019 3077 4031 3080
rect 3973 3071 4031 3077
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 4430 3068 4436 3120
rect 4488 3108 4494 3120
rect 5169 3111 5227 3117
rect 5169 3108 5181 3111
rect 4488 3080 5181 3108
rect 4488 3068 4494 3080
rect 5169 3077 5181 3080
rect 5215 3108 5227 3111
rect 5718 3108 5724 3120
rect 5215 3080 5724 3108
rect 5215 3077 5227 3080
rect 5169 3071 5227 3077
rect 5718 3068 5724 3080
rect 5776 3068 5782 3120
rect 16390 3068 16396 3120
rect 16448 3108 16454 3120
rect 16485 3111 16543 3117
rect 16485 3108 16497 3111
rect 16448 3080 16497 3108
rect 16448 3068 16454 3080
rect 16485 3077 16497 3080
rect 16531 3108 16543 3111
rect 18506 3108 18512 3120
rect 16531 3080 18512 3108
rect 16531 3077 16543 3080
rect 16485 3071 16543 3077
rect 18506 3068 18512 3080
rect 18564 3108 18570 3120
rect 19981 3111 20039 3117
rect 19981 3108 19993 3111
rect 18564 3080 19993 3108
rect 18564 3068 18570 3080
rect 19981 3077 19993 3080
rect 20027 3077 20039 3111
rect 19981 3071 20039 3077
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 4614 3040 4620 3052
rect 2832 3012 4620 3040
rect 2832 3000 2838 3012
rect 4614 3000 4620 3012
rect 4672 3040 4678 3052
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 4672 3012 5457 3040
rect 4672 3000 4678 3012
rect 5445 3009 5457 3012
rect 5491 3040 5503 3043
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5491 3012 5825 3040
rect 5491 3009 5503 3012
rect 5445 3003 5503 3009
rect 5813 3009 5825 3012
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 19521 3043 19579 3049
rect 19521 3040 19533 3043
rect 19116 3012 19533 3040
rect 19116 3000 19122 3012
rect 19521 3009 19533 3012
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 3142 2972 3148 2984
rect 2731 2944 3148 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 1596 2904 1624 2935
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 4525 2975 4583 2981
rect 4525 2972 4537 2975
rect 3651 2944 4537 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 4525 2941 4537 2944
rect 4571 2972 4583 2975
rect 5166 2972 5172 2984
rect 4571 2944 5172 2972
rect 4571 2941 4583 2944
rect 4525 2935 4583 2941
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 8352 2944 8677 2972
rect 8352 2932 8358 2944
rect 8665 2941 8677 2944
rect 8711 2972 8723 2975
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 8711 2944 9413 2972
rect 8711 2941 8723 2944
rect 8665 2935 8723 2941
rect 9401 2941 9413 2944
rect 9447 2941 9459 2975
rect 9401 2935 9459 2941
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 13262 2972 13268 2984
rect 12483 2944 13268 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13725 2975 13783 2981
rect 13725 2941 13737 2975
rect 13771 2972 13783 2975
rect 14458 2972 14464 2984
rect 13771 2944 14464 2972
rect 13771 2941 13783 2944
rect 13725 2935 13783 2941
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 18012 2944 18521 2972
rect 18012 2932 18018 2944
rect 18509 2941 18521 2944
rect 18555 2972 18567 2975
rect 19337 2975 19395 2981
rect 19337 2972 19349 2975
rect 18555 2944 19349 2972
rect 18555 2941 18567 2944
rect 18509 2935 18567 2941
rect 19337 2941 19349 2944
rect 19383 2941 19395 2975
rect 19337 2935 19395 2941
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 20533 2975 20591 2981
rect 19484 2944 19529 2972
rect 19484 2932 19490 2944
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 21376 2972 21404 3139
rect 21542 3136 21548 3148
rect 21600 3136 21606 3188
rect 26510 3136 26516 3188
rect 26568 3176 26574 3188
rect 27249 3179 27307 3185
rect 27249 3176 27261 3179
rect 26568 3148 27261 3176
rect 26568 3136 26574 3148
rect 27249 3145 27261 3148
rect 27295 3145 27307 3179
rect 27249 3139 27307 3145
rect 23658 2972 23664 2984
rect 20579 2944 21404 2972
rect 23619 2944 23664 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 23658 2932 23664 2944
rect 23716 2972 23722 2984
rect 24397 2975 24455 2981
rect 24397 2972 24409 2975
rect 23716 2944 24409 2972
rect 23716 2932 23722 2944
rect 24397 2941 24409 2944
rect 24443 2941 24455 2975
rect 26326 2972 26332 2984
rect 26287 2944 26332 2972
rect 24397 2935 24455 2941
rect 26326 2932 26332 2944
rect 26384 2972 26390 2984
rect 26881 2975 26939 2981
rect 26881 2972 26893 2975
rect 26384 2944 26893 2972
rect 26384 2932 26390 2944
rect 26881 2941 26893 2944
rect 26927 2941 26939 2975
rect 27430 2972 27436 2984
rect 27391 2944 27436 2972
rect 26881 2935 26939 2941
rect 27430 2932 27436 2944
rect 27488 2972 27494 2984
rect 27985 2975 28043 2981
rect 27985 2972 27997 2975
rect 27488 2944 27997 2972
rect 27488 2932 27494 2944
rect 27985 2941 27997 2944
rect 28031 2941 28043 2975
rect 27985 2935 28043 2941
rect 2225 2907 2283 2913
rect 2225 2904 2237 2907
rect 1596 2876 2237 2904
rect 2225 2873 2237 2876
rect 2271 2904 2283 2907
rect 8941 2907 8999 2913
rect 2271 2876 4476 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 1762 2836 1768 2848
rect 1723 2808 1768 2836
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 2866 2836 2872 2848
rect 2827 2808 2872 2836
rect 2866 2796 2872 2808
rect 2924 2796 2930 2848
rect 4448 2845 4476 2876
rect 8941 2873 8953 2907
rect 8987 2904 8999 2907
rect 10594 2904 10600 2916
rect 8987 2876 10600 2904
rect 8987 2873 8999 2876
rect 8941 2867 8999 2873
rect 10594 2864 10600 2876
rect 10652 2864 10658 2916
rect 12713 2907 12771 2913
rect 12713 2873 12725 2907
rect 12759 2904 12771 2907
rect 13446 2904 13452 2916
rect 12759 2876 13452 2904
rect 12759 2873 12771 2876
rect 12713 2867 12771 2873
rect 13446 2864 13452 2876
rect 13504 2864 13510 2916
rect 14001 2907 14059 2913
rect 14001 2873 14013 2907
rect 14047 2904 14059 2907
rect 14918 2904 14924 2916
rect 14047 2876 14924 2904
rect 14047 2873 14059 2876
rect 14001 2867 14059 2873
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 18782 2864 18788 2916
rect 18840 2904 18846 2916
rect 19444 2904 19472 2932
rect 18840 2876 19472 2904
rect 18840 2864 18846 2876
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 20809 2907 20867 2913
rect 20809 2904 20821 2907
rect 20680 2876 20821 2904
rect 20680 2864 20686 2876
rect 20809 2873 20821 2876
rect 20855 2873 20867 2907
rect 20809 2867 20867 2873
rect 23937 2907 23995 2913
rect 23937 2873 23949 2907
rect 23983 2904 23995 2907
rect 24854 2904 24860 2916
rect 23983 2876 24860 2904
rect 23983 2873 23995 2876
rect 23937 2867 23995 2873
rect 24854 2864 24860 2876
rect 24912 2864 24918 2916
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2836 4491 2839
rect 5350 2836 5356 2848
rect 4479 2808 5356 2836
rect 4479 2805 4491 2808
rect 4433 2799 4491 2805
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 26510 2836 26516 2848
rect 26471 2808 26516 2836
rect 26510 2796 26516 2808
rect 26568 2796 26574 2848
rect 27614 2836 27620 2848
rect 27575 2808 27620 2836
rect 27614 2796 27620 2808
rect 27672 2796 27678 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 2590 2592 2596 2644
rect 2648 2632 2654 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 2648 2604 3801 2632
rect 2648 2592 2654 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5350 2632 5356 2644
rect 4939 2604 5356 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 1486 2496 1492 2508
rect 1447 2468 1492 2496
rect 1486 2456 1492 2468
rect 1544 2456 1550 2508
rect 1756 2499 1814 2505
rect 1756 2465 1768 2499
rect 1802 2496 1814 2499
rect 2038 2496 2044 2508
rect 1802 2468 2044 2496
rect 1802 2465 1814 2468
rect 1756 2459 1814 2465
rect 2038 2456 2044 2468
rect 2096 2496 2102 2508
rect 3145 2499 3203 2505
rect 3145 2496 3157 2499
rect 2096 2468 3157 2496
rect 2096 2456 2102 2468
rect 3145 2465 3157 2468
rect 3191 2465 3203 2499
rect 3804 2496 3832 2595
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 11514 2632 11520 2644
rect 11195 2604 11520 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 5810 2564 5816 2576
rect 5771 2536 5816 2564
rect 5810 2524 5816 2536
rect 5868 2524 5874 2576
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3804 2468 4077 2496
rect 3145 2459 3203 2465
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4982 2456 4988 2508
rect 5040 2496 5046 2508
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 5040 2468 5549 2496
rect 5040 2456 5046 2468
rect 5537 2465 5549 2468
rect 5583 2496 5595 2499
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5583 2468 6285 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 7653 2499 7711 2505
rect 7653 2496 7665 2499
rect 6972 2468 7665 2496
rect 6972 2456 6978 2468
rect 7653 2465 7665 2468
rect 7699 2465 7711 2499
rect 7653 2459 7711 2465
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 11164 2496 11192 2595
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 19058 2632 19064 2644
rect 19019 2604 19064 2632
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 21726 2592 21732 2644
rect 21784 2632 21790 2644
rect 21913 2635 21971 2641
rect 21913 2632 21925 2635
rect 21784 2604 21925 2632
rect 21784 2592 21790 2604
rect 21913 2601 21925 2604
rect 21959 2601 21971 2635
rect 21913 2595 21971 2601
rect 23477 2635 23535 2641
rect 23477 2601 23489 2635
rect 23523 2632 23535 2635
rect 24026 2632 24032 2644
rect 23523 2604 24032 2632
rect 23523 2601 23535 2604
rect 23477 2595 23535 2601
rect 13449 2567 13507 2573
rect 13449 2533 13461 2567
rect 13495 2564 13507 2567
rect 13722 2564 13728 2576
rect 13495 2536 13728 2564
rect 13495 2533 13507 2536
rect 13449 2527 13507 2533
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 10367 2468 11192 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12492 2468 13185 2496
rect 12492 2456 12498 2468
rect 13173 2465 13185 2468
rect 13219 2496 13231 2499
rect 13909 2499 13967 2505
rect 13909 2496 13921 2499
rect 13219 2468 13921 2496
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 13909 2465 13921 2468
rect 13955 2465 13967 2499
rect 13909 2459 13967 2465
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 15749 2499 15807 2505
rect 15749 2496 15761 2499
rect 15344 2468 15761 2496
rect 15344 2456 15350 2468
rect 15749 2465 15761 2468
rect 15795 2496 15807 2499
rect 16485 2499 16543 2505
rect 16485 2496 16497 2499
rect 15795 2468 16497 2496
rect 15795 2465 15807 2468
rect 15749 2459 15807 2465
rect 16485 2465 16497 2468
rect 16531 2465 16543 2499
rect 18064 2496 18092 2592
rect 18598 2564 18604 2576
rect 18559 2536 18604 2564
rect 18598 2524 18604 2536
rect 18656 2524 18662 2576
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18064 2468 18337 2496
rect 16485 2459 16543 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 19613 2499 19671 2505
rect 19613 2496 19625 2499
rect 19392 2468 19625 2496
rect 19392 2456 19398 2468
rect 19613 2465 19625 2468
rect 19659 2496 19671 2499
rect 20349 2499 20407 2505
rect 20349 2496 20361 2499
rect 19659 2468 20361 2496
rect 19659 2465 19671 2468
rect 19613 2459 19671 2465
rect 20349 2465 20361 2468
rect 20395 2465 20407 2499
rect 20349 2459 20407 2465
rect 21177 2499 21235 2505
rect 21177 2465 21189 2499
rect 21223 2496 21235 2499
rect 21744 2496 21772 2592
rect 21223 2468 21772 2496
rect 22649 2499 22707 2505
rect 21223 2465 21235 2468
rect 21177 2459 21235 2465
rect 22649 2465 22661 2499
rect 22695 2496 22707 2499
rect 23492 2496 23520 2595
rect 24026 2592 24032 2604
rect 24084 2592 24090 2644
rect 25682 2496 25688 2508
rect 22695 2468 23520 2496
rect 25595 2468 25688 2496
rect 22695 2465 22707 2468
rect 22649 2459 22707 2465
rect 25682 2456 25688 2468
rect 25740 2496 25746 2508
rect 26237 2499 26295 2505
rect 26237 2496 26249 2499
rect 25740 2468 26249 2496
rect 25740 2456 25746 2468
rect 26237 2465 26249 2468
rect 26283 2465 26295 2499
rect 26237 2459 26295 2465
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4890 2428 4896 2440
rect 4387 2400 4896 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6420 2400 7113 2428
rect 6420 2388 6426 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 12066 2428 12072 2440
rect 10643 2400 12072 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2428 16083 2431
rect 17770 2428 17776 2440
rect 16071 2400 17776 2428
rect 16071 2397 16083 2400
rect 16025 2391 16083 2397
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 19150 2388 19156 2440
rect 19208 2428 19214 2440
rect 19797 2431 19855 2437
rect 19797 2428 19809 2431
rect 19208 2400 19809 2428
rect 19208 2388 19214 2400
rect 19797 2397 19809 2400
rect 19843 2397 19855 2431
rect 19797 2391 19855 2397
rect 21453 2431 21511 2437
rect 21453 2397 21465 2431
rect 21499 2428 21511 2431
rect 22002 2428 22008 2440
rect 21499 2400 22008 2428
rect 21499 2397 21511 2400
rect 21453 2391 21511 2397
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23474 2428 23480 2440
rect 22971 2400 23480 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 2774 2320 2780 2372
rect 2832 2360 2838 2372
rect 2869 2363 2927 2369
rect 2869 2360 2881 2363
rect 2832 2332 2881 2360
rect 2832 2320 2838 2332
rect 2869 2329 2881 2332
rect 2915 2329 2927 2363
rect 2869 2323 2927 2329
rect 1486 2252 1492 2304
rect 1544 2292 1550 2304
rect 5169 2295 5227 2301
rect 5169 2292 5181 2295
rect 1544 2264 5181 2292
rect 1544 2252 1550 2264
rect 5169 2261 5181 2264
rect 5215 2292 5227 2295
rect 6546 2292 6552 2304
rect 5215 2264 6552 2292
rect 5215 2261 5227 2264
rect 5169 2255 5227 2261
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 25866 2292 25872 2304
rect 25827 2264 25872 2292
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 27065 2295 27123 2301
rect 27065 2261 27077 2295
rect 27111 2292 27123 2295
rect 29178 2292 29184 2304
rect 27111 2264 29184 2292
rect 27111 2261 27123 2264
rect 27065 2255 27123 2261
rect 29178 2252 29184 2264
rect 29236 2252 29242 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
rect 3510 552 3516 604
rect 3568 592 3574 604
rect 7282 592 7288 604
rect 3568 564 7288 592
rect 3568 552 3574 564
rect 7282 552 7288 564
rect 7340 552 7346 604
<< via1 >>
rect 3424 22176 3476 22228
rect 8300 22176 8352 22228
rect 3056 22108 3108 22160
rect 15660 22108 15712 22160
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 2964 20748 3016 20800
rect 17960 20748 18012 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 22468 20544 22520 20596
rect 25964 20247 26016 20256
rect 25964 20213 25973 20247
rect 25973 20213 26007 20247
rect 26007 20213 26016 20247
rect 25964 20204 26016 20213
rect 27804 20204 27856 20256
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 2596 19116 2648 19168
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 2136 18844 2188 18896
rect 3516 18844 3568 18896
rect 3608 18776 3660 18828
rect 9588 18776 9640 18828
rect 19156 18776 19208 18828
rect 22100 18776 22152 18828
rect 24492 18819 24544 18828
rect 2596 18751 2648 18760
rect 2596 18717 2605 18751
rect 2605 18717 2639 18751
rect 2639 18717 2648 18751
rect 2596 18708 2648 18717
rect 9772 18708 9824 18760
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 8208 18683 8260 18692
rect 8208 18649 8217 18683
rect 8217 18649 8251 18683
rect 8251 18649 8260 18683
rect 8208 18640 8260 18649
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 11704 18572 11756 18624
rect 12624 18615 12676 18624
rect 12624 18581 12633 18615
rect 12633 18581 12667 18615
rect 12667 18581 12676 18615
rect 12624 18572 12676 18581
rect 15292 18572 15344 18624
rect 19984 18615 20036 18624
rect 19984 18581 19993 18615
rect 19993 18581 20027 18615
rect 20027 18581 20036 18615
rect 19984 18572 20036 18581
rect 21088 18615 21140 18624
rect 21088 18581 21097 18615
rect 21097 18581 21131 18615
rect 21131 18581 21140 18615
rect 24492 18785 24526 18819
rect 24526 18785 24544 18819
rect 24492 18776 24544 18785
rect 21088 18572 21140 18581
rect 22192 18572 22244 18624
rect 24584 18572 24636 18624
rect 25596 18615 25648 18624
rect 25596 18581 25605 18615
rect 25605 18581 25639 18615
rect 25639 18581 25648 18615
rect 25596 18572 25648 18581
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 19984 18368 20036 18420
rect 20352 18368 20404 18420
rect 3516 18343 3568 18352
rect 3516 18309 3525 18343
rect 3525 18309 3559 18343
rect 3559 18309 3568 18343
rect 3516 18300 3568 18309
rect 15292 18300 15344 18352
rect 1768 18232 1820 18284
rect 2596 18275 2648 18284
rect 2596 18241 2605 18275
rect 2605 18241 2639 18275
rect 2639 18241 2648 18275
rect 2596 18232 2648 18241
rect 3608 18275 3660 18284
rect 3608 18241 3617 18275
rect 3617 18241 3651 18275
rect 3651 18241 3660 18275
rect 3608 18232 3660 18241
rect 11520 18232 11572 18284
rect 12624 18275 12676 18284
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 18604 18300 18656 18352
rect 19340 18300 19392 18352
rect 19156 18275 19208 18284
rect 19156 18241 19165 18275
rect 19165 18241 19199 18275
rect 19199 18241 19208 18275
rect 19156 18232 19208 18241
rect 3056 18164 3108 18216
rect 8208 18164 8260 18216
rect 12900 18207 12952 18216
rect 12900 18173 12923 18207
rect 12923 18173 12952 18207
rect 12900 18164 12952 18173
rect 18328 18164 18380 18216
rect 21088 18275 21140 18284
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 21088 18232 21140 18241
rect 24492 18232 24544 18284
rect 25044 18232 25096 18284
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 8576 18096 8628 18148
rect 9772 18096 9824 18148
rect 12164 18139 12216 18148
rect 12164 18105 12173 18139
rect 12173 18105 12207 18139
rect 12207 18105 12216 18139
rect 12164 18096 12216 18105
rect 14280 18096 14332 18148
rect 15476 18139 15528 18148
rect 15476 18105 15485 18139
rect 15485 18105 15519 18139
rect 15519 18105 15528 18139
rect 15476 18096 15528 18105
rect 19064 18139 19116 18148
rect 2596 18028 2648 18080
rect 3056 18071 3108 18080
rect 3056 18037 3065 18071
rect 3065 18037 3099 18071
rect 3099 18037 3108 18071
rect 3056 18028 3108 18037
rect 9588 18028 9640 18080
rect 15016 18071 15068 18080
rect 15016 18037 15025 18071
rect 15025 18037 15059 18071
rect 15059 18037 15068 18071
rect 15016 18028 15068 18037
rect 15200 18028 15252 18080
rect 16580 18028 16632 18080
rect 19064 18105 19073 18139
rect 19073 18105 19107 18139
rect 19107 18105 19116 18139
rect 19064 18096 19116 18105
rect 18328 18028 18380 18080
rect 18880 18028 18932 18080
rect 22100 18028 22152 18080
rect 24584 18071 24636 18080
rect 24584 18037 24593 18071
rect 24593 18037 24627 18071
rect 24627 18037 24636 18071
rect 25596 18096 25648 18148
rect 25136 18071 25188 18080
rect 24584 18028 24636 18037
rect 25136 18037 25145 18071
rect 25145 18037 25179 18071
rect 25179 18037 25188 18071
rect 25136 18028 25188 18037
rect 26240 18028 26292 18080
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 12900 17824 12952 17876
rect 14648 17824 14700 17876
rect 15016 17824 15068 17876
rect 18880 17756 18932 17808
rect 1768 17688 1820 17740
rect 4436 17688 4488 17740
rect 7748 17688 7800 17740
rect 11704 17688 11756 17740
rect 15200 17688 15252 17740
rect 18420 17688 18472 17740
rect 24216 17824 24268 17876
rect 22652 17688 22704 17740
rect 24952 17688 25004 17740
rect 1676 17663 1728 17672
rect 1676 17629 1685 17663
rect 1685 17629 1719 17663
rect 1719 17629 1728 17663
rect 1676 17620 1728 17629
rect 3792 17620 3844 17672
rect 7656 17620 7708 17672
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 9772 17620 9824 17672
rect 11520 17620 11572 17672
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 17592 17663 17644 17672
rect 17592 17629 17601 17663
rect 17601 17629 17635 17663
rect 17635 17629 17644 17663
rect 17592 17620 17644 17629
rect 19248 17663 19300 17672
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 21548 17663 21600 17672
rect 21548 17629 21557 17663
rect 21557 17629 21591 17663
rect 21591 17629 21600 17663
rect 21548 17620 21600 17629
rect 22008 17620 22060 17672
rect 25320 17663 25372 17672
rect 25320 17629 25329 17663
rect 25329 17629 25363 17663
rect 25363 17629 25372 17663
rect 25320 17620 25372 17629
rect 27160 17688 27212 17740
rect 26148 17620 26200 17672
rect 26792 17620 26844 17672
rect 9496 17552 9548 17604
rect 19156 17552 19208 17604
rect 22192 17552 22244 17604
rect 23572 17552 23624 17604
rect 24584 17552 24636 17604
rect 26332 17552 26384 17604
rect 2688 17484 2740 17536
rect 4436 17484 4488 17536
rect 5540 17484 5592 17536
rect 8576 17484 8628 17536
rect 10048 17527 10100 17536
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10048 17484 10100 17493
rect 10324 17527 10376 17536
rect 10324 17493 10333 17527
rect 10333 17493 10367 17527
rect 10367 17493 10376 17527
rect 10324 17484 10376 17493
rect 15108 17527 15160 17536
rect 15108 17493 15117 17527
rect 15117 17493 15151 17527
rect 15151 17493 15160 17527
rect 15108 17484 15160 17493
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 21456 17484 21508 17536
rect 24860 17527 24912 17536
rect 24860 17493 24869 17527
rect 24869 17493 24903 17527
rect 24903 17493 24912 17527
rect 24860 17484 24912 17493
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 1400 17280 1452 17332
rect 1676 17280 1728 17332
rect 3792 17323 3844 17332
rect 3792 17289 3801 17323
rect 3801 17289 3835 17323
rect 3835 17289 3844 17323
rect 3792 17280 3844 17289
rect 4436 17323 4488 17332
rect 4436 17289 4445 17323
rect 4445 17289 4479 17323
rect 4479 17289 4488 17323
rect 4436 17280 4488 17289
rect 7748 17323 7800 17332
rect 7748 17289 7757 17323
rect 7757 17289 7791 17323
rect 7791 17289 7800 17323
rect 7748 17280 7800 17289
rect 11520 17280 11572 17332
rect 18420 17323 18472 17332
rect 18420 17289 18429 17323
rect 18429 17289 18463 17323
rect 18463 17289 18472 17323
rect 18420 17280 18472 17289
rect 19248 17280 19300 17332
rect 20352 17323 20404 17332
rect 20352 17289 20361 17323
rect 20361 17289 20395 17323
rect 20395 17289 20404 17323
rect 20352 17280 20404 17289
rect 21364 17280 21416 17332
rect 22652 17323 22704 17332
rect 22652 17289 22661 17323
rect 22661 17289 22695 17323
rect 22695 17289 22704 17323
rect 22652 17280 22704 17289
rect 24216 17323 24268 17332
rect 24216 17289 24225 17323
rect 24225 17289 24259 17323
rect 24259 17289 24268 17323
rect 24216 17280 24268 17289
rect 25320 17280 25372 17332
rect 2044 17144 2096 17196
rect 5448 17212 5500 17264
rect 8484 17212 8536 17264
rect 2688 17187 2740 17196
rect 2688 17153 2697 17187
rect 2697 17153 2731 17187
rect 2731 17153 2740 17187
rect 2688 17144 2740 17153
rect 2964 17144 3016 17196
rect 5540 17187 5592 17196
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 10048 17144 10100 17196
rect 11704 17212 11756 17264
rect 13728 17212 13780 17264
rect 14924 17187 14976 17196
rect 14924 17153 14933 17187
rect 14933 17153 14967 17187
rect 14967 17153 14976 17187
rect 14924 17144 14976 17153
rect 15108 17144 15160 17196
rect 18144 17144 18196 17196
rect 18972 17144 19024 17196
rect 19156 17144 19208 17196
rect 19432 17144 19484 17196
rect 21548 17212 21600 17264
rect 24952 17255 25004 17264
rect 24952 17221 24961 17255
rect 24961 17221 24995 17255
rect 24995 17221 25004 17255
rect 24952 17212 25004 17221
rect 26792 17255 26844 17264
rect 26792 17221 26801 17255
rect 26801 17221 26835 17255
rect 26835 17221 26844 17255
rect 26792 17212 26844 17221
rect 26332 17187 26384 17196
rect 26332 17153 26341 17187
rect 26341 17153 26375 17187
rect 26375 17153 26384 17187
rect 26332 17144 26384 17153
rect 1952 17076 2004 17128
rect 8576 17119 8628 17128
rect 8576 17085 8585 17119
rect 8585 17085 8619 17119
rect 8619 17085 8628 17119
rect 8576 17076 8628 17085
rect 14648 17119 14700 17128
rect 14648 17085 14657 17119
rect 14657 17085 14691 17119
rect 14691 17085 14700 17119
rect 14648 17076 14700 17085
rect 21364 17119 21416 17128
rect 21364 17085 21373 17119
rect 21373 17085 21407 17119
rect 21407 17085 21416 17119
rect 21364 17076 21416 17085
rect 25136 17076 25188 17128
rect 5264 17051 5316 17060
rect 1768 16983 1820 16992
rect 1768 16949 1777 16983
rect 1777 16949 1811 16983
rect 1811 16949 1820 16983
rect 1768 16940 1820 16949
rect 5264 17017 5273 17051
rect 5273 17017 5307 17051
rect 5307 17017 5316 17051
rect 5264 17008 5316 17017
rect 10324 17051 10376 17060
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 4896 16940 4948 16949
rect 5356 16983 5408 16992
rect 5356 16949 5365 16983
rect 5365 16949 5399 16983
rect 5399 16949 5408 16983
rect 5356 16940 5408 16949
rect 7656 16940 7708 16992
rect 10324 17017 10333 17051
rect 10333 17017 10367 17051
rect 10367 17017 10376 17051
rect 10324 17008 10376 17017
rect 21272 17051 21324 17060
rect 21272 17017 21281 17051
rect 21281 17017 21315 17051
rect 21315 17017 21324 17051
rect 21272 17008 21324 17017
rect 26240 17051 26292 17060
rect 26240 17017 26249 17051
rect 26249 17017 26283 17051
rect 26283 17017 26292 17051
rect 26240 17008 26292 17017
rect 29184 17008 29236 17060
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 9588 16940 9640 16992
rect 10692 16940 10744 16992
rect 14740 16983 14792 16992
rect 14740 16949 14749 16983
rect 14749 16949 14783 16983
rect 14783 16949 14792 16983
rect 14740 16940 14792 16949
rect 15200 16940 15252 16992
rect 15384 16940 15436 16992
rect 16304 16940 16356 16992
rect 18788 16983 18840 16992
rect 18788 16949 18797 16983
rect 18797 16949 18831 16983
rect 18831 16949 18840 16983
rect 18788 16940 18840 16949
rect 26424 16940 26476 16992
rect 27160 16983 27212 16992
rect 27160 16949 27169 16983
rect 27169 16949 27203 16983
rect 27203 16949 27212 16983
rect 27160 16940 27212 16949
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 5356 16736 5408 16788
rect 8668 16736 8720 16788
rect 10048 16736 10100 16788
rect 11612 16779 11664 16788
rect 2688 16668 2740 16720
rect 5264 16711 5316 16720
rect 5264 16677 5273 16711
rect 5273 16677 5307 16711
rect 5307 16677 5316 16711
rect 5264 16668 5316 16677
rect 5540 16668 5592 16720
rect 9496 16711 9548 16720
rect 9496 16677 9505 16711
rect 9505 16677 9539 16711
rect 9539 16677 9548 16711
rect 9496 16668 9548 16677
rect 2412 16600 2464 16652
rect 4068 16600 4120 16652
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 2964 16575 3016 16584
rect 2964 16541 2973 16575
rect 2973 16541 3007 16575
rect 3007 16541 3016 16575
rect 2964 16532 3016 16541
rect 8116 16532 8168 16584
rect 8300 16600 8352 16652
rect 8668 16600 8720 16652
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 9128 16532 9180 16584
rect 11612 16745 11621 16779
rect 11621 16745 11655 16779
rect 11655 16745 11664 16779
rect 11612 16736 11664 16745
rect 14740 16736 14792 16788
rect 15660 16711 15712 16720
rect 15660 16677 15669 16711
rect 15669 16677 15703 16711
rect 15703 16677 15712 16711
rect 15660 16668 15712 16677
rect 11704 16643 11756 16652
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 11704 16600 11756 16609
rect 15936 16736 15988 16788
rect 17592 16736 17644 16788
rect 18788 16736 18840 16788
rect 18880 16779 18932 16788
rect 18880 16745 18889 16779
rect 18889 16745 18923 16779
rect 18923 16745 18932 16779
rect 18880 16736 18932 16745
rect 21272 16736 21324 16788
rect 27160 16736 27212 16788
rect 23480 16668 23532 16720
rect 24952 16668 25004 16720
rect 25412 16668 25464 16720
rect 9680 16532 9732 16584
rect 10324 16575 10376 16584
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 11980 16532 12032 16584
rect 15016 16532 15068 16584
rect 20812 16600 20864 16652
rect 21272 16600 21324 16652
rect 21640 16575 21692 16584
rect 1860 16464 1912 16516
rect 15200 16464 15252 16516
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 21548 16464 21600 16516
rect 21824 16532 21876 16584
rect 23572 16600 23624 16652
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 19708 16396 19760 16448
rect 26240 16464 26292 16516
rect 24676 16396 24728 16448
rect 27160 16396 27212 16448
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 1860 16235 1912 16244
rect 1860 16201 1869 16235
rect 1869 16201 1903 16235
rect 1903 16201 1912 16235
rect 1860 16192 1912 16201
rect 2688 16235 2740 16244
rect 2688 16201 2697 16235
rect 2697 16201 2731 16235
rect 2731 16201 2740 16235
rect 2688 16192 2740 16201
rect 4068 16235 4120 16244
rect 4068 16201 4077 16235
rect 4077 16201 4111 16235
rect 4111 16201 4120 16235
rect 4068 16192 4120 16201
rect 5540 16235 5592 16244
rect 5540 16201 5549 16235
rect 5549 16201 5583 16235
rect 5583 16201 5592 16235
rect 5540 16192 5592 16201
rect 8576 16192 8628 16244
rect 9496 16235 9548 16244
rect 1768 16124 1820 16176
rect 2964 16124 3016 16176
rect 5448 16124 5500 16176
rect 8668 16124 8720 16176
rect 9496 16201 9505 16235
rect 9505 16201 9539 16235
rect 9539 16201 9548 16235
rect 9496 16192 9548 16201
rect 10324 16192 10376 16244
rect 11612 16192 11664 16244
rect 15016 16235 15068 16244
rect 15016 16201 15025 16235
rect 15025 16201 15059 16235
rect 15059 16201 15068 16235
rect 15016 16192 15068 16201
rect 19432 16192 19484 16244
rect 20628 16235 20680 16244
rect 20628 16201 20637 16235
rect 20637 16201 20671 16235
rect 20671 16201 20680 16235
rect 20628 16192 20680 16201
rect 21364 16192 21416 16244
rect 23480 16235 23532 16244
rect 23480 16201 23489 16235
rect 23489 16201 23523 16235
rect 23523 16201 23532 16235
rect 23480 16192 23532 16201
rect 24952 16124 25004 16176
rect 25596 16124 25648 16176
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 11980 16099 12032 16108
rect 10508 16056 10560 16065
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 13360 16056 13412 16108
rect 3148 15988 3200 16040
rect 4988 15988 5040 16040
rect 10876 15988 10928 16040
rect 13544 15988 13596 16040
rect 21548 16056 21600 16108
rect 24216 16056 24268 16108
rect 24676 16099 24728 16108
rect 24676 16065 24685 16099
rect 24685 16065 24719 16099
rect 24719 16065 24728 16099
rect 24676 16056 24728 16065
rect 26332 16056 26384 16108
rect 27160 16056 27212 16108
rect 2872 15920 2924 15972
rect 3516 15920 3568 15972
rect 13728 15920 13780 15972
rect 15844 15988 15896 16040
rect 19340 15988 19392 16040
rect 24768 15988 24820 16040
rect 16304 15920 16356 15972
rect 3608 15852 3660 15904
rect 8116 15895 8168 15904
rect 8116 15861 8125 15895
rect 8125 15861 8159 15895
rect 8159 15861 8168 15895
rect 8116 15852 8168 15861
rect 8300 15852 8352 15904
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 11704 15895 11756 15904
rect 9956 15852 10008 15861
rect 11704 15861 11713 15895
rect 11713 15861 11747 15895
rect 11747 15861 11756 15895
rect 11704 15852 11756 15861
rect 13268 15895 13320 15904
rect 13268 15861 13277 15895
rect 13277 15861 13311 15895
rect 13311 15861 13320 15895
rect 13268 15852 13320 15861
rect 15660 15852 15712 15904
rect 17500 15920 17552 15972
rect 20720 15920 20772 15972
rect 21824 15963 21876 15972
rect 21824 15929 21833 15963
rect 21833 15929 21867 15963
rect 21867 15929 21876 15963
rect 21824 15920 21876 15929
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 21364 15852 21416 15904
rect 21916 15895 21968 15904
rect 21916 15861 21925 15895
rect 21925 15861 21959 15895
rect 21959 15861 21968 15895
rect 21916 15852 21968 15861
rect 22836 15895 22888 15904
rect 22836 15861 22845 15895
rect 22845 15861 22879 15895
rect 22879 15861 22888 15895
rect 22836 15852 22888 15861
rect 24032 15895 24084 15904
rect 24032 15861 24041 15895
rect 24041 15861 24075 15895
rect 24075 15861 24084 15895
rect 24032 15852 24084 15861
rect 24492 15895 24544 15904
rect 24492 15861 24501 15895
rect 24501 15861 24535 15895
rect 24535 15861 24544 15895
rect 24492 15852 24544 15861
rect 25136 15852 25188 15904
rect 25872 15920 25924 15972
rect 25596 15895 25648 15904
rect 25596 15861 25605 15895
rect 25605 15861 25639 15895
rect 25639 15861 25648 15895
rect 25596 15852 25648 15861
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 2412 15691 2464 15700
rect 2412 15657 2421 15691
rect 2421 15657 2455 15691
rect 2455 15657 2464 15691
rect 2412 15648 2464 15657
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 9956 15648 10008 15700
rect 10508 15648 10560 15700
rect 13360 15691 13412 15700
rect 13360 15657 13369 15691
rect 13369 15657 13403 15691
rect 13403 15657 13412 15691
rect 13360 15648 13412 15657
rect 15844 15691 15896 15700
rect 15844 15657 15853 15691
rect 15853 15657 15887 15691
rect 15887 15657 15896 15691
rect 15844 15648 15896 15657
rect 19340 15691 19392 15700
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 20628 15648 20680 15700
rect 21548 15691 21600 15700
rect 21548 15657 21557 15691
rect 21557 15657 21591 15691
rect 21591 15657 21600 15691
rect 21548 15648 21600 15657
rect 21640 15648 21692 15700
rect 22836 15648 22888 15700
rect 24492 15648 24544 15700
rect 25596 15648 25648 15700
rect 2780 15623 2832 15632
rect 2780 15589 2789 15623
rect 2789 15589 2823 15623
rect 2823 15589 2832 15623
rect 2780 15580 2832 15589
rect 4068 15580 4120 15632
rect 6276 15580 6328 15632
rect 6828 15580 6880 15632
rect 17132 15580 17184 15632
rect 24676 15580 24728 15632
rect 27068 15580 27120 15632
rect 2412 15512 2464 15564
rect 5448 15512 5500 15564
rect 9772 15512 9824 15564
rect 13728 15555 13780 15564
rect 13728 15521 13737 15555
rect 13737 15521 13771 15555
rect 13771 15521 13780 15555
rect 13728 15512 13780 15521
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 12992 15444 13044 15496
rect 12900 15376 12952 15428
rect 15844 15444 15896 15496
rect 16304 15487 16356 15496
rect 16304 15453 16313 15487
rect 16313 15453 16347 15487
rect 16347 15453 16356 15487
rect 16304 15444 16356 15453
rect 16764 15444 16816 15496
rect 19340 15512 19392 15564
rect 22652 15512 22704 15564
rect 24768 15512 24820 15564
rect 27252 15512 27304 15564
rect 21180 15444 21232 15496
rect 22284 15487 22336 15496
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 25412 15487 25464 15496
rect 22284 15444 22336 15453
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 25412 15444 25464 15453
rect 27160 15487 27212 15496
rect 27160 15453 27169 15487
rect 27169 15453 27203 15487
rect 27203 15453 27212 15487
rect 27160 15444 27212 15453
rect 1676 15351 1728 15360
rect 1676 15317 1685 15351
rect 1685 15317 1719 15351
rect 1719 15317 1728 15351
rect 3700 15351 3752 15360
rect 1676 15308 1728 15317
rect 3700 15317 3709 15351
rect 3709 15317 3743 15351
rect 3743 15317 3752 15351
rect 3700 15308 3752 15317
rect 7564 15351 7616 15360
rect 7564 15317 7573 15351
rect 7573 15317 7607 15351
rect 7607 15317 7616 15351
rect 7564 15308 7616 15317
rect 15200 15308 15252 15360
rect 18512 15351 18564 15360
rect 18512 15317 18521 15351
rect 18521 15317 18555 15351
rect 18555 15317 18564 15351
rect 18512 15308 18564 15317
rect 23572 15351 23624 15360
rect 23572 15317 23581 15351
rect 23581 15317 23615 15351
rect 23615 15317 23624 15351
rect 23572 15308 23624 15317
rect 24308 15308 24360 15360
rect 25044 15308 25096 15360
rect 26332 15308 26384 15360
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 2964 15104 3016 15156
rect 3608 15147 3660 15156
rect 3608 15113 3617 15147
rect 3617 15113 3651 15147
rect 3651 15113 3660 15147
rect 3608 15104 3660 15113
rect 4068 15104 4120 15156
rect 6276 15147 6328 15156
rect 6276 15113 6285 15147
rect 6285 15113 6319 15147
rect 6319 15113 6328 15147
rect 6276 15104 6328 15113
rect 9588 15104 9640 15156
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 12900 15147 12952 15156
rect 12900 15113 12909 15147
rect 12909 15113 12943 15147
rect 12943 15113 12952 15147
rect 12900 15104 12952 15113
rect 16764 15147 16816 15156
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 3700 14968 3752 15020
rect 4620 14968 4672 15020
rect 6644 15036 6696 15088
rect 6276 14968 6328 15020
rect 9312 15036 9364 15088
rect 9864 15036 9916 15088
rect 13728 15079 13780 15088
rect 13728 15045 13737 15079
rect 13737 15045 13771 15079
rect 13771 15045 13780 15079
rect 13728 15036 13780 15045
rect 16764 15113 16773 15147
rect 16773 15113 16807 15147
rect 16807 15113 16816 15147
rect 16764 15104 16816 15113
rect 17132 15147 17184 15156
rect 17132 15113 17141 15147
rect 17141 15113 17175 15147
rect 17175 15113 17184 15147
rect 17132 15104 17184 15113
rect 19892 15104 19944 15156
rect 21180 15147 21232 15156
rect 21180 15113 21189 15147
rect 21189 15113 21223 15147
rect 21223 15113 21232 15147
rect 21180 15104 21232 15113
rect 21916 15104 21968 15156
rect 22744 15147 22796 15156
rect 22744 15113 22753 15147
rect 22753 15113 22787 15147
rect 22787 15113 22796 15147
rect 22744 15104 22796 15113
rect 24676 15104 24728 15156
rect 25596 15104 25648 15156
rect 25872 15147 25924 15156
rect 25872 15113 25881 15147
rect 25881 15113 25915 15147
rect 25915 15113 25924 15147
rect 25872 15104 25924 15113
rect 25412 15036 25464 15088
rect 10232 14968 10284 15020
rect 12164 14968 12216 15020
rect 14188 14968 14240 15020
rect 15108 14968 15160 15020
rect 18512 14968 18564 15020
rect 19064 15011 19116 15020
rect 19064 14977 19073 15011
rect 19073 14977 19107 15011
rect 19107 14977 19116 15011
rect 19064 14968 19116 14977
rect 20720 14968 20772 15020
rect 21272 14968 21324 15020
rect 22284 15011 22336 15020
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 26332 14968 26384 15020
rect 1676 14943 1728 14952
rect 1676 14909 1710 14943
rect 1710 14909 1728 14943
rect 1676 14900 1728 14909
rect 5448 14900 5500 14952
rect 9404 14900 9456 14952
rect 10876 14900 10928 14952
rect 14556 14900 14608 14952
rect 18420 14943 18472 14952
rect 1124 14832 1176 14884
rect 7012 14832 7064 14884
rect 12992 14832 13044 14884
rect 18420 14909 18429 14943
rect 18429 14909 18463 14943
rect 18463 14909 18472 14943
rect 18420 14900 18472 14909
rect 18512 14875 18564 14884
rect 18512 14841 18521 14875
rect 18521 14841 18555 14875
rect 18555 14841 18564 14875
rect 18512 14832 18564 14841
rect 21732 14900 21784 14952
rect 21916 14832 21968 14884
rect 3700 14764 3752 14816
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 11336 14764 11388 14816
rect 13176 14764 13228 14816
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 17408 14807 17460 14816
rect 17408 14773 17417 14807
rect 17417 14773 17451 14807
rect 17451 14773 17460 14807
rect 17408 14764 17460 14773
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 20720 14807 20772 14816
rect 20720 14773 20729 14807
rect 20729 14773 20763 14807
rect 20763 14773 20772 14807
rect 20720 14764 20772 14773
rect 23112 14807 23164 14816
rect 23112 14773 23121 14807
rect 23121 14773 23155 14807
rect 23155 14773 23164 14807
rect 23112 14764 23164 14773
rect 25688 14807 25740 14816
rect 25688 14773 25697 14807
rect 25697 14773 25731 14807
rect 25731 14773 25740 14807
rect 25688 14764 25740 14773
rect 26608 14764 26660 14816
rect 27068 14764 27120 14816
rect 27252 14807 27304 14816
rect 27252 14773 27261 14807
rect 27261 14773 27295 14807
rect 27295 14773 27304 14807
rect 27252 14764 27304 14773
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 1676 14560 1728 14612
rect 2412 14603 2464 14612
rect 2412 14569 2421 14603
rect 2421 14569 2455 14603
rect 2455 14569 2464 14603
rect 2412 14560 2464 14569
rect 5172 14560 5224 14612
rect 6552 14560 6604 14612
rect 7196 14560 7248 14612
rect 9956 14560 10008 14612
rect 10600 14560 10652 14612
rect 11336 14560 11388 14612
rect 12992 14603 13044 14612
rect 12992 14569 13001 14603
rect 13001 14569 13035 14603
rect 13035 14569 13044 14603
rect 12992 14560 13044 14569
rect 15752 14560 15804 14612
rect 16304 14560 16356 14612
rect 17132 14560 17184 14612
rect 18052 14560 18104 14612
rect 19340 14603 19392 14612
rect 19340 14569 19349 14603
rect 19349 14569 19383 14603
rect 19383 14569 19392 14603
rect 19340 14560 19392 14569
rect 21824 14560 21876 14612
rect 27160 14560 27212 14612
rect 2872 14535 2924 14544
rect 2872 14501 2881 14535
rect 2881 14501 2915 14535
rect 2915 14501 2924 14535
rect 2872 14492 2924 14501
rect 4712 14492 4764 14544
rect 6828 14492 6880 14544
rect 13268 14492 13320 14544
rect 3608 14424 3660 14476
rect 5448 14424 5500 14476
rect 6276 14424 6328 14476
rect 9496 14467 9548 14476
rect 9496 14433 9505 14467
rect 9505 14433 9539 14467
rect 9539 14433 9548 14467
rect 9496 14424 9548 14433
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 12164 14424 12216 14476
rect 14004 14424 14056 14476
rect 18236 14467 18288 14476
rect 18236 14433 18245 14467
rect 18245 14433 18279 14467
rect 18279 14433 18288 14467
rect 18236 14424 18288 14433
rect 18696 14467 18748 14476
rect 18696 14433 18705 14467
rect 18705 14433 18739 14467
rect 18739 14433 18748 14467
rect 18696 14424 18748 14433
rect 21824 14424 21876 14476
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 3700 14399 3752 14408
rect 3700 14365 3709 14399
rect 3709 14365 3743 14399
rect 3743 14365 3752 14399
rect 3700 14356 3752 14365
rect 5632 14356 5684 14408
rect 7564 14356 7616 14408
rect 10140 14399 10192 14408
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 16856 14399 16908 14408
rect 1400 14220 1452 14272
rect 5540 14288 5592 14340
rect 5816 14288 5868 14340
rect 6460 14288 6512 14340
rect 9772 14288 9824 14340
rect 10324 14288 10376 14340
rect 16856 14365 16865 14399
rect 16865 14365 16899 14399
rect 16899 14365 16908 14399
rect 16856 14356 16908 14365
rect 18788 14399 18840 14408
rect 18788 14365 18797 14399
rect 18797 14365 18831 14399
rect 18831 14365 18840 14399
rect 18788 14356 18840 14365
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 22284 14399 22336 14408
rect 22284 14365 22293 14399
rect 22293 14365 22327 14399
rect 22327 14365 22336 14399
rect 22284 14356 22336 14365
rect 23112 14356 23164 14408
rect 19156 14288 19208 14340
rect 19340 14288 19392 14340
rect 22008 14288 22060 14340
rect 5080 14220 5132 14272
rect 5448 14263 5500 14272
rect 5448 14229 5457 14263
rect 5457 14229 5491 14263
rect 5491 14229 5500 14263
rect 5448 14220 5500 14229
rect 8116 14220 8168 14272
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 14096 14263 14148 14272
rect 14096 14229 14105 14263
rect 14105 14229 14139 14263
rect 14139 14229 14148 14263
rect 14096 14220 14148 14229
rect 15660 14220 15712 14272
rect 18328 14263 18380 14272
rect 18328 14229 18337 14263
rect 18337 14229 18371 14263
rect 18371 14229 18380 14263
rect 18328 14220 18380 14229
rect 24308 14263 24360 14272
rect 24308 14229 24317 14263
rect 24317 14229 24351 14263
rect 24351 14229 24360 14263
rect 24308 14220 24360 14229
rect 26608 14220 26660 14272
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 2412 14016 2464 14068
rect 2688 14016 2740 14068
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 8852 14059 8904 14068
rect 8852 14025 8861 14059
rect 8861 14025 8895 14059
rect 8895 14025 8904 14059
rect 8852 14016 8904 14025
rect 10048 14016 10100 14068
rect 10324 14059 10376 14068
rect 10324 14025 10333 14059
rect 10333 14025 10367 14059
rect 10367 14025 10376 14059
rect 10324 14016 10376 14025
rect 14096 14059 14148 14068
rect 14096 14025 14105 14059
rect 14105 14025 14139 14059
rect 14139 14025 14148 14059
rect 14096 14016 14148 14025
rect 16304 14059 16356 14068
rect 3608 13991 3660 14000
rect 3608 13957 3617 13991
rect 3617 13957 3651 13991
rect 3651 13957 3660 13991
rect 3608 13948 3660 13957
rect 2872 13880 2924 13932
rect 2964 13880 3016 13932
rect 5448 13880 5500 13932
rect 10232 13948 10284 14000
rect 12164 13991 12216 14000
rect 12164 13957 12173 13991
rect 12173 13957 12207 13991
rect 12207 13957 12216 13991
rect 12164 13948 12216 13957
rect 13820 13991 13872 14000
rect 13820 13957 13829 13991
rect 13829 13957 13863 13991
rect 13863 13957 13872 13991
rect 13820 13948 13872 13957
rect 15200 13948 15252 14000
rect 16304 14025 16313 14059
rect 16313 14025 16347 14059
rect 16347 14025 16356 14059
rect 16304 14016 16356 14025
rect 16672 14016 16724 14068
rect 17132 14059 17184 14068
rect 17132 14025 17141 14059
rect 17141 14025 17175 14059
rect 17175 14025 17184 14059
rect 17132 14016 17184 14025
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 16856 13948 16908 14000
rect 18880 13948 18932 14000
rect 21272 14059 21324 14068
rect 21272 14025 21281 14059
rect 21281 14025 21315 14059
rect 21315 14025 21324 14059
rect 21272 14016 21324 14025
rect 21824 14016 21876 14068
rect 24216 14059 24268 14068
rect 6368 13880 6420 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 2780 13812 2832 13864
rect 3240 13744 3292 13796
rect 5080 13744 5132 13796
rect 8116 13744 8168 13796
rect 15752 13923 15804 13932
rect 15752 13889 15761 13923
rect 15761 13889 15795 13923
rect 15795 13889 15804 13923
rect 15752 13880 15804 13889
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 18236 13880 18288 13932
rect 20720 13880 20772 13932
rect 22008 13880 22060 13932
rect 12532 13812 12584 13864
rect 15660 13855 15712 13864
rect 5172 13719 5224 13728
rect 5172 13685 5181 13719
rect 5181 13685 5215 13719
rect 5215 13685 5224 13719
rect 5172 13676 5224 13685
rect 5632 13676 5684 13728
rect 9036 13744 9088 13796
rect 11980 13744 12032 13796
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 18696 13812 18748 13864
rect 19156 13855 19208 13864
rect 19156 13821 19165 13855
rect 19165 13821 19199 13855
rect 19199 13821 19208 13855
rect 19156 13812 19208 13821
rect 21180 13812 21232 13864
rect 24216 14025 24225 14059
rect 24225 14025 24259 14059
rect 24259 14025 24268 14059
rect 24216 14016 24268 14025
rect 26884 13948 26936 14000
rect 23388 13812 23440 13864
rect 24308 13855 24360 13864
rect 16856 13744 16908 13796
rect 19064 13744 19116 13796
rect 19432 13787 19484 13796
rect 19432 13753 19444 13787
rect 19444 13753 19484 13787
rect 24308 13821 24317 13855
rect 24317 13821 24351 13855
rect 24351 13821 24360 13855
rect 24308 13812 24360 13821
rect 26516 13855 26568 13864
rect 26516 13821 26525 13855
rect 26525 13821 26559 13855
rect 26559 13821 26568 13855
rect 26516 13812 26568 13821
rect 19432 13744 19484 13753
rect 9588 13676 9640 13728
rect 21548 13676 21600 13728
rect 25872 13676 25924 13728
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 2964 13515 3016 13524
rect 2964 13481 2973 13515
rect 2973 13481 3007 13515
rect 3007 13481 3016 13515
rect 2964 13472 3016 13481
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 1492 13336 1544 13388
rect 2320 13336 2372 13388
rect 5632 13379 5684 13388
rect 5632 13345 5641 13379
rect 5641 13345 5675 13379
rect 5675 13345 5684 13379
rect 5632 13336 5684 13345
rect 7104 13336 7156 13388
rect 9496 13472 9548 13524
rect 13268 13472 13320 13524
rect 17224 13515 17276 13524
rect 17224 13481 17233 13515
rect 17233 13481 17267 13515
rect 17267 13481 17276 13515
rect 17224 13472 17276 13481
rect 18788 13472 18840 13524
rect 21364 13515 21416 13524
rect 21364 13481 21373 13515
rect 21373 13481 21407 13515
rect 21407 13481 21416 13515
rect 21364 13472 21416 13481
rect 23112 13515 23164 13524
rect 23112 13481 23121 13515
rect 23121 13481 23155 13515
rect 23155 13481 23164 13515
rect 23112 13472 23164 13481
rect 25228 13515 25280 13524
rect 25228 13481 25237 13515
rect 25237 13481 25271 13515
rect 25271 13481 25280 13515
rect 25228 13472 25280 13481
rect 12256 13447 12308 13456
rect 12256 13413 12290 13447
rect 12290 13413 12308 13447
rect 12256 13404 12308 13413
rect 16856 13404 16908 13456
rect 8484 13336 8536 13388
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 15476 13336 15528 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 25320 13404 25372 13456
rect 15752 13336 15804 13345
rect 5540 13268 5592 13320
rect 6276 13268 6328 13320
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 5356 13200 5408 13252
rect 17316 13311 17368 13320
rect 17316 13277 17325 13311
rect 17325 13277 17359 13311
rect 17359 13277 17368 13311
rect 17316 13268 17368 13277
rect 19524 13336 19576 13388
rect 21548 13336 21600 13388
rect 21824 13336 21876 13388
rect 19248 13311 19300 13320
rect 19248 13277 19257 13311
rect 19257 13277 19291 13311
rect 19291 13277 19300 13311
rect 19248 13268 19300 13277
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 25320 13311 25372 13320
rect 25320 13277 25329 13311
rect 25329 13277 25363 13311
rect 25363 13277 25372 13311
rect 25320 13268 25372 13277
rect 18696 13200 18748 13252
rect 25780 13200 25832 13252
rect 3240 13175 3292 13184
rect 3240 13141 3249 13175
rect 3249 13141 3283 13175
rect 3283 13141 3292 13175
rect 3240 13132 3292 13141
rect 5448 13132 5500 13184
rect 9036 13175 9088 13184
rect 9036 13141 9045 13175
rect 9045 13141 9079 13175
rect 9079 13141 9088 13175
rect 9036 13132 9088 13141
rect 10140 13132 10192 13184
rect 10784 13132 10836 13184
rect 13360 13175 13412 13184
rect 13360 13141 13369 13175
rect 13369 13141 13403 13175
rect 13403 13141 13412 13175
rect 13360 13132 13412 13141
rect 14280 13132 14332 13184
rect 24676 13132 24728 13184
rect 25872 13175 25924 13184
rect 25872 13141 25881 13175
rect 25881 13141 25915 13175
rect 25915 13141 25924 13175
rect 25872 13132 25924 13141
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 2136 12928 2188 12980
rect 2320 12971 2372 12980
rect 2320 12937 2329 12971
rect 2329 12937 2363 12971
rect 2363 12937 2372 12971
rect 2320 12928 2372 12937
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 5080 12928 5132 12980
rect 5724 12928 5776 12980
rect 4252 12860 4304 12912
rect 5632 12860 5684 12912
rect 6276 12928 6328 12980
rect 7104 12971 7156 12980
rect 7104 12937 7113 12971
rect 7113 12937 7147 12971
rect 7147 12937 7156 12971
rect 7104 12928 7156 12937
rect 9680 12928 9732 12980
rect 12256 12928 12308 12980
rect 13360 12928 13412 12980
rect 13728 12971 13780 12980
rect 13728 12937 13737 12971
rect 13737 12937 13771 12971
rect 13771 12937 13780 12971
rect 13728 12928 13780 12937
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 6460 12860 6512 12912
rect 11980 12860 12032 12912
rect 12808 12860 12860 12912
rect 15568 12860 15620 12912
rect 5448 12835 5500 12844
rect 5448 12801 5457 12835
rect 5457 12801 5491 12835
rect 5491 12801 5500 12835
rect 5448 12792 5500 12801
rect 5540 12835 5592 12844
rect 5540 12801 5549 12835
rect 5549 12801 5583 12835
rect 5583 12801 5592 12835
rect 5540 12792 5592 12801
rect 5724 12792 5776 12844
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 13728 12792 13780 12844
rect 16856 12928 16908 12980
rect 17316 12971 17368 12980
rect 17316 12937 17325 12971
rect 17325 12937 17359 12971
rect 17359 12937 17368 12971
rect 17316 12928 17368 12937
rect 18788 12971 18840 12980
rect 18788 12937 18797 12971
rect 18797 12937 18831 12971
rect 18831 12937 18840 12971
rect 18788 12928 18840 12937
rect 21824 12971 21876 12980
rect 21824 12937 21833 12971
rect 21833 12937 21867 12971
rect 21867 12937 21876 12971
rect 21824 12928 21876 12937
rect 25320 12971 25372 12980
rect 25320 12937 25329 12971
rect 25329 12937 25363 12971
rect 25363 12937 25372 12971
rect 25320 12928 25372 12937
rect 19524 12860 19576 12912
rect 21548 12860 21600 12912
rect 24308 12860 24360 12912
rect 17224 12792 17276 12844
rect 19432 12835 19484 12844
rect 19432 12801 19441 12835
rect 19441 12801 19475 12835
rect 19475 12801 19484 12835
rect 19432 12792 19484 12801
rect 23940 12792 23992 12844
rect 4804 12724 4856 12776
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 14372 12767 14424 12776
rect 14372 12733 14381 12767
rect 14381 12733 14415 12767
rect 14415 12733 14424 12767
rect 14372 12724 14424 12733
rect 15108 12724 15160 12776
rect 24400 12792 24452 12844
rect 24676 12767 24728 12776
rect 24676 12733 24685 12767
rect 24685 12733 24719 12767
rect 24719 12733 24728 12767
rect 25228 12860 25280 12912
rect 25320 12792 25372 12844
rect 25504 12792 25556 12844
rect 24676 12724 24728 12733
rect 1492 12656 1544 12708
rect 2688 12699 2740 12708
rect 2688 12665 2697 12699
rect 2697 12665 2731 12699
rect 2731 12665 2740 12699
rect 2688 12656 2740 12665
rect 7932 12656 7984 12708
rect 8484 12656 8536 12708
rect 9220 12656 9272 12708
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 9036 12588 9088 12640
rect 14464 12656 14516 12708
rect 15568 12656 15620 12708
rect 18972 12656 19024 12708
rect 25504 12656 25556 12708
rect 25872 12656 25924 12708
rect 26148 12656 26200 12708
rect 17960 12588 18012 12640
rect 24308 12588 24360 12640
rect 27160 12631 27212 12640
rect 27160 12597 27169 12631
rect 27169 12597 27203 12631
rect 27203 12597 27212 12631
rect 27160 12588 27212 12597
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 2320 12384 2372 12436
rect 6368 12427 6420 12436
rect 6368 12393 6377 12427
rect 6377 12393 6411 12427
rect 6411 12393 6420 12427
rect 6368 12384 6420 12393
rect 7748 12384 7800 12436
rect 7932 12384 7984 12436
rect 12808 12427 12860 12436
rect 12808 12393 12817 12427
rect 12817 12393 12851 12427
rect 12851 12393 12860 12427
rect 12808 12384 12860 12393
rect 14372 12384 14424 12436
rect 15568 12427 15620 12436
rect 15568 12393 15577 12427
rect 15577 12393 15611 12427
rect 15611 12393 15620 12427
rect 15568 12384 15620 12393
rect 15844 12384 15896 12436
rect 17684 12384 17736 12436
rect 18236 12384 18288 12436
rect 19432 12384 19484 12436
rect 23480 12384 23532 12436
rect 25044 12384 25096 12436
rect 25504 12427 25556 12436
rect 25504 12393 25513 12427
rect 25513 12393 25547 12427
rect 25547 12393 25556 12427
rect 25504 12384 25556 12393
rect 25596 12384 25648 12436
rect 26240 12427 26292 12436
rect 26240 12393 26249 12427
rect 26249 12393 26283 12427
rect 26283 12393 26292 12427
rect 26240 12384 26292 12393
rect 2780 12316 2832 12368
rect 15752 12316 15804 12368
rect 1492 12248 1544 12300
rect 1676 12291 1728 12300
rect 1676 12257 1710 12291
rect 1710 12257 1728 12291
rect 1676 12248 1728 12257
rect 2688 12248 2740 12300
rect 4988 12291 5040 12300
rect 4988 12257 4997 12291
rect 4997 12257 5031 12291
rect 5031 12257 5040 12291
rect 4988 12248 5040 12257
rect 5724 12248 5776 12300
rect 7840 12248 7892 12300
rect 10600 12248 10652 12300
rect 17776 12248 17828 12300
rect 18880 12248 18932 12300
rect 21548 12248 21600 12300
rect 21916 12291 21968 12300
rect 21916 12257 21950 12291
rect 21950 12257 21968 12291
rect 21916 12248 21968 12257
rect 24400 12248 24452 12300
rect 24768 12291 24820 12300
rect 24768 12257 24777 12291
rect 24777 12257 24811 12291
rect 24811 12257 24820 12291
rect 24768 12248 24820 12257
rect 7288 12180 7340 12232
rect 9036 12180 9088 12232
rect 9956 12180 10008 12232
rect 6276 12112 6328 12164
rect 9588 12112 9640 12164
rect 17868 12180 17920 12232
rect 25596 12180 25648 12232
rect 26884 12180 26936 12232
rect 24124 12112 24176 12164
rect 25688 12112 25740 12164
rect 26608 12112 26660 12164
rect 2780 12087 2832 12096
rect 2780 12053 2789 12087
rect 2789 12053 2823 12087
rect 2823 12053 2832 12087
rect 7932 12087 7984 12096
rect 2780 12044 2832 12053
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 8116 12044 8168 12096
rect 9680 12087 9732 12096
rect 9680 12053 9689 12087
rect 9689 12053 9723 12087
rect 9723 12053 9732 12087
rect 9680 12044 9732 12053
rect 16488 12087 16540 12096
rect 16488 12053 16497 12087
rect 16497 12053 16531 12087
rect 16531 12053 16540 12087
rect 16488 12044 16540 12053
rect 17132 12087 17184 12096
rect 17132 12053 17141 12087
rect 17141 12053 17175 12087
rect 17175 12053 17184 12087
rect 17132 12044 17184 12053
rect 19156 12044 19208 12096
rect 23020 12087 23072 12096
rect 23020 12053 23029 12087
rect 23029 12053 23063 12087
rect 23063 12053 23072 12087
rect 23020 12044 23072 12053
rect 24952 12044 25004 12096
rect 25136 12044 25188 12096
rect 25872 12087 25924 12096
rect 25872 12053 25881 12087
rect 25881 12053 25915 12087
rect 25915 12053 25924 12087
rect 25872 12044 25924 12053
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 2688 11840 2740 11892
rect 4988 11840 5040 11892
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 9036 11840 9088 11892
rect 17684 11840 17736 11892
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 5264 11772 5316 11824
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 6276 11704 6328 11756
rect 7932 11772 7984 11824
rect 9588 11704 9640 11756
rect 12808 11747 12860 11756
rect 12808 11713 12817 11747
rect 12817 11713 12851 11747
rect 12851 11713 12860 11747
rect 12808 11704 12860 11713
rect 15844 11704 15896 11756
rect 17868 11704 17920 11756
rect 19432 11840 19484 11892
rect 19616 11840 19668 11892
rect 21916 11840 21968 11892
rect 24768 11840 24820 11892
rect 21548 11772 21600 11824
rect 23020 11772 23072 11824
rect 25044 11840 25096 11892
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 19340 11704 19392 11756
rect 24308 11747 24360 11756
rect 24308 11713 24317 11747
rect 24317 11713 24351 11747
rect 24351 11713 24360 11747
rect 24308 11704 24360 11713
rect 26516 11772 26568 11824
rect 24952 11704 25004 11756
rect 25872 11704 25924 11756
rect 7656 11636 7708 11688
rect 7932 11636 7984 11688
rect 8024 11568 8076 11620
rect 9680 11636 9732 11688
rect 8392 11568 8444 11620
rect 16396 11636 16448 11688
rect 16488 11636 16540 11688
rect 24124 11636 24176 11688
rect 25964 11636 26016 11688
rect 13728 11568 13780 11620
rect 16304 11611 16356 11620
rect 16304 11577 16313 11611
rect 16313 11577 16347 11611
rect 16347 11577 16356 11611
rect 16304 11568 16356 11577
rect 19708 11611 19760 11620
rect 19708 11577 19742 11611
rect 19742 11577 19760 11611
rect 19708 11568 19760 11577
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 9496 11500 9548 11552
rect 10600 11500 10652 11552
rect 10876 11500 10928 11552
rect 12900 11500 12952 11552
rect 14096 11500 14148 11552
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 18880 11543 18932 11552
rect 18880 11509 18889 11543
rect 18889 11509 18923 11543
rect 18923 11509 18932 11543
rect 18880 11500 18932 11509
rect 20812 11543 20864 11552
rect 20812 11509 20821 11543
rect 20821 11509 20855 11543
rect 20855 11509 20864 11543
rect 20812 11500 20864 11509
rect 23848 11543 23900 11552
rect 23848 11509 23857 11543
rect 23857 11509 23891 11543
rect 23891 11509 23900 11543
rect 23848 11500 23900 11509
rect 25596 11543 25648 11552
rect 25596 11509 25605 11543
rect 25605 11509 25639 11543
rect 25639 11509 25648 11543
rect 25596 11500 25648 11509
rect 25780 11543 25832 11552
rect 25780 11509 25789 11543
rect 25789 11509 25823 11543
rect 25823 11509 25832 11543
rect 25780 11500 25832 11509
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2504 11296 2556 11348
rect 8024 11296 8076 11348
rect 9496 11339 9548 11348
rect 9496 11305 9505 11339
rect 9505 11305 9539 11339
rect 9539 11305 9548 11339
rect 9496 11296 9548 11305
rect 10876 11296 10928 11348
rect 19248 11296 19300 11348
rect 3424 11271 3476 11280
rect 3424 11237 3433 11271
rect 3433 11237 3467 11271
rect 3467 11237 3476 11271
rect 3424 11228 3476 11237
rect 7840 11228 7892 11280
rect 15844 11228 15896 11280
rect 18696 11228 18748 11280
rect 20812 11228 20864 11280
rect 5080 11203 5132 11212
rect 5080 11169 5089 11203
rect 5089 11169 5123 11203
rect 5123 11169 5132 11203
rect 5080 11160 5132 11169
rect 12900 11160 12952 11212
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 21548 11160 21600 11212
rect 22284 11296 22336 11348
rect 23296 11339 23348 11348
rect 23296 11305 23305 11339
rect 23305 11305 23339 11339
rect 23339 11305 23348 11339
rect 23296 11296 23348 11305
rect 24308 11296 24360 11348
rect 24400 11339 24452 11348
rect 24400 11305 24409 11339
rect 24409 11305 24443 11339
rect 24443 11305 24452 11339
rect 25320 11339 25372 11348
rect 24400 11296 24452 11305
rect 25320 11305 25329 11339
rect 25329 11305 25363 11339
rect 25363 11305 25372 11339
rect 25320 11296 25372 11305
rect 25780 11296 25832 11348
rect 26976 11339 27028 11348
rect 22192 11271 22244 11280
rect 22192 11237 22226 11271
rect 22226 11237 22244 11271
rect 22192 11228 22244 11237
rect 23020 11228 23072 11280
rect 24860 11228 24912 11280
rect 25044 11228 25096 11280
rect 25504 11228 25556 11280
rect 26976 11305 26985 11339
rect 26985 11305 27019 11339
rect 27019 11305 27028 11339
rect 26976 11296 27028 11305
rect 26884 11271 26936 11280
rect 26884 11237 26893 11271
rect 26893 11237 26927 11271
rect 26927 11237 26936 11271
rect 26884 11228 26936 11237
rect 25872 11203 25924 11212
rect 25872 11169 25881 11203
rect 25881 11169 25915 11203
rect 25915 11169 25924 11203
rect 25872 11160 25924 11169
rect 2596 11092 2648 11144
rect 2780 11092 2832 11144
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 2320 11024 2372 11076
rect 9956 11067 10008 11076
rect 9956 11033 9965 11067
rect 9965 11033 9999 11067
rect 9999 11033 10008 11067
rect 9956 11024 10008 11033
rect 10968 11092 11020 11144
rect 12440 11092 12492 11144
rect 5724 10999 5776 11008
rect 5724 10965 5733 10999
rect 5733 10965 5767 10999
rect 5767 10965 5776 10999
rect 5724 10956 5776 10965
rect 10324 10956 10376 11008
rect 13820 11024 13872 11076
rect 11336 10956 11388 11008
rect 24952 11092 25004 11144
rect 27160 11160 27212 11212
rect 24860 11067 24912 11076
rect 24860 11033 24869 11067
rect 24869 11033 24903 11067
rect 24903 11033 24912 11067
rect 24860 11024 24912 11033
rect 16948 10956 17000 11008
rect 17040 10956 17092 11008
rect 17868 10956 17920 11008
rect 19248 10956 19300 11008
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 1676 10752 1728 10804
rect 2504 10752 2556 10804
rect 4160 10795 4212 10804
rect 4160 10761 4169 10795
rect 4169 10761 4203 10795
rect 4203 10761 4212 10795
rect 4160 10752 4212 10761
rect 4436 10752 4488 10804
rect 2596 10684 2648 10736
rect 5080 10752 5132 10804
rect 11060 10752 11112 10804
rect 12348 10752 12400 10804
rect 12900 10795 12952 10804
rect 12900 10761 12909 10795
rect 12909 10761 12943 10795
rect 12943 10761 12952 10795
rect 12900 10752 12952 10761
rect 15844 10752 15896 10804
rect 18604 10752 18656 10804
rect 22008 10795 22060 10804
rect 22008 10761 22017 10795
rect 22017 10761 22051 10795
rect 22051 10761 22060 10795
rect 22008 10752 22060 10761
rect 22284 10795 22336 10804
rect 22284 10761 22293 10795
rect 22293 10761 22327 10795
rect 22327 10761 22336 10795
rect 22284 10752 22336 10761
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 23480 10752 23532 10761
rect 24952 10795 25004 10804
rect 24952 10761 24961 10795
rect 24961 10761 24995 10795
rect 24995 10761 25004 10795
rect 24952 10752 25004 10761
rect 25320 10795 25372 10804
rect 25320 10761 25329 10795
rect 25329 10761 25363 10795
rect 25363 10761 25372 10795
rect 25320 10752 25372 10761
rect 25872 10795 25924 10804
rect 25872 10761 25881 10795
rect 25881 10761 25915 10795
rect 25915 10761 25924 10795
rect 25872 10752 25924 10761
rect 26884 10752 26936 10804
rect 26976 10752 27028 10804
rect 5264 10616 5316 10668
rect 4620 10591 4672 10600
rect 4620 10557 4629 10591
rect 4629 10557 4663 10591
rect 4663 10557 4672 10591
rect 4620 10548 4672 10557
rect 3056 10480 3108 10532
rect 5172 10480 5224 10532
rect 2780 10455 2832 10464
rect 2780 10421 2789 10455
rect 2789 10421 2823 10455
rect 2823 10421 2832 10455
rect 14372 10684 14424 10736
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 9588 10616 9640 10668
rect 10784 10616 10836 10668
rect 10968 10616 11020 10668
rect 17500 10684 17552 10736
rect 18696 10727 18748 10736
rect 18696 10693 18705 10727
rect 18705 10693 18739 10727
rect 18739 10693 18748 10727
rect 18696 10684 18748 10693
rect 26608 10727 26660 10736
rect 16396 10616 16448 10668
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 18604 10616 18656 10668
rect 18788 10616 18840 10668
rect 23848 10616 23900 10668
rect 26608 10693 26617 10727
rect 26617 10693 26651 10727
rect 26651 10693 26660 10727
rect 26608 10684 26660 10693
rect 5540 10548 5592 10600
rect 5816 10548 5868 10600
rect 10416 10548 10468 10600
rect 16580 10548 16632 10600
rect 17132 10548 17184 10600
rect 24768 10548 24820 10600
rect 26424 10591 26476 10600
rect 26424 10557 26433 10591
rect 26433 10557 26467 10591
rect 26467 10557 26476 10591
rect 26424 10548 26476 10557
rect 5540 10455 5592 10464
rect 2780 10412 2832 10421
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 11336 10412 11388 10464
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 16396 10455 16448 10464
rect 13452 10412 13504 10421
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 16948 10412 17000 10464
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 23664 10455 23716 10464
rect 23664 10421 23673 10455
rect 23673 10421 23707 10455
rect 23707 10421 23716 10455
rect 23664 10412 23716 10421
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 2780 10208 2832 10260
rect 5172 10208 5224 10260
rect 5264 10140 5316 10192
rect 3240 10072 3292 10124
rect 5080 10072 5132 10124
rect 6644 10208 6696 10260
rect 6828 10208 6880 10260
rect 7196 10208 7248 10260
rect 10048 10208 10100 10260
rect 15384 10208 15436 10260
rect 17132 10208 17184 10260
rect 19524 10208 19576 10260
rect 21824 10208 21876 10260
rect 23848 10208 23900 10260
rect 25504 10251 25556 10260
rect 25504 10217 25513 10251
rect 25513 10217 25547 10251
rect 25547 10217 25556 10251
rect 25504 10208 25556 10217
rect 26700 10251 26752 10260
rect 26700 10217 26709 10251
rect 26709 10217 26743 10251
rect 26743 10217 26752 10251
rect 26700 10208 26752 10217
rect 10324 10183 10376 10192
rect 10324 10149 10333 10183
rect 10333 10149 10367 10183
rect 10367 10149 10376 10183
rect 10324 10140 10376 10149
rect 13912 10183 13964 10192
rect 13912 10149 13921 10183
rect 13921 10149 13955 10183
rect 13955 10149 13964 10183
rect 13912 10140 13964 10149
rect 14280 10140 14332 10192
rect 10784 10072 10836 10124
rect 12716 10072 12768 10124
rect 15660 10115 15712 10124
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 3332 10004 3384 10056
rect 3056 9936 3108 9988
rect 5632 10047 5684 10056
rect 1676 9911 1728 9920
rect 1676 9877 1685 9911
rect 1685 9877 1719 9911
rect 1719 9877 1728 9911
rect 1676 9868 1728 9877
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 10600 10047 10652 10056
rect 7104 10004 7156 10013
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 15752 10072 15804 10124
rect 17040 10140 17092 10192
rect 24952 10140 25004 10192
rect 18052 10072 18104 10124
rect 18328 10072 18380 10124
rect 21916 10115 21968 10124
rect 21916 10081 21950 10115
rect 21950 10081 21968 10115
rect 21916 10072 21968 10081
rect 25596 10072 25648 10124
rect 27344 10072 27396 10124
rect 13728 10004 13780 10056
rect 14004 10047 14056 10056
rect 14004 10013 14013 10047
rect 14013 10013 14047 10047
rect 14047 10013 14056 10047
rect 14004 10004 14056 10013
rect 14096 10047 14148 10056
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 15844 10047 15896 10056
rect 14096 10004 14148 10013
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 18696 10047 18748 10056
rect 18696 10013 18705 10047
rect 18705 10013 18739 10047
rect 18739 10013 18748 10047
rect 18696 10004 18748 10013
rect 19248 10004 19300 10056
rect 21640 10047 21692 10056
rect 21640 10013 21649 10047
rect 21649 10013 21683 10047
rect 21683 10013 21692 10047
rect 21640 10004 21692 10013
rect 24860 10047 24912 10056
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 25044 10047 25096 10056
rect 25044 10013 25053 10047
rect 25053 10013 25087 10047
rect 25087 10013 25096 10047
rect 25044 10004 25096 10013
rect 11336 9936 11388 9988
rect 14648 9979 14700 9988
rect 14648 9945 14657 9979
rect 14657 9945 14691 9979
rect 14691 9945 14700 9979
rect 14648 9936 14700 9945
rect 5816 9868 5868 9920
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 12348 9868 12400 9920
rect 12900 9868 12952 9920
rect 17960 9868 18012 9920
rect 23480 9868 23532 9920
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 2780 9707 2832 9716
rect 2780 9673 2789 9707
rect 2789 9673 2823 9707
rect 2823 9673 2832 9707
rect 2780 9664 2832 9673
rect 3240 9664 3292 9716
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 3240 9571 3292 9580
rect 2136 9528 2188 9537
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 5080 9664 5132 9716
rect 5816 9707 5868 9716
rect 5816 9673 5825 9707
rect 5825 9673 5859 9707
rect 5859 9673 5868 9707
rect 5816 9664 5868 9673
rect 10324 9664 10376 9716
rect 13176 9664 13228 9716
rect 5724 9596 5776 9648
rect 6828 9596 6880 9648
rect 5172 9528 5224 9580
rect 1676 9460 1728 9512
rect 6644 9460 6696 9512
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9588 9503 9640 9512
rect 9312 9460 9364 9469
rect 5632 9392 5684 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 5172 9324 5224 9376
rect 6368 9324 6420 9376
rect 6828 9324 6880 9376
rect 7012 9392 7064 9444
rect 9588 9469 9622 9503
rect 9622 9469 9640 9503
rect 9588 9460 9640 9469
rect 10692 9460 10744 9512
rect 11520 9460 11572 9512
rect 12900 9503 12952 9512
rect 10600 9392 10652 9444
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 14004 9664 14056 9716
rect 18604 9664 18656 9716
rect 15384 9639 15436 9648
rect 15384 9605 15393 9639
rect 15393 9605 15427 9639
rect 15427 9605 15436 9639
rect 15384 9596 15436 9605
rect 17868 9639 17920 9648
rect 17868 9605 17877 9639
rect 17877 9605 17911 9639
rect 17911 9605 17920 9639
rect 17868 9596 17920 9605
rect 18328 9639 18380 9648
rect 18328 9605 18337 9639
rect 18337 9605 18371 9639
rect 18371 9605 18380 9639
rect 18328 9596 18380 9605
rect 18788 9596 18840 9648
rect 14096 9528 14148 9580
rect 14740 9528 14792 9580
rect 15844 9528 15896 9580
rect 19708 9596 19760 9648
rect 20536 9596 20588 9648
rect 21640 9664 21692 9716
rect 21916 9664 21968 9716
rect 21364 9528 21416 9580
rect 21456 9528 21508 9580
rect 23204 9664 23256 9716
rect 25412 9664 25464 9716
rect 27344 9707 27396 9716
rect 27344 9673 27353 9707
rect 27353 9673 27387 9707
rect 27387 9673 27396 9707
rect 27344 9664 27396 9673
rect 24860 9596 24912 9648
rect 26608 9639 26660 9648
rect 26608 9605 26617 9639
rect 26617 9605 26651 9639
rect 26651 9605 26660 9639
rect 26608 9596 26660 9605
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 12256 9324 12308 9376
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 12992 9324 13044 9376
rect 14648 9460 14700 9512
rect 18880 9460 18932 9512
rect 19524 9460 19576 9512
rect 24952 9528 25004 9580
rect 25412 9528 25464 9580
rect 23756 9460 23808 9512
rect 26332 9460 26384 9512
rect 19156 9392 19208 9444
rect 21916 9392 21968 9444
rect 22100 9392 22152 9444
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 14188 9324 14240 9376
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 18788 9367 18840 9376
rect 18788 9333 18797 9367
rect 18797 9333 18831 9367
rect 18831 9333 18840 9367
rect 18788 9324 18840 9333
rect 19064 9367 19116 9376
rect 19064 9333 19073 9367
rect 19073 9333 19107 9367
rect 19107 9333 19116 9367
rect 19064 9324 19116 9333
rect 19524 9367 19576 9376
rect 19524 9333 19533 9367
rect 19533 9333 19567 9367
rect 19567 9333 19576 9367
rect 19524 9324 19576 9333
rect 23572 9392 23624 9444
rect 25504 9392 25556 9444
rect 25044 9367 25096 9376
rect 25044 9333 25053 9367
rect 25053 9333 25087 9367
rect 25087 9333 25096 9367
rect 25044 9324 25096 9333
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 2688 9163 2740 9172
rect 2688 9129 2697 9163
rect 2697 9129 2731 9163
rect 2731 9129 2740 9163
rect 2688 9120 2740 9129
rect 9220 9120 9272 9172
rect 10048 9120 10100 9172
rect 11336 9120 11388 9172
rect 11704 9163 11756 9172
rect 11704 9129 11713 9163
rect 11713 9129 11747 9163
rect 11747 9129 11756 9163
rect 11704 9120 11756 9129
rect 12900 9120 12952 9172
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 14004 9120 14056 9172
rect 14740 9163 14792 9172
rect 14740 9129 14749 9163
rect 14749 9129 14783 9163
rect 14783 9129 14792 9163
rect 14740 9120 14792 9129
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 15752 9120 15804 9129
rect 16396 9120 16448 9172
rect 18696 9120 18748 9172
rect 18880 9163 18932 9172
rect 18880 9129 18889 9163
rect 18889 9129 18923 9163
rect 18923 9129 18932 9163
rect 18880 9120 18932 9129
rect 24860 9163 24912 9172
rect 24860 9129 24869 9163
rect 24869 9129 24903 9163
rect 24903 9129 24912 9163
rect 24860 9120 24912 9129
rect 25228 9163 25280 9172
rect 25228 9129 25237 9163
rect 25237 9129 25271 9163
rect 25271 9129 25280 9163
rect 25228 9120 25280 9129
rect 25320 9163 25372 9172
rect 25320 9129 25329 9163
rect 25329 9129 25363 9163
rect 25363 9129 25372 9163
rect 26700 9163 26752 9172
rect 25320 9120 25372 9129
rect 26700 9129 26709 9163
rect 26709 9129 26743 9163
rect 26743 9129 26752 9163
rect 26700 9120 26752 9129
rect 10692 9052 10744 9104
rect 12716 9095 12768 9104
rect 1676 8984 1728 9036
rect 2136 8984 2188 9036
rect 2504 9027 2556 9036
rect 2504 8993 2513 9027
rect 2513 8993 2547 9027
rect 2547 8993 2556 9027
rect 2504 8984 2556 8993
rect 10600 8984 10652 9036
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 6644 8916 6696 8968
rect 11428 8916 11480 8968
rect 12256 8984 12308 9036
rect 12716 9061 12725 9095
rect 12725 9061 12759 9095
rect 12759 9061 12768 9095
rect 12716 9052 12768 9061
rect 12992 8984 13044 9036
rect 13176 8984 13228 9036
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 19064 9052 19116 9104
rect 25044 9052 25096 9104
rect 11888 8916 11940 8925
rect 16396 8959 16448 8968
rect 16396 8925 16405 8959
rect 16405 8925 16439 8959
rect 16439 8925 16448 8959
rect 16396 8916 16448 8925
rect 16488 8959 16540 8968
rect 16488 8925 16497 8959
rect 16497 8925 16531 8959
rect 16531 8925 16540 8959
rect 16488 8916 16540 8925
rect 17868 8916 17920 8968
rect 18144 8984 18196 9036
rect 19800 8984 19852 9036
rect 23388 8984 23440 9036
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 12808 8848 12860 8900
rect 18880 8916 18932 8968
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 22008 8959 22060 8968
rect 22008 8925 22017 8959
rect 22017 8925 22051 8959
rect 22051 8925 22060 8959
rect 22008 8916 22060 8925
rect 23848 8959 23900 8968
rect 18328 8848 18380 8900
rect 21824 8848 21876 8900
rect 23848 8925 23857 8959
rect 23857 8925 23891 8959
rect 23891 8925 23900 8959
rect 23848 8916 23900 8925
rect 25504 8959 25556 8968
rect 25504 8925 25513 8959
rect 25513 8925 25547 8959
rect 25547 8925 25556 8959
rect 25504 8916 25556 8925
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2872 8780 2924 8832
rect 3700 8823 3752 8832
rect 3700 8789 3709 8823
rect 3709 8789 3743 8823
rect 3743 8789 3752 8823
rect 3700 8780 3752 8789
rect 7012 8823 7064 8832
rect 7012 8789 7021 8823
rect 7021 8789 7055 8823
rect 7055 8789 7064 8823
rect 7012 8780 7064 8789
rect 12348 8780 12400 8832
rect 14188 8780 14240 8832
rect 14280 8780 14332 8832
rect 14648 8780 14700 8832
rect 15844 8780 15896 8832
rect 17500 8823 17552 8832
rect 17500 8789 17509 8823
rect 17509 8789 17543 8823
rect 17543 8789 17552 8823
rect 17500 8780 17552 8789
rect 21548 8823 21600 8832
rect 21548 8789 21557 8823
rect 21557 8789 21591 8823
rect 21591 8789 21600 8823
rect 21548 8780 21600 8789
rect 23756 8823 23808 8832
rect 23756 8789 23765 8823
rect 23765 8789 23799 8823
rect 23799 8789 23808 8823
rect 23756 8780 23808 8789
rect 24676 8780 24728 8832
rect 25872 8823 25924 8832
rect 25872 8789 25881 8823
rect 25881 8789 25915 8823
rect 25915 8789 25924 8823
rect 25872 8780 25924 8789
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 7012 8576 7064 8628
rect 13360 8576 13412 8628
rect 14096 8576 14148 8628
rect 16304 8576 16356 8628
rect 17868 8576 17920 8628
rect 18052 8576 18104 8628
rect 18696 8576 18748 8628
rect 1584 8551 1636 8560
rect 1584 8517 1593 8551
rect 1593 8517 1627 8551
rect 1627 8517 1636 8551
rect 1584 8508 1636 8517
rect 9312 8508 9364 8560
rect 3700 8440 3752 8492
rect 2044 8372 2096 8424
rect 4068 8372 4120 8424
rect 2504 8304 2556 8356
rect 3884 8304 3936 8356
rect 3608 8279 3660 8288
rect 3608 8245 3617 8279
rect 3617 8245 3651 8279
rect 3651 8245 3660 8279
rect 3608 8236 3660 8245
rect 6276 8440 6328 8492
rect 6552 8440 6604 8492
rect 6644 8372 6696 8424
rect 10048 8415 10100 8424
rect 10048 8381 10057 8415
rect 10057 8381 10091 8415
rect 10091 8381 10100 8415
rect 10048 8372 10100 8381
rect 13176 8508 13228 8560
rect 10232 8372 10284 8424
rect 6552 8347 6604 8356
rect 6552 8313 6561 8347
rect 6561 8313 6595 8347
rect 6595 8313 6604 8347
rect 6552 8304 6604 8313
rect 10600 8304 10652 8356
rect 15292 8304 15344 8356
rect 15476 8347 15528 8356
rect 15476 8313 15485 8347
rect 15485 8313 15519 8347
rect 15519 8313 15528 8347
rect 16488 8372 16540 8424
rect 19432 8483 19484 8492
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 19708 8576 19760 8628
rect 20536 8619 20588 8628
rect 20536 8585 20545 8619
rect 20545 8585 20579 8619
rect 20579 8585 20588 8619
rect 20536 8576 20588 8585
rect 21824 8576 21876 8628
rect 22008 8576 22060 8628
rect 23388 8619 23440 8628
rect 23388 8585 23397 8619
rect 23397 8585 23431 8619
rect 23431 8585 23440 8619
rect 23388 8576 23440 8585
rect 24492 8619 24544 8628
rect 24492 8585 24501 8619
rect 24501 8585 24535 8619
rect 24535 8585 24544 8619
rect 24492 8576 24544 8585
rect 25228 8576 25280 8628
rect 25412 8619 25464 8628
rect 25412 8585 25421 8619
rect 25421 8585 25455 8619
rect 25455 8585 25464 8619
rect 25412 8576 25464 8585
rect 26516 8619 26568 8628
rect 26516 8585 26525 8619
rect 26525 8585 26559 8619
rect 26559 8585 26568 8619
rect 26516 8576 26568 8585
rect 27160 8619 27212 8628
rect 27160 8585 27169 8619
rect 27169 8585 27203 8619
rect 27203 8585 27212 8619
rect 27160 8576 27212 8585
rect 21916 8440 21968 8492
rect 22100 8440 22152 8492
rect 25320 8483 25372 8492
rect 25320 8449 25329 8483
rect 25329 8449 25363 8483
rect 25363 8449 25372 8483
rect 25320 8440 25372 8449
rect 25964 8440 26016 8492
rect 26148 8440 26200 8492
rect 18788 8372 18840 8424
rect 18880 8415 18932 8424
rect 18880 8381 18889 8415
rect 18889 8381 18923 8415
rect 18923 8381 18932 8415
rect 18880 8372 18932 8381
rect 19616 8372 19668 8424
rect 15476 8304 15528 8313
rect 15936 8347 15988 8356
rect 15936 8313 15970 8347
rect 15970 8313 15988 8347
rect 15936 8304 15988 8313
rect 17224 8304 17276 8356
rect 21824 8372 21876 8424
rect 23848 8372 23900 8424
rect 25872 8372 25924 8424
rect 24492 8304 24544 8356
rect 4712 8236 4764 8288
rect 6644 8236 6696 8288
rect 11888 8279 11940 8288
rect 11888 8245 11897 8279
rect 11897 8245 11931 8279
rect 11931 8245 11940 8279
rect 11888 8236 11940 8245
rect 22376 8236 22428 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 3608 8032 3660 8084
rect 4068 8032 4120 8084
rect 4344 8032 4396 8084
rect 11428 8075 11480 8084
rect 11428 8041 11437 8075
rect 11437 8041 11471 8075
rect 11471 8041 11480 8075
rect 11428 8032 11480 8041
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 12716 8032 12768 8084
rect 16396 8032 16448 8084
rect 17500 8032 17552 8084
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 19248 8032 19300 8084
rect 19616 8032 19668 8084
rect 19708 8075 19760 8084
rect 19708 8041 19717 8075
rect 19717 8041 19751 8075
rect 19751 8041 19760 8075
rect 19708 8032 19760 8041
rect 22008 8032 22060 8084
rect 22376 8075 22428 8084
rect 22376 8041 22385 8075
rect 22385 8041 22419 8075
rect 22419 8041 22428 8075
rect 22376 8032 22428 8041
rect 23940 8032 23992 8084
rect 25136 8032 25188 8084
rect 25872 8075 25924 8084
rect 25872 8041 25881 8075
rect 25881 8041 25915 8075
rect 25915 8041 25924 8075
rect 25872 8032 25924 8041
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 4620 7964 4672 8016
rect 10324 8007 10376 8016
rect 10324 7973 10333 8007
rect 10333 7973 10367 8007
rect 10367 7973 10376 8007
rect 10324 7964 10376 7973
rect 17868 7964 17920 8016
rect 21916 8007 21968 8016
rect 21916 7973 21925 8007
rect 21925 7973 21959 8007
rect 21959 7973 21968 8007
rect 21916 7964 21968 7973
rect 6276 7896 6328 7948
rect 9036 7896 9088 7948
rect 10048 7896 10100 7948
rect 17132 7939 17184 7948
rect 17132 7905 17141 7939
rect 17141 7905 17175 7939
rect 17175 7905 17184 7939
rect 17132 7896 17184 7905
rect 21364 7896 21416 7948
rect 23112 7896 23164 7948
rect 26332 7964 26384 8016
rect 25044 7896 25096 7948
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 2688 7760 2740 7812
rect 3884 7828 3936 7880
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 10508 7828 10560 7880
rect 17040 7828 17092 7880
rect 17224 7828 17276 7880
rect 22836 7871 22888 7880
rect 22836 7837 22845 7871
rect 22845 7837 22879 7871
rect 22879 7837 22888 7871
rect 22836 7828 22888 7837
rect 22928 7828 22980 7880
rect 23388 7828 23440 7880
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 6644 7692 6696 7744
rect 16396 7692 16448 7744
rect 16488 7692 16540 7744
rect 17408 7692 17460 7744
rect 24124 7735 24176 7744
rect 24124 7701 24133 7735
rect 24133 7701 24167 7735
rect 24167 7701 24176 7735
rect 24124 7692 24176 7701
rect 25504 7735 25556 7744
rect 25504 7701 25513 7735
rect 25513 7701 25547 7735
rect 25547 7701 25556 7735
rect 25504 7692 25556 7701
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 4344 7488 4396 7540
rect 6276 7531 6328 7540
rect 6276 7497 6285 7531
rect 6285 7497 6319 7531
rect 6319 7497 6328 7531
rect 6276 7488 6328 7497
rect 6552 7488 6604 7540
rect 17500 7488 17552 7540
rect 18420 7488 18472 7540
rect 17224 7463 17276 7472
rect 17224 7429 17233 7463
rect 17233 7429 17267 7463
rect 17267 7429 17276 7463
rect 17224 7420 17276 7429
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 6644 7352 6696 7404
rect 12256 7352 12308 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 15200 7352 15252 7404
rect 21824 7488 21876 7540
rect 25044 7531 25096 7540
rect 25044 7497 25053 7531
rect 25053 7497 25087 7531
rect 25087 7497 25096 7531
rect 25044 7488 25096 7497
rect 26516 7488 26568 7540
rect 27620 7531 27672 7540
rect 27620 7497 27629 7531
rect 27629 7497 27663 7531
rect 27663 7497 27672 7531
rect 27620 7488 27672 7497
rect 22836 7420 22888 7472
rect 26332 7420 26384 7472
rect 19432 7352 19484 7404
rect 22284 7352 22336 7404
rect 22928 7352 22980 7404
rect 24124 7352 24176 7404
rect 1952 7284 2004 7336
rect 9128 7284 9180 7336
rect 10324 7284 10376 7336
rect 16304 7284 16356 7336
rect 23940 7284 23992 7336
rect 2044 7259 2096 7268
rect 2044 7225 2053 7259
rect 2053 7225 2087 7259
rect 2087 7225 2096 7259
rect 2044 7216 2096 7225
rect 7012 7216 7064 7268
rect 9588 7216 9640 7268
rect 11888 7216 11940 7268
rect 16396 7216 16448 7268
rect 17776 7216 17828 7268
rect 23388 7216 23440 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 3884 7148 3936 7157
rect 3976 7148 4028 7200
rect 4712 7148 4764 7200
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 13912 7148 13964 7200
rect 15200 7191 15252 7200
rect 15200 7157 15209 7191
rect 15209 7157 15243 7191
rect 15243 7157 15252 7191
rect 15200 7148 15252 7157
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 18696 7191 18748 7200
rect 18696 7157 18705 7191
rect 18705 7157 18739 7191
rect 18739 7157 18748 7191
rect 18696 7148 18748 7157
rect 22468 7191 22520 7200
rect 22468 7157 22477 7191
rect 22477 7157 22511 7191
rect 22511 7157 22520 7191
rect 22468 7148 22520 7157
rect 23112 7191 23164 7200
rect 23112 7157 23121 7191
rect 23121 7157 23155 7191
rect 23155 7157 23164 7191
rect 23112 7148 23164 7157
rect 27436 7327 27488 7336
rect 27436 7293 27445 7327
rect 27445 7293 27479 7327
rect 27479 7293 27488 7327
rect 27436 7284 27488 7293
rect 24308 7148 24360 7200
rect 24676 7191 24728 7200
rect 24676 7157 24685 7191
rect 24685 7157 24719 7191
rect 24719 7157 24728 7191
rect 24676 7148 24728 7157
rect 25228 7148 25280 7200
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 9128 6987 9180 6996
rect 9128 6953 9137 6987
rect 9137 6953 9171 6987
rect 9171 6953 9180 6987
rect 9128 6944 9180 6953
rect 9680 6944 9732 6996
rect 17132 6944 17184 6996
rect 17776 6987 17828 6996
rect 17776 6953 17785 6987
rect 17785 6953 17819 6987
rect 17819 6953 17828 6987
rect 17776 6944 17828 6953
rect 19156 6987 19208 6996
rect 19156 6953 19165 6987
rect 19165 6953 19199 6987
rect 19199 6953 19208 6987
rect 19156 6944 19208 6953
rect 19616 6944 19668 6996
rect 20536 6944 20588 6996
rect 22468 6944 22520 6996
rect 23296 6944 23348 6996
rect 17868 6876 17920 6928
rect 22284 6876 22336 6928
rect 22836 6919 22888 6928
rect 22836 6885 22845 6919
rect 22845 6885 22879 6919
rect 22879 6885 22888 6919
rect 22836 6876 22888 6885
rect 2136 6808 2188 6860
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 2688 6808 2740 6860
rect 6828 6851 6880 6860
rect 6828 6817 6837 6851
rect 6837 6817 6871 6851
rect 6871 6817 6880 6851
rect 6828 6808 6880 6817
rect 11612 6851 11664 6860
rect 11612 6817 11621 6851
rect 11621 6817 11655 6851
rect 11655 6817 11664 6851
rect 11612 6808 11664 6817
rect 11796 6808 11848 6860
rect 12624 6808 12676 6860
rect 13452 6808 13504 6860
rect 19248 6851 19300 6860
rect 19248 6817 19257 6851
rect 19257 6817 19291 6851
rect 19291 6817 19300 6851
rect 19248 6808 19300 6817
rect 23204 6808 23256 6860
rect 24216 6808 24268 6860
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 27344 6808 27396 6860
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 10140 6783 10192 6792
rect 2596 6672 2648 6724
rect 6552 6672 6604 6724
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10416 6740 10468 6792
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 13820 6783 13872 6792
rect 13820 6749 13829 6783
rect 13829 6749 13863 6783
rect 13863 6749 13872 6783
rect 13820 6740 13872 6749
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 15016 6740 15068 6792
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 23572 6783 23624 6792
rect 23572 6749 23581 6783
rect 23581 6749 23615 6783
rect 23615 6749 23624 6783
rect 23572 6740 23624 6749
rect 9772 6672 9824 6724
rect 13360 6715 13412 6724
rect 13360 6681 13369 6715
rect 13369 6681 13403 6715
rect 13403 6681 13412 6715
rect 13360 6672 13412 6681
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 3884 6604 3936 6656
rect 6736 6604 6788 6656
rect 7380 6604 7432 6656
rect 13084 6604 13136 6656
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 16488 6604 16540 6656
rect 16672 6647 16724 6656
rect 16672 6613 16681 6647
rect 16681 6613 16715 6647
rect 16715 6613 16724 6647
rect 16672 6604 16724 6613
rect 18512 6604 18564 6656
rect 25228 6647 25280 6656
rect 25228 6613 25237 6647
rect 25237 6613 25271 6647
rect 25271 6613 25280 6647
rect 25228 6604 25280 6613
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 2136 6400 2188 6452
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 2872 6400 2924 6452
rect 6828 6400 6880 6452
rect 6920 6400 6972 6452
rect 10140 6400 10192 6452
rect 11796 6400 11848 6452
rect 11888 6400 11940 6452
rect 13912 6400 13964 6452
rect 15752 6400 15804 6452
rect 16488 6400 16540 6452
rect 19156 6443 19208 6452
rect 19156 6409 19165 6443
rect 19165 6409 19199 6443
rect 19199 6409 19208 6443
rect 19156 6400 19208 6409
rect 19248 6400 19300 6452
rect 23296 6400 23348 6452
rect 23480 6400 23532 6452
rect 27344 6443 27396 6452
rect 27344 6409 27353 6443
rect 27353 6409 27387 6443
rect 27387 6409 27396 6443
rect 27344 6400 27396 6409
rect 6552 6375 6604 6384
rect 6552 6341 6561 6375
rect 6561 6341 6595 6375
rect 6595 6341 6604 6375
rect 6552 6332 6604 6341
rect 7012 6264 7064 6316
rect 3240 6196 3292 6248
rect 1952 6128 2004 6180
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 10416 6332 10468 6384
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 11336 6264 11388 6316
rect 23572 6332 23624 6384
rect 24124 6332 24176 6384
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13403 6307
rect 13403 6273 13412 6307
rect 13360 6264 13412 6273
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 13084 6196 13136 6248
rect 13820 6264 13872 6316
rect 15200 6264 15252 6316
rect 16672 6264 16724 6316
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 19616 6307 19668 6316
rect 18604 6264 18656 6273
rect 19616 6273 19625 6307
rect 19625 6273 19659 6307
rect 19659 6273 19668 6307
rect 19616 6264 19668 6273
rect 23204 6264 23256 6316
rect 25228 6332 25280 6384
rect 26608 6375 26660 6384
rect 26608 6341 26617 6375
rect 26617 6341 26651 6375
rect 26651 6341 26660 6375
rect 26608 6332 26660 6341
rect 15568 6239 15620 6248
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 18696 6196 18748 6248
rect 19432 6196 19484 6248
rect 23480 6239 23532 6248
rect 23480 6205 23489 6239
rect 23489 6205 23523 6239
rect 23523 6205 23532 6239
rect 23480 6196 23532 6205
rect 24768 6196 24820 6248
rect 26424 6239 26476 6248
rect 26424 6205 26433 6239
rect 26433 6205 26467 6239
rect 26467 6205 26476 6239
rect 26424 6196 26476 6205
rect 3884 6171 3936 6180
rect 3884 6137 3893 6171
rect 3893 6137 3927 6171
rect 3927 6137 3936 6171
rect 3884 6128 3936 6137
rect 4988 6128 5040 6180
rect 7564 6128 7616 6180
rect 10048 6128 10100 6180
rect 10508 6171 10560 6180
rect 10508 6137 10517 6171
rect 10517 6137 10551 6171
rect 10551 6137 10560 6171
rect 10508 6128 10560 6137
rect 12808 6171 12860 6180
rect 12808 6137 12817 6171
rect 12817 6137 12851 6171
rect 12851 6137 12860 6171
rect 12808 6128 12860 6137
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 2504 6060 2556 6112
rect 5356 6103 5408 6112
rect 5356 6069 5365 6103
rect 5365 6069 5399 6103
rect 5399 6069 5408 6103
rect 5356 6060 5408 6069
rect 11612 6103 11664 6112
rect 11612 6069 11621 6103
rect 11621 6069 11655 6103
rect 11655 6069 11664 6103
rect 11612 6060 11664 6069
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 15844 6128 15896 6180
rect 24216 6128 24268 6180
rect 13360 6060 13412 6112
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 17960 6060 18012 6112
rect 20812 6060 20864 6112
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 1400 5856 1452 5908
rect 2412 5856 2464 5908
rect 2688 5788 2740 5840
rect 6920 5856 6972 5908
rect 7012 5899 7064 5908
rect 7012 5865 7021 5899
rect 7021 5865 7055 5899
rect 7055 5865 7064 5899
rect 7012 5856 7064 5865
rect 7380 5856 7432 5908
rect 8024 5856 8076 5908
rect 9588 5856 9640 5908
rect 11612 5856 11664 5908
rect 12256 5899 12308 5908
rect 12256 5865 12265 5899
rect 12265 5865 12299 5899
rect 12299 5865 12308 5899
rect 12256 5856 12308 5865
rect 13176 5856 13228 5908
rect 15660 5856 15712 5908
rect 18512 5856 18564 5908
rect 19432 5899 19484 5908
rect 19432 5865 19441 5899
rect 19441 5865 19475 5899
rect 19475 5865 19484 5899
rect 19432 5856 19484 5865
rect 24124 5899 24176 5908
rect 24124 5865 24133 5899
rect 24133 5865 24167 5899
rect 24167 5865 24176 5899
rect 24124 5856 24176 5865
rect 17960 5788 18012 5840
rect 22744 5788 22796 5840
rect 4160 5720 4212 5772
rect 5448 5720 5500 5772
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 15200 5720 15252 5772
rect 15752 5720 15804 5772
rect 21364 5720 21416 5772
rect 2412 5652 2464 5704
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4528 5652 4580 5661
rect 4988 5652 5040 5704
rect 7012 5652 7064 5704
rect 7932 5652 7984 5704
rect 5356 5584 5408 5636
rect 9496 5652 9548 5704
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 13084 5695 13136 5704
rect 13084 5661 13093 5695
rect 13093 5661 13127 5695
rect 13127 5661 13136 5695
rect 13084 5652 13136 5661
rect 15384 5652 15436 5704
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 19064 5695 19116 5704
rect 19064 5661 19073 5695
rect 19073 5661 19107 5695
rect 19107 5661 19116 5695
rect 19064 5652 19116 5661
rect 23388 5720 23440 5772
rect 24676 5720 24728 5772
rect 27068 5720 27120 5772
rect 26700 5627 26752 5636
rect 26700 5593 26709 5627
rect 26709 5593 26743 5627
rect 26743 5593 26752 5627
rect 26700 5584 26752 5593
rect 2596 5516 2648 5568
rect 12992 5516 13044 5568
rect 13452 5559 13504 5568
rect 13452 5525 13461 5559
rect 13461 5525 13495 5559
rect 13495 5525 13504 5559
rect 13452 5516 13504 5525
rect 14556 5516 14608 5568
rect 15016 5559 15068 5568
rect 15016 5525 15025 5559
rect 15025 5525 15059 5559
rect 15059 5525 15068 5559
rect 15016 5516 15068 5525
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 19156 5516 19208 5568
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 2412 5355 2464 5364
rect 2412 5321 2421 5355
rect 2421 5321 2455 5355
rect 2455 5321 2464 5355
rect 2412 5312 2464 5321
rect 4068 5312 4120 5364
rect 4988 5355 5040 5364
rect 4988 5321 4997 5355
rect 4997 5321 5031 5355
rect 5031 5321 5040 5355
rect 4988 5312 5040 5321
rect 5448 5312 5500 5364
rect 7564 5355 7616 5364
rect 7564 5321 7573 5355
rect 7573 5321 7607 5355
rect 7607 5321 7616 5355
rect 7564 5312 7616 5321
rect 8024 5312 8076 5364
rect 8576 5355 8628 5364
rect 8576 5321 8585 5355
rect 8585 5321 8619 5355
rect 8619 5321 8628 5355
rect 8576 5312 8628 5321
rect 3056 5176 3108 5228
rect 3976 5176 4028 5228
rect 4620 5219 4672 5228
rect 4620 5185 4629 5219
rect 4629 5185 4663 5219
rect 4663 5185 4672 5219
rect 4620 5176 4672 5185
rect 9496 5312 9548 5364
rect 12164 5355 12216 5364
rect 12164 5321 12173 5355
rect 12173 5321 12207 5355
rect 12207 5321 12216 5355
rect 12164 5312 12216 5321
rect 15200 5312 15252 5364
rect 15384 5355 15436 5364
rect 15384 5321 15393 5355
rect 15393 5321 15427 5355
rect 15427 5321 15436 5355
rect 15384 5312 15436 5321
rect 15660 5355 15712 5364
rect 15660 5321 15669 5355
rect 15669 5321 15703 5355
rect 15703 5321 15712 5355
rect 15660 5312 15712 5321
rect 17868 5355 17920 5364
rect 17868 5321 17877 5355
rect 17877 5321 17911 5355
rect 17911 5321 17920 5355
rect 17868 5312 17920 5321
rect 18880 5355 18932 5364
rect 18880 5321 18889 5355
rect 18889 5321 18923 5355
rect 18923 5321 18932 5355
rect 18880 5312 18932 5321
rect 22744 5355 22796 5364
rect 22744 5321 22753 5355
rect 22753 5321 22787 5355
rect 22787 5321 22796 5355
rect 22744 5312 22796 5321
rect 23388 5355 23440 5364
rect 23388 5321 23397 5355
rect 23397 5321 23431 5355
rect 23431 5321 23440 5355
rect 23388 5312 23440 5321
rect 27068 5312 27120 5364
rect 14372 5244 14424 5296
rect 19064 5244 19116 5296
rect 12256 5176 12308 5228
rect 15844 5176 15896 5228
rect 18604 5176 18656 5228
rect 20812 5176 20864 5228
rect 5080 5108 5132 5160
rect 19064 5108 19116 5160
rect 2044 5083 2096 5092
rect 2044 5049 2053 5083
rect 2053 5049 2087 5083
rect 2087 5049 2096 5083
rect 2044 5040 2096 5049
rect 4436 5083 4488 5092
rect 4436 5049 4445 5083
rect 4445 5049 4479 5083
rect 4479 5049 4488 5083
rect 4436 5040 4488 5049
rect 4528 5040 4580 5092
rect 8024 5083 8076 5092
rect 8024 5049 8033 5083
rect 8033 5049 8067 5083
rect 8067 5049 8076 5083
rect 8024 5040 8076 5049
rect 13084 5040 13136 5092
rect 15108 5040 15160 5092
rect 19248 5083 19300 5092
rect 19248 5049 19257 5083
rect 19257 5049 19291 5083
rect 19291 5049 19300 5083
rect 19248 5040 19300 5049
rect 21364 5151 21416 5160
rect 21364 5117 21373 5151
rect 21373 5117 21407 5151
rect 21407 5117 21416 5151
rect 21364 5108 21416 5117
rect 26424 5151 26476 5160
rect 26424 5117 26433 5151
rect 26433 5117 26467 5151
rect 26467 5117 26476 5151
rect 26424 5108 26476 5117
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 8208 4972 8260 5024
rect 26608 5015 26660 5024
rect 26608 4981 26617 5015
rect 26617 4981 26651 5015
rect 26651 4981 26660 5015
rect 26608 4972 26660 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 2688 4768 2740 4820
rect 4528 4768 4580 4820
rect 11336 4768 11388 4820
rect 12532 4811 12584 4820
rect 12532 4777 12541 4811
rect 12541 4777 12575 4811
rect 12575 4777 12584 4811
rect 12532 4768 12584 4777
rect 2872 4700 2924 4752
rect 3240 4632 3292 4684
rect 3884 4632 3936 4684
rect 7104 4675 7156 4684
rect 7104 4641 7138 4675
rect 7138 4641 7156 4675
rect 7104 4632 7156 4641
rect 10140 4700 10192 4752
rect 9772 4632 9824 4684
rect 12900 4768 12952 4820
rect 15292 4768 15344 4820
rect 15844 4768 15896 4820
rect 18880 4768 18932 4820
rect 19248 4811 19300 4820
rect 19248 4777 19257 4811
rect 19257 4777 19291 4811
rect 19291 4777 19300 4811
rect 19248 4768 19300 4777
rect 19892 4768 19944 4820
rect 21364 4811 21416 4820
rect 21364 4777 21373 4811
rect 21373 4777 21407 4811
rect 21407 4777 21416 4811
rect 21364 4768 21416 4777
rect 12992 4743 13044 4752
rect 12992 4709 13001 4743
rect 13001 4709 13035 4743
rect 13035 4709 13044 4743
rect 12992 4700 13044 4709
rect 19432 4700 19484 4752
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 26516 4675 26568 4684
rect 4068 4564 4120 4616
rect 4620 4564 4672 4616
rect 5448 4564 5500 4616
rect 6552 4564 6604 4616
rect 12716 4564 12768 4616
rect 14372 4564 14424 4616
rect 16304 4564 16356 4616
rect 19248 4564 19300 4616
rect 26516 4641 26525 4675
rect 26525 4641 26559 4675
rect 26559 4641 26568 4675
rect 26516 4632 26568 4641
rect 27344 4632 27396 4684
rect 1492 4496 1544 4548
rect 1952 4496 2004 4548
rect 1400 4428 1452 4480
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 3884 4471 3936 4480
rect 3884 4437 3893 4471
rect 3893 4437 3927 4471
rect 3927 4437 3936 4471
rect 3884 4428 3936 4437
rect 8208 4471 8260 4480
rect 8208 4437 8217 4471
rect 8217 4437 8251 4471
rect 8251 4437 8260 4471
rect 8208 4428 8260 4437
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 3056 4224 3108 4276
rect 4252 4224 4304 4276
rect 4436 4224 4488 4276
rect 7104 4267 7156 4276
rect 7104 4233 7113 4267
rect 7113 4233 7147 4267
rect 7147 4233 7156 4267
rect 7104 4224 7156 4233
rect 8024 4267 8076 4276
rect 8024 4233 8033 4267
rect 8033 4233 8067 4267
rect 8067 4233 8076 4267
rect 8024 4224 8076 4233
rect 9772 4267 9824 4276
rect 9772 4233 9781 4267
rect 9781 4233 9815 4267
rect 9815 4233 9824 4267
rect 9772 4224 9824 4233
rect 10140 4267 10192 4276
rect 10140 4233 10149 4267
rect 10149 4233 10183 4267
rect 10183 4233 10192 4267
rect 10140 4224 10192 4233
rect 12716 4267 12768 4276
rect 12716 4233 12725 4267
rect 12725 4233 12759 4267
rect 12759 4233 12768 4267
rect 12716 4224 12768 4233
rect 12900 4224 12952 4276
rect 14372 4267 14424 4276
rect 14372 4233 14381 4267
rect 14381 4233 14415 4267
rect 14415 4233 14424 4267
rect 14372 4224 14424 4233
rect 15752 4224 15804 4276
rect 19064 4267 19116 4276
rect 19064 4233 19073 4267
rect 19073 4233 19107 4267
rect 19107 4233 19116 4267
rect 19064 4224 19116 4233
rect 19892 4224 19944 4276
rect 27344 4267 27396 4276
rect 27344 4233 27353 4267
rect 27353 4233 27387 4267
rect 27387 4233 27396 4267
rect 27344 4224 27396 4233
rect 8208 4156 8260 4208
rect 4620 4088 4672 4140
rect 5448 4088 5500 4140
rect 12992 4088 13044 4140
rect 16304 4156 16356 4208
rect 1492 4063 1544 4072
rect 1492 4029 1501 4063
rect 1501 4029 1535 4063
rect 1535 4029 1544 4063
rect 1492 4020 1544 4029
rect 3240 4063 3292 4072
rect 3240 4029 3249 4063
rect 3249 4029 3283 4063
rect 3283 4029 3292 4063
rect 3240 4020 3292 4029
rect 4252 4020 4304 4072
rect 9588 4020 9640 4072
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 19248 4088 19300 4140
rect 19432 4088 19484 4140
rect 26424 4063 26476 4072
rect 26424 4029 26433 4063
rect 26433 4029 26467 4063
rect 26467 4029 26476 4063
rect 26424 4020 26476 4029
rect 27528 4063 27580 4072
rect 27528 4029 27537 4063
rect 27537 4029 27571 4063
rect 27571 4029 27580 4063
rect 27528 4020 27580 4029
rect 2320 3952 2372 4004
rect 2780 3952 2832 4004
rect 8392 3995 8444 4004
rect 8392 3961 8401 3995
rect 8401 3961 8435 3995
rect 8435 3961 8444 3995
rect 8392 3952 8444 3961
rect 18972 3952 19024 4004
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 5080 3884 5132 3893
rect 6552 3927 6604 3936
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 18880 3927 18932 3936
rect 18880 3893 18889 3927
rect 18889 3893 18923 3927
rect 18923 3893 18932 3927
rect 18880 3884 18932 3893
rect 19616 3884 19668 3936
rect 26608 3927 26660 3936
rect 26608 3893 26617 3927
rect 26617 3893 26651 3927
rect 26651 3893 26660 3927
rect 26608 3884 26660 3893
rect 27712 3927 27764 3936
rect 27712 3893 27721 3927
rect 27721 3893 27755 3927
rect 27755 3893 27764 3927
rect 27712 3884 27764 3893
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2320 3680 2372 3689
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 4068 3723 4120 3732
rect 4068 3689 4077 3723
rect 4077 3689 4111 3723
rect 4111 3689 4120 3723
rect 4068 3680 4120 3689
rect 8392 3680 8444 3732
rect 15844 3723 15896 3732
rect 15844 3689 15853 3723
rect 15853 3689 15887 3723
rect 15887 3689 15896 3723
rect 15844 3680 15896 3689
rect 19432 3680 19484 3732
rect 4252 3612 4304 3664
rect 2504 3587 2556 3596
rect 2504 3553 2513 3587
rect 2513 3553 2547 3587
rect 2547 3553 2556 3587
rect 4436 3587 4488 3596
rect 2504 3544 2556 3553
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 5632 3587 5684 3596
rect 5632 3553 5641 3587
rect 5641 3553 5675 3587
rect 5675 3553 5684 3587
rect 5632 3544 5684 3553
rect 16304 3587 16356 3596
rect 16304 3553 16338 3587
rect 16338 3553 16356 3587
rect 16304 3544 16356 3553
rect 17776 3544 17828 3596
rect 19064 3544 19116 3596
rect 26516 3587 26568 3596
rect 26516 3553 26525 3587
rect 26525 3553 26559 3587
rect 26559 3553 26568 3587
rect 26516 3544 26568 3553
rect 3700 3476 3752 3528
rect 4344 3476 4396 3528
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 7748 3476 7800 3528
rect 14556 3476 14608 3528
rect 18512 3519 18564 3528
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 16396 3340 16448 3392
rect 17776 3340 17828 3392
rect 26792 3340 26844 3392
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 3884 3136 3936 3188
rect 5632 3136 5684 3188
rect 13268 3179 13320 3188
rect 13268 3145 13277 3179
rect 13277 3145 13311 3179
rect 13311 3145 13320 3179
rect 13268 3136 13320 3145
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 16304 3136 16356 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 18788 3179 18840 3188
rect 18788 3145 18797 3179
rect 18797 3145 18831 3179
rect 18831 3145 18840 3179
rect 18788 3136 18840 3145
rect 18972 3179 19024 3188
rect 18972 3145 18981 3179
rect 18981 3145 19015 3179
rect 19015 3145 19024 3179
rect 18972 3136 19024 3145
rect 4344 3068 4396 3120
rect 4436 3068 4488 3120
rect 5724 3068 5776 3120
rect 16396 3068 16448 3120
rect 18512 3068 18564 3120
rect 2780 3000 2832 3052
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 19064 3000 19116 3052
rect 3148 2932 3200 2984
rect 5172 2932 5224 2984
rect 8300 2932 8352 2984
rect 13268 2932 13320 2984
rect 14464 2932 14516 2984
rect 17960 2932 18012 2984
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 21548 3136 21600 3188
rect 26516 3136 26568 3188
rect 23664 2975 23716 2984
rect 23664 2941 23673 2975
rect 23673 2941 23707 2975
rect 23707 2941 23716 2975
rect 23664 2932 23716 2941
rect 26332 2975 26384 2984
rect 26332 2941 26341 2975
rect 26341 2941 26375 2975
rect 26375 2941 26384 2975
rect 26332 2932 26384 2941
rect 27436 2975 27488 2984
rect 27436 2941 27445 2975
rect 27445 2941 27479 2975
rect 27479 2941 27488 2975
rect 27436 2932 27488 2941
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 2872 2839 2924 2848
rect 2872 2805 2881 2839
rect 2881 2805 2915 2839
rect 2915 2805 2924 2839
rect 2872 2796 2924 2805
rect 10600 2864 10652 2916
rect 13452 2864 13504 2916
rect 14924 2864 14976 2916
rect 18788 2864 18840 2916
rect 20628 2864 20680 2916
rect 24860 2864 24912 2916
rect 5356 2796 5408 2848
rect 26516 2839 26568 2848
rect 26516 2805 26525 2839
rect 26525 2805 26559 2839
rect 26559 2805 26568 2839
rect 26516 2796 26568 2805
rect 27620 2839 27672 2848
rect 27620 2805 27629 2839
rect 27629 2805 27663 2839
rect 27663 2805 27672 2839
rect 27620 2796 27672 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 2596 2592 2648 2644
rect 1492 2499 1544 2508
rect 1492 2465 1501 2499
rect 1501 2465 1535 2499
rect 1535 2465 1544 2499
rect 1492 2456 1544 2465
rect 2044 2456 2096 2508
rect 5356 2592 5408 2644
rect 5816 2567 5868 2576
rect 5816 2533 5825 2567
rect 5825 2533 5859 2567
rect 5859 2533 5868 2567
rect 5816 2524 5868 2533
rect 4988 2456 5040 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 11520 2592 11572 2644
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 19064 2635 19116 2644
rect 19064 2601 19073 2635
rect 19073 2601 19107 2635
rect 19107 2601 19116 2635
rect 19064 2592 19116 2601
rect 21732 2592 21784 2644
rect 13728 2524 13780 2576
rect 12440 2456 12492 2508
rect 15292 2456 15344 2508
rect 18604 2567 18656 2576
rect 18604 2533 18613 2567
rect 18613 2533 18647 2567
rect 18647 2533 18656 2567
rect 18604 2524 18656 2533
rect 19340 2456 19392 2508
rect 24032 2592 24084 2644
rect 25688 2499 25740 2508
rect 25688 2465 25697 2499
rect 25697 2465 25731 2499
rect 25731 2465 25740 2499
rect 25688 2456 25740 2465
rect 4896 2388 4948 2440
rect 6368 2388 6420 2440
rect 12072 2388 12124 2440
rect 17776 2388 17828 2440
rect 19156 2388 19208 2440
rect 22008 2388 22060 2440
rect 23480 2388 23532 2440
rect 2780 2320 2832 2372
rect 1492 2252 1544 2304
rect 6552 2252 6604 2304
rect 25872 2295 25924 2304
rect 25872 2261 25881 2295
rect 25881 2261 25915 2295
rect 25915 2261 25924 2295
rect 25872 2252 25924 2261
rect 29184 2252 29236 2304
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
rect 3516 552 3568 604
rect 7288 552 7340 604
<< metal2 >>
rect 2778 23624 2834 23633
rect 2778 23559 2834 23568
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17746 1808 18226
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1688 17338 1716 17614
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1122 16416 1178 16425
rect 1122 16351 1178 16360
rect 1136 14890 1164 16351
rect 1412 15026 1440 17274
rect 1780 16998 1808 17682
rect 1964 17134 1992 18566
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 2056 17202 2084 18022
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1780 16182 1808 16934
rect 1860 16516 1912 16522
rect 1860 16458 1912 16464
rect 1872 16250 1900 16458
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1768 16176 1820 16182
rect 1768 16118 1820 16124
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1400 15020 1452 15026
rect 1452 14980 1532 15008
rect 1400 14962 1452 14968
rect 1124 14884 1176 14890
rect 1124 14826 1176 14832
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 13870 1440 14214
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1504 13394 1532 14980
rect 1688 14958 1716 15302
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1688 14618 1716 14894
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 2042 14104 2098 14113
rect 2042 14039 2098 14048
rect 2056 13870 2084 14039
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1504 12714 1532 13330
rect 2148 12986 2176 18838
rect 2608 18766 2636 19110
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2608 18290 2636 18702
rect 2596 18284 2648 18290
rect 2596 18226 2648 18232
rect 2596 18080 2648 18086
rect 2792 18068 2820 23559
rect 7470 23520 7526 24000
rect 22466 23520 22522 24000
rect 24950 23624 25006 23633
rect 24950 23559 25006 23568
rect 3054 23080 3110 23089
rect 3054 23015 3110 23024
rect 3068 22166 3096 23015
rect 3422 22400 3478 22409
rect 3422 22335 3478 22344
rect 3436 22234 3464 22335
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 3056 22160 3108 22166
rect 3056 22102 3108 22108
rect 4342 21856 4398 21865
rect 4342 21791 4398 21800
rect 2962 21312 3018 21321
rect 2962 21247 3018 21256
rect 2976 20806 3004 21247
rect 2964 20800 3016 20806
rect 2964 20742 3016 20748
rect 3330 20632 3386 20641
rect 3330 20567 3386 20576
rect 2870 20088 2926 20097
rect 2870 20023 2926 20032
rect 2648 18040 2820 18068
rect 2596 18022 2648 18028
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2424 15706 2452 16594
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2424 14618 2452 15506
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2332 12986 2360 13330
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 1492 12708 1544 12714
rect 1492 12650 1544 12656
rect 1504 12306 1532 12650
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1596 11665 1624 12582
rect 2332 12442 2360 12922
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1582 11656 1638 11665
rect 1582 11591 1638 11600
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 10441 1624 11494
rect 1688 11354 1716 12242
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1688 10810 1716 11290
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1582 10432 1638 10441
rect 1582 10367 1638 10376
rect 1674 10024 1730 10033
rect 1674 9959 1730 9968
rect 1688 9926 1716 9959
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9518 1716 9862
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 2042 9072 2098 9081
rect 1676 9036 1728 9042
rect 2148 9042 2176 9522
rect 2042 9007 2098 9016
rect 2136 9036 2188 9042
rect 1676 8978 1728 8984
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 8673 1624 8774
rect 1582 8664 1638 8673
rect 1582 8599 1638 8608
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 662 7848 718 7857
rect 662 7783 718 7792
rect 676 480 704 7783
rect 1596 7449 1624 8502
rect 1688 8090 1716 8978
rect 2056 8634 2084 9007
rect 2136 8978 2188 8984
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2056 8430 2084 8570
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1582 7440 1638 7449
rect 1582 7375 1638 7384
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 2042 7304 2098 7313
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6905 1624 7142
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1398 6760 1454 6769
rect 1398 6695 1454 6704
rect 1412 6254 1440 6695
rect 1964 6662 1992 7278
rect 2042 7239 2044 7248
rect 2096 7239 2098 7248
rect 2044 7210 2096 7216
rect 2134 7168 2190 7177
rect 2134 7103 2190 7112
rect 2148 6866 2176 7103
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1596 6361 1624 6598
rect 1582 6352 1638 6361
rect 1582 6287 1638 6296
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5914 1440 6190
rect 1964 6186 1992 6598
rect 2148 6458 2176 6802
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 1952 6180 2004 6186
rect 1952 6122 2004 6128
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1596 5681 1624 6054
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1596 5030 1624 5063
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1964 4554 1992 6122
rect 2042 5128 2098 5137
rect 2042 5063 2044 5072
rect 2096 5063 2098 5072
rect 2044 5034 2096 5040
rect 1492 4548 1544 4554
rect 1492 4490 1544 4496
rect 1952 4548 2004 4554
rect 1952 4490 2004 4496
rect 1400 4480 1452 4486
rect 1400 4422 1452 4428
rect 1412 3369 1440 4422
rect 1504 4078 1532 4490
rect 2332 4162 2360 11018
rect 2424 9194 2452 14010
rect 2608 11665 2636 18022
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 17202 2728 17478
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2700 16250 2728 16662
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2884 15978 2912 20023
rect 3146 18320 3202 18329
rect 3146 18255 3202 18264
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3068 18086 3096 18158
rect 3056 18080 3108 18086
rect 3054 18048 3056 18057
rect 3108 18048 3110 18057
rect 3054 17983 3110 17992
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2976 16590 3004 17138
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2964 16176 3016 16182
rect 2964 16118 3016 16124
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 2792 14090 2820 15574
rect 2976 15502 3004 16118
rect 3160 16046 3188 18255
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2976 15162 3004 15438
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2700 14074 2820 14090
rect 2688 14068 2820 14074
rect 2740 14062 2820 14068
rect 2688 14010 2740 14016
rect 2884 13938 2912 14486
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2976 13938 3004 14350
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2780 13864 2832 13870
rect 2778 13832 2780 13841
rect 2832 13832 2834 13841
rect 2778 13767 2834 13776
rect 2884 13705 2912 13874
rect 2870 13696 2926 13705
rect 2870 13631 2926 13640
rect 2884 12889 2912 13631
rect 2976 13530 3004 13874
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 3252 13190 3280 13738
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 2870 12880 2926 12889
rect 2870 12815 2926 12824
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2700 12306 2728 12650
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2700 11898 2728 12242
rect 2792 12102 2820 12310
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2594 11656 2650 11665
rect 2594 11591 2650 11600
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11354 2544 11494
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2516 10810 2544 11290
rect 2792 11150 2820 12038
rect 3252 11914 3280 13126
rect 3068 11886 3280 11914
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2608 10742 2636 11086
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 3068 10690 3096 11886
rect 3344 11642 3372 20567
rect 4066 19408 4122 19417
rect 4066 19343 4122 19352
rect 3516 18896 3568 18902
rect 3516 18838 3568 18844
rect 3528 18358 3556 18838
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3516 18352 3568 18358
rect 3514 18320 3516 18329
rect 3568 18320 3570 18329
rect 3620 18290 3648 18770
rect 3514 18255 3570 18264
rect 3608 18284 3660 18290
rect 3608 18226 3660 18232
rect 4080 17785 4108 19343
rect 4066 17776 4122 17785
rect 4066 17711 4122 17720
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 3804 17338 3832 17614
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4080 16250 4108 16594
rect 4356 16561 4384 21791
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 7484 20369 7512 23520
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 7470 20360 7526 20369
rect 7470 20295 7526 20304
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 8206 18728 8262 18737
rect 8206 18663 8208 18672
rect 8260 18663 8262 18672
rect 8208 18634 8260 18640
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 8220 18222 8248 18634
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 4448 17542 4476 17682
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 4448 17338 4476 17478
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 4802 17096 4858 17105
rect 4802 17031 4858 17040
rect 5264 17060 5316 17066
rect 4342 16552 4398 16561
rect 4342 16487 4398 16496
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3252 11614 3372 11642
rect 3252 11529 3280 11614
rect 3332 11552 3384 11558
rect 3238 11520 3294 11529
rect 3332 11494 3384 11500
rect 3238 11455 3294 11464
rect 3068 10662 3188 10690
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10266 2820 10406
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2686 9888 2742 9897
rect 2686 9823 2742 9832
rect 2424 9166 2636 9194
rect 2700 9178 2728 9823
rect 2792 9722 2820 10202
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2608 9058 2636 9166
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2504 9036 2556 9042
rect 2608 9030 2820 9058
rect 2504 8978 2556 8984
rect 2516 8362 2544 8978
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2594 8120 2650 8129
rect 2594 8055 2650 8064
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 5914 2452 7686
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2516 6225 2544 6802
rect 2608 6730 2636 8055
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2700 6866 2728 7754
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2502 6216 2558 6225
rect 2502 6151 2558 6160
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2424 5370 2452 5646
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2332 4134 2452 4162
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1398 3360 1454 3369
rect 1398 3295 1454 3304
rect 1504 2514 1532 4014
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 2332 3738 2360 3946
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2424 3641 2452 4134
rect 2516 3913 2544 6054
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2502 3904 2558 3913
rect 2502 3839 2558 3848
rect 2410 3632 2466 3641
rect 2410 3567 2466 3576
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 2689 1624 3334
rect 2516 3194 2544 3538
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1582 2680 1638 2689
rect 1582 2615 1638 2624
rect 1492 2508 1544 2514
rect 1492 2450 1544 2456
rect 1504 2310 1532 2450
rect 1492 2304 1544 2310
rect 1492 2246 1544 2252
rect 1780 1465 1808 2790
rect 2608 2650 2636 5510
rect 2700 4826 2728 5782
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2792 4457 2820 9030
rect 2884 8838 2912 9998
rect 3068 9994 3096 10474
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 6905 2912 8774
rect 2870 6896 2926 6905
rect 2870 6831 2926 6840
rect 2884 6458 2912 6831
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2870 5672 2926 5681
rect 2870 5607 2926 5616
rect 2884 4758 2912 5607
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 2964 4480 3016 4486
rect 2778 4448 2834 4457
rect 2964 4422 3016 4428
rect 2778 4383 2834 4392
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 1766 1456 1822 1465
rect 1766 1391 1822 1400
rect 2056 480 2084 2450
rect 2700 1442 2728 3334
rect 2792 3058 2820 3946
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2792 2378 2820 2994
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2884 2145 2912 2790
rect 2870 2136 2926 2145
rect 2870 2071 2926 2080
rect 2700 1414 2820 1442
rect 662 0 718 480
rect 2042 0 2098 480
rect 2792 377 2820 1414
rect 2976 921 3004 4422
rect 3068 4282 3096 5170
rect 3160 5001 3188 10662
rect 3252 10130 3280 11455
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3252 9722 3280 10066
rect 3344 10062 3372 11494
rect 3436 11286 3464 11698
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3238 9616 3294 9625
rect 3436 9586 3464 9862
rect 3238 9551 3240 9560
rect 3292 9551 3294 9560
rect 3424 9580 3476 9586
rect 3240 9522 3292 9528
rect 3424 9522 3476 9528
rect 3528 7993 3556 15914
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3620 15162 3648 15846
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3790 15328 3846 15337
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3712 15026 3740 15302
rect 3790 15263 3846 15272
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3620 14006 3648 14418
rect 3712 14414 3740 14758
rect 3700 14408 3752 14414
rect 3698 14376 3700 14385
rect 3752 14376 3754 14385
rect 3698 14311 3754 14320
rect 3608 14000 3660 14006
rect 3606 13968 3608 13977
rect 3660 13968 3662 13977
rect 3606 13903 3662 13912
rect 3606 12336 3662 12345
rect 3606 12271 3662 12280
rect 3620 8378 3648 12271
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3712 8498 3740 8774
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3698 8392 3754 8401
rect 3620 8350 3698 8378
rect 3698 8327 3754 8336
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3620 8090 3648 8230
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3514 7984 3570 7993
rect 3514 7919 3570 7928
rect 3240 6248 3292 6254
rect 3238 6216 3240 6225
rect 3292 6216 3294 6225
rect 3238 6151 3294 6160
rect 3146 4992 3202 5001
rect 3146 4927 3202 4936
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3160 3738 3188 4927
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3252 4078 3280 4626
rect 3240 4072 3292 4078
rect 3238 4040 3240 4049
rect 3292 4040 3294 4049
rect 3238 3975 3294 3984
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3160 2990 3188 3674
rect 3712 3534 3740 8327
rect 3804 5953 3832 15263
rect 4080 15162 4108 15574
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 4158 11112 4214 11121
rect 4158 11047 4214 11056
rect 4172 10810 4200 11047
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 3882 9480 3938 9489
rect 3882 9415 3938 9424
rect 3896 8362 3924 9415
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 8430 4108 8910
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 4080 8090 4108 8366
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3896 7206 3924 7822
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3896 6662 3924 7142
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6186 3924 6598
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3790 5944 3846 5953
rect 3790 5879 3846 5888
rect 3988 5234 4016 7142
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4068 5364 4120 5370
rect 4172 5352 4200 5714
rect 4120 5324 4200 5352
rect 4068 5306 4120 5312
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3896 4486 3924 4626
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3896 3194 3924 4422
rect 4080 3738 4108 4558
rect 4264 4282 4292 12854
rect 4356 8090 4384 16487
rect 4434 15872 4490 15881
rect 4434 15807 4490 15816
rect 4448 10810 4476 15807
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4632 13433 4660 14962
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4724 14074 4752 14486
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4618 13424 4674 13433
rect 4618 13359 4674 13368
rect 4816 12986 4844 17031
rect 5264 17002 5316 17008
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4816 12782 4844 12922
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4620 10600 4672 10606
rect 4618 10568 4620 10577
rect 4672 10568 4674 10577
rect 4618 10503 4674 10512
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4356 7546 4384 8026
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4632 7449 4660 7958
rect 4724 7886 4752 8230
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4618 7440 4674 7449
rect 4618 7375 4620 7384
rect 4672 7375 4674 7384
rect 4620 7346 4672 7352
rect 4632 7177 4660 7346
rect 4724 7206 4752 7822
rect 4712 7200 4764 7206
rect 4618 7168 4674 7177
rect 4712 7142 4764 7148
rect 4618 7103 4674 7112
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4540 5098 4568 5646
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4448 4282 4476 5034
rect 4540 4826 4568 5034
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4632 4622 4660 5170
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4264 4078 4292 4218
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4264 3670 4292 4014
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 4356 3126 4384 3470
rect 4448 3126 4476 3538
rect 4632 3534 4660 4082
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4632 3058 4660 3470
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 4908 2530 4936 16934
rect 5276 16726 5304 17002
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5368 16794 5396 16934
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5264 16720 5316 16726
rect 5264 16662 5316 16668
rect 5460 16658 5488 17206
rect 5552 17202 5580 17478
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5552 16726 5580 17138
rect 7668 16998 7696 17614
rect 7760 17338 7788 17682
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5460 16182 5488 16594
rect 5552 16250 5580 16662
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 5000 12424 5028 15982
rect 5460 15570 5488 16118
rect 6840 15638 6868 16390
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5460 14958 5488 15506
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 6288 15162 6316 15574
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6288 15026 6316 15098
rect 6644 15088 6696 15094
rect 6644 15030 6696 15036
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 14618 5212 14758
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5460 14482 5488 14894
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5448 14476 5500 14482
rect 5368 14436 5448 14464
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 13802 5120 14214
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5092 12986 5120 13738
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5000 12396 5120 12424
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5000 11898 5028 12242
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5092 11778 5120 12396
rect 5184 12209 5212 13670
rect 5368 13258 5396 14436
rect 5448 14418 5500 14424
rect 5552 14346 5580 14758
rect 5722 14648 5778 14657
rect 5722 14583 5778 14592
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5460 13938 5488 14214
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5644 13734 5672 14350
rect 5632 13728 5684 13734
rect 5552 13688 5632 13716
rect 5552 13326 5580 13688
rect 5632 13670 5684 13676
rect 5736 13530 5764 14583
rect 6288 14482 6316 14962
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5630 13424 5686 13433
rect 5630 13359 5632 13368
rect 5684 13359 5686 13368
rect 5632 13330 5684 13336
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12850 5488 13126
rect 5552 12850 5580 13262
rect 5644 12918 5672 13330
rect 5736 12986 5764 13466
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5170 12200 5226 12209
rect 5170 12135 5226 12144
rect 5000 11750 5120 11778
rect 5264 11824 5316 11830
rect 5264 11766 5316 11772
rect 5000 6338 5028 11750
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5092 10810 5120 11154
rect 5276 11150 5304 11766
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5184 10538 5212 11086
rect 5276 10674 5304 11086
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5184 10266 5212 10474
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5276 10198 5304 10610
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5092 9722 5120 10066
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5184 9382 5212 9522
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5000 6310 5120 6338
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 5000 5710 5028 6122
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 5370 5028 5646
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5092 5166 5120 6310
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5092 3505 5120 3878
rect 5078 3496 5134 3505
rect 5078 3431 5134 3440
rect 5184 2990 5212 9318
rect 5368 8945 5396 12718
rect 5736 12306 5764 12786
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10674 5764 10950
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5540 10600 5592 10606
rect 5460 10548 5540 10554
rect 5460 10542 5592 10548
rect 5460 10526 5580 10542
rect 5460 9874 5488 10526
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 10033 5580 10406
rect 5736 10282 5764 10610
rect 5828 10606 5856 14282
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 6288 13326 6316 14418
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6472 14113 6500 14282
rect 6458 14104 6514 14113
rect 6564 14074 6592 14554
rect 6458 14039 6514 14048
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 6288 12986 6316 13262
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6380 12442 6408 13874
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6472 12458 6500 12854
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6463 12430 6500 12458
rect 6463 12356 6491 12430
rect 6463 12328 6500 12356
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 6288 11762 6316 12106
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5644 10254 5764 10282
rect 5644 10062 5672 10254
rect 5632 10056 5684 10062
rect 5538 10024 5594 10033
rect 5632 9998 5684 10004
rect 5538 9959 5594 9968
rect 5460 9846 5580 9874
rect 5354 8936 5410 8945
rect 5354 8871 5410 8880
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5368 5642 5396 6054
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5368 5273 5396 5578
rect 5460 5370 5488 5714
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5354 5264 5410 5273
rect 5354 5199 5410 5208
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 4146 5488 4558
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5368 2854 5396 2885
rect 5356 2848 5408 2854
rect 5552 2802 5580 9846
rect 5644 9450 5672 9998
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5828 9722 5856 9862
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5724 9648 5776 9654
rect 6472 9636 6500 12328
rect 6656 10266 6684 15030
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14550 6868 14758
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6840 9654 6868 10202
rect 7024 10062 7052 14826
rect 7196 14816 7248 14822
rect 7194 14784 7196 14793
rect 7248 14784 7250 14793
rect 7194 14719 7250 14728
rect 7208 14618 7236 14719
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7116 12986 7144 13330
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7208 10266 7236 14554
rect 7576 14414 7604 15302
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7300 12238 7328 12269
rect 7288 12232 7340 12238
rect 7286 12200 7288 12209
rect 7340 12200 7342 12209
rect 7286 12135 7342 12144
rect 7300 11898 7328 12135
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7668 11694 7696 16934
rect 8312 16658 8340 22170
rect 15660 22160 15712 22166
rect 15660 22102 15712 22108
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8588 17678 8616 18090
rect 9600 18086 9628 18770
rect 9772 18760 9824 18766
rect 9770 18728 9772 18737
rect 9824 18728 9826 18737
rect 9770 18663 9826 18672
rect 11794 18728 11850 18737
rect 11794 18663 11850 18672
rect 9784 18154 9812 18663
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 8576 17672 8628 17678
rect 8496 17620 8576 17626
rect 8496 17614 8628 17620
rect 9310 17640 9366 17649
rect 8496 17598 8616 17614
rect 8496 17270 8524 17598
rect 9310 17575 9366 17584
rect 9496 17604 9548 17610
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8116 16584 8168 16590
rect 8496 16572 8524 17206
rect 8588 17134 8616 17478
rect 9324 17241 9352 17575
rect 9496 17546 9548 17552
rect 9310 17232 9366 17241
rect 9310 17167 9366 17176
rect 8576 17128 8628 17134
rect 9508 17105 9536 17546
rect 8576 17070 8628 17076
rect 9494 17096 9550 17105
rect 9494 17031 9550 17040
rect 9600 16998 9628 18022
rect 9784 17678 9812 18090
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 11532 17678 11560 18226
rect 11716 17746 11744 18566
rect 11808 18193 11836 18663
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 12636 18290 12664 18566
rect 15304 18358 15332 18566
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12900 18216 12952 18222
rect 11794 18184 11850 18193
rect 12900 18158 12952 18164
rect 11794 18119 11850 18128
rect 12164 18148 12216 18154
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 9588 16992 9640 16998
rect 9640 16940 9720 16946
rect 9588 16934 9720 16940
rect 8680 16794 8708 16934
rect 9600 16918 9720 16934
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 9496 16720 9548 16726
rect 8666 16688 8722 16697
rect 9496 16662 9548 16668
rect 8666 16623 8668 16632
rect 8720 16623 8722 16632
rect 8668 16594 8720 16600
rect 8576 16584 8628 16590
rect 8496 16544 8576 16572
rect 8116 16526 8168 16532
rect 8576 16526 8628 16532
rect 8128 15910 8156 16526
rect 8588 16250 8616 16526
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8680 16182 8708 16594
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8128 15473 8156 15846
rect 8114 15464 8170 15473
rect 8114 15399 8170 15408
rect 8312 14362 8340 15846
rect 8220 14334 8340 14362
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8128 13802 8156 14214
rect 8220 13841 8248 14334
rect 8206 13832 8262 13841
rect 8116 13796 8168 13802
rect 8206 13767 8262 13776
rect 8116 13738 8168 13744
rect 8128 12850 8156 13738
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7944 12442 7972 12650
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7760 11898 7788 12378
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7852 11558 7880 12242
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 7944 11830 7972 12038
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7944 11694 7972 11766
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7852 11286 7880 11494
rect 8036 11354 8064 11562
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 6828 9648 6880 9654
rect 6472 9608 6592 9636
rect 5724 9590 5776 9596
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5630 3632 5686 3641
rect 5630 3567 5632 3576
rect 5684 3567 5686 3576
rect 5632 3538 5684 3544
rect 5644 3194 5672 3538
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5736 3126 5764 9590
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6288 8276 6316 8434
rect 6380 8401 6408 9318
rect 6564 8498 6592 9608
rect 7024 9602 7052 9998
rect 6828 9590 6880 9596
rect 6932 9574 7052 9602
rect 6644 9512 6696 9518
rect 6932 9500 6960 9574
rect 6644 9454 6696 9460
rect 6840 9472 6960 9500
rect 6656 8974 6684 9454
rect 6840 9382 6868 9472
rect 7116 9466 7144 9998
rect 7024 9450 7144 9466
rect 7012 9444 7144 9450
rect 7064 9438 7144 9444
rect 7012 9386 7064 9392
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6840 9217 6868 9318
rect 6826 9208 6882 9217
rect 6826 9143 6882 9152
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6656 8430 6684 8910
rect 7024 8838 7052 9386
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8634 7052 8774
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6644 8424 6696 8430
rect 6366 8392 6422 8401
rect 6644 8366 6696 8372
rect 6366 8327 6422 8336
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6288 8248 6408 8276
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 6288 7546 6316 7890
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 6380 3505 6408 8248
rect 6564 7546 6592 8298
rect 6656 8294 6684 8366
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7750 6684 8230
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6564 6730 6592 7482
rect 6656 7410 6684 7686
rect 7286 7576 7342 7585
rect 7286 7511 7342 7520
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6564 6390 6592 6666
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6552 4616 6604 4622
rect 6656 4604 6684 7346
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 6769 6868 6802
rect 6920 6792 6972 6798
rect 6826 6760 6882 6769
rect 6920 6734 6972 6740
rect 6826 6695 6882 6704
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6604 4576 6684 4604
rect 6552 4558 6604 4564
rect 6564 3942 6592 4558
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6366 3496 6422 3505
rect 6366 3431 6422 3440
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5408 2796 5580 2802
rect 5356 2790 5580 2796
rect 5368 2774 5580 2790
rect 5814 2816 5870 2825
rect 5368 2650 5396 2774
rect 5814 2751 5870 2760
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5828 2582 5856 2751
rect 5816 2576 5868 2582
rect 4908 2514 5028 2530
rect 5816 2518 5868 2524
rect 4908 2508 5040 2514
rect 4908 2502 4988 2508
rect 4988 2450 5040 2456
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 2962 912 3018 921
rect 2962 847 3018 856
rect 3516 604 3568 610
rect 3516 546 3568 552
rect 3528 480 3556 546
rect 4908 480 4936 2382
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 6380 480 6408 2382
rect 6564 2310 6592 3878
rect 6748 2666 6776 6598
rect 6840 6458 6868 6695
rect 6932 6458 6960 6734
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6932 5914 6960 6394
rect 7024 6322 7052 7210
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7024 5914 7052 6258
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7024 5030 7052 5646
rect 7102 5264 7158 5273
rect 7102 5199 7158 5208
rect 7012 5024 7064 5030
rect 7010 4992 7012 5001
rect 7064 4992 7066 5001
rect 7010 4927 7066 4936
rect 7116 4690 7144 5199
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7116 4282 7144 4626
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 6748 2638 6960 2666
rect 6932 2514 6960 2638
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 7300 610 7328 7511
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 6254 7420 6598
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 5914 7420 6190
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7576 5370 7604 6122
rect 8022 5944 8078 5953
rect 8022 5879 8024 5888
rect 8076 5879 8078 5888
rect 8024 5850 8076 5856
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7944 5545 7972 5646
rect 7930 5536 7986 5545
rect 7930 5471 7986 5480
rect 8036 5370 8064 5850
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8036 4282 8064 5034
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7288 604 7340 610
rect 7288 546 7340 552
rect 7760 480 7788 3470
rect 8128 3074 8156 12038
rect 8220 6497 8248 13767
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8496 12714 8524 13330
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8404 9625 8432 11562
rect 8390 9616 8446 9625
rect 8390 9551 8446 9560
rect 8680 6633 8708 16118
rect 9140 15706 9168 16526
rect 9508 16250 9536 16662
rect 9692 16590 9720 16918
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9784 16436 9812 17614
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10060 17202 10088 17478
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10060 16794 10088 17138
rect 10336 17066 10364 17478
rect 11532 17338 11560 17614
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11716 17270 11744 17682
rect 11704 17264 11756 17270
rect 11610 17232 11666 17241
rect 11704 17206 11756 17212
rect 11610 17167 11666 17176
rect 10324 17060 10376 17066
rect 10324 17002 10376 17008
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 9692 16408 9812 16436
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9692 15502 9720 16408
rect 10336 16250 10364 16526
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 15706 9996 15846
rect 10520 15706 10548 16050
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9692 15178 9720 15438
rect 9600 15162 9720 15178
rect 9784 15162 9812 15506
rect 9588 15156 9720 15162
rect 9640 15150 9720 15156
rect 9772 15156 9824 15162
rect 9588 15098 9640 15104
rect 9772 15098 9824 15104
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 9324 14822 9352 15030
rect 9404 14952 9456 14958
rect 9586 14920 9642 14929
rect 9456 14900 9586 14906
rect 9404 14894 9586 14900
rect 9416 14878 9586 14894
rect 9586 14855 9642 14864
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14278 9352 14758
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8864 13977 8892 14010
rect 8850 13968 8906 13977
rect 8850 13903 8906 13912
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9048 13190 9076 13738
rect 9508 13530 9536 14418
rect 9784 14346 9812 15098
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9876 14929 9904 15030
rect 9862 14920 9918 14929
rect 9862 14855 9918 14864
rect 9968 14618 9996 15642
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 10060 14074 10088 14418
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10060 13977 10088 14010
rect 10046 13968 10102 13977
rect 10046 13903 10102 13912
rect 9588 13728 9640 13734
rect 10152 13705 10180 14350
rect 10244 14006 10272 14962
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10612 14521 10640 14554
rect 10598 14512 10654 14521
rect 10598 14447 10654 14456
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10336 14074 10364 14282
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 9588 13670 9640 13676
rect 10138 13696 10194 13705
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 12646 9076 13126
rect 9600 12968 9628 13670
rect 10138 13631 10194 13640
rect 10152 13190 10180 13631
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 9680 12980 9732 12986
rect 9600 12940 9680 12968
rect 9680 12922 9732 12928
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9048 12238 9076 12582
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9048 11898 9076 12174
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9232 10713 9260 12650
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9600 11762 9628 12106
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9692 11694 9720 12038
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 11354 9536 11494
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9968 11082 9996 12174
rect 10612 11558 10640 12242
rect 10600 11552 10652 11558
rect 10598 11520 10600 11529
rect 10652 11520 10654 11529
rect 10598 11455 10654 11464
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9218 10704 9274 10713
rect 9218 10639 9274 10648
rect 9588 10668 9640 10674
rect 9232 9518 9260 10639
rect 9588 10610 9640 10616
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9518 9352 9862
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 7954 9076 9318
rect 9232 9178 9260 9454
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9324 8566 9352 9454
rect 9508 9081 9536 10406
rect 9600 9518 9628 10610
rect 9968 9897 9996 11018
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 10266 10088 10406
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9954 9888 10010 9897
rect 9954 9823 10010 9832
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9494 9072 9550 9081
rect 9494 9007 9550 9016
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9862 7984 9918 7993
rect 9036 7948 9088 7954
rect 9862 7919 9918 7928
rect 9036 7890 9088 7896
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 7002 9168 7278
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 8666 6624 8722 6633
rect 8666 6559 8722 6568
rect 8206 6488 8262 6497
rect 8206 6423 8262 6432
rect 8220 5030 8248 6423
rect 9600 6322 9628 7210
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9600 6066 9628 6258
rect 9508 6038 9628 6066
rect 9508 5710 9536 6038
rect 9588 5908 9640 5914
rect 9692 5896 9720 6938
rect 9770 6760 9826 6769
rect 9770 6695 9772 6704
rect 9824 6695 9826 6704
rect 9772 6666 9824 6672
rect 9770 6624 9826 6633
rect 9770 6559 9826 6568
rect 9640 5868 9720 5896
rect 9588 5850 9640 5856
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 8574 5400 8630 5409
rect 9508 5370 9536 5646
rect 8574 5335 8576 5344
rect 8628 5335 8630 5344
rect 9496 5364 9548 5370
rect 8576 5306 8628 5312
rect 9496 5306 9548 5312
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 9784 4808 9812 6559
rect 9876 6254 9904 7919
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9968 5137 9996 9823
rect 10060 9178 10088 10202
rect 10336 10198 10364 10950
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10428 10470 10456 10542
rect 10416 10464 10468 10470
rect 10612 10418 10640 11455
rect 10416 10406 10468 10412
rect 10520 10390 10640 10418
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10336 9722 10364 10134
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 10232 8424 10284 8430
rect 10284 8372 10364 8378
rect 10232 8366 10364 8372
rect 10060 7954 10088 8366
rect 10244 8350 10364 8366
rect 10336 8022 10364 8350
rect 10324 8016 10376 8022
rect 10322 7984 10324 7993
rect 10376 7984 10378 7993
rect 10048 7948 10100 7954
rect 10322 7919 10378 7928
rect 10048 7890 10100 7896
rect 10336 7342 10364 7919
rect 10520 7886 10548 10390
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10612 9450 10640 9998
rect 10704 9518 10732 16934
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 11624 16794 11652 17167
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11624 16250 11652 16730
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11624 16153 11652 16186
rect 11610 16144 11666 16153
rect 11610 16079 11666 16088
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 14958 10916 15982
rect 11716 15910 11744 16594
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 10796 14521 10824 14758
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 11348 14657 11376 14758
rect 11334 14648 11390 14657
rect 11334 14583 11336 14592
rect 11388 14583 11390 14592
rect 11336 14554 11388 14560
rect 11348 14523 11376 14554
rect 10782 14512 10838 14521
rect 10782 14447 10838 14456
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11716 13569 11744 15846
rect 11702 13560 11758 13569
rect 11702 13495 11758 13504
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 11132 10824 13126
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11354 10916 11494
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 10876 11348 10928 11354
rect 10928 11308 11100 11336
rect 10876 11290 10928 11296
rect 10888 11225 10916 11290
rect 10968 11144 11020 11150
rect 10796 11104 10916 11132
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10796 10130 10824 10610
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10612 9042 10640 9386
rect 10690 9208 10746 9217
rect 10690 9143 10746 9152
rect 10704 9110 10732 9143
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10612 8362 10640 8978
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10428 6798 10456 7142
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10416 6792 10468 6798
rect 10888 6769 10916 11104
rect 10968 11086 11020 11092
rect 10980 10674 11008 11086
rect 11072 10810 11100 11308
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 11348 10577 11376 10950
rect 11334 10568 11390 10577
rect 11334 10503 11390 10512
rect 11518 10568 11574 10577
rect 11518 10503 11574 10512
rect 11348 10470 11376 10503
rect 11336 10464 11388 10470
rect 11334 10432 11336 10441
rect 11388 10432 11390 10441
rect 10956 10364 11252 10384
rect 11334 10367 11390 10376
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 11532 10033 11560 10503
rect 11518 10024 11574 10033
rect 11336 9988 11388 9994
rect 11518 9959 11574 9968
rect 11336 9930 11388 9936
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 11348 9178 11376 9930
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 11440 8090 11468 8910
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 10416 6734 10468 6740
rect 10874 6760 10930 6769
rect 10152 6458 10180 6734
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10428 6390 10456 6734
rect 10874 6695 10930 6704
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10506 6352 10562 6361
rect 10506 6287 10562 6296
rect 11336 6316 11388 6322
rect 10520 6186 10548 6287
rect 11336 6258 11388 6264
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10060 5710 10088 6122
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 10048 5704 10100 5710
rect 10046 5672 10048 5681
rect 10100 5672 10102 5681
rect 10046 5607 10102 5616
rect 9954 5128 10010 5137
rect 9954 5063 10010 5072
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 11348 4826 11376 6258
rect 9692 4780 9812 4808
rect 11336 4820 11388 4826
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8220 4214 8248 4422
rect 8208 4208 8260 4214
rect 9692 4162 9720 4780
rect 11336 4762 11388 4768
rect 10140 4752 10192 4758
rect 10140 4694 10192 4700
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9784 4282 9812 4626
rect 10152 4321 10180 4694
rect 10138 4312 10194 4321
rect 9772 4276 9824 4282
rect 10138 4247 10140 4256
rect 9772 4218 9824 4224
rect 10192 4247 10194 4256
rect 10140 4218 10192 4224
rect 8208 4150 8260 4156
rect 9600 4134 9720 4162
rect 9600 4078 9628 4134
rect 9588 4072 9640 4078
rect 8390 4040 8446 4049
rect 9588 4014 9640 4020
rect 8390 3975 8392 3984
rect 8444 3975 8446 3984
rect 8392 3946 8444 3952
rect 8404 3738 8432 3946
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8128 3046 8340 3074
rect 8312 2990 8340 3046
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 9218 2816 9274 2825
rect 9218 2751 9274 2760
rect 9232 480 9260 2751
rect 10612 480 10640 2858
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 11532 2650 11560 9454
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11716 8090 11744 9114
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11808 6866 11836 18119
rect 12164 18090 12216 18096
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11992 16114 12020 16526
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 12176 15026 12204 18090
rect 12912 17882 12940 18158
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 16114 13400 16390
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12912 15162 12940 15370
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 13004 14890 13032 15438
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 13004 14618 13032 14826
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12176 14006 12204 14418
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 12544 13870 12572 14214
rect 13188 14113 13216 14758
rect 13280 14634 13308 15846
rect 13372 15706 13400 16050
rect 13544 16040 13596 16046
rect 13542 16008 13544 16017
rect 13596 16008 13598 16017
rect 13740 15978 13768 17206
rect 13542 15943 13598 15952
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13740 15094 13768 15506
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 14188 15020 14240 15026
rect 14108 14980 14188 15008
rect 13910 14648 13966 14657
rect 13280 14606 13400 14634
rect 13268 14544 13320 14550
rect 13266 14512 13268 14521
rect 13320 14512 13322 14521
rect 13266 14447 13322 14456
rect 13174 14104 13230 14113
rect 13174 14039 13230 14048
rect 12622 13968 12678 13977
rect 12622 13903 12678 13912
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11992 13394 12020 13738
rect 12254 13696 12310 13705
rect 12254 13631 12310 13640
rect 12268 13462 12296 13631
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11992 12918 12020 13330
rect 12268 12986 12296 13398
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12348 10804 12400 10810
rect 12452 10792 12480 11086
rect 12400 10764 12572 10792
rect 12348 10746 12400 10752
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12256 9376 12308 9382
rect 12360 9353 12388 9862
rect 12256 9318 12308 9324
rect 12346 9344 12402 9353
rect 12268 9042 12296 9318
rect 12346 9279 12402 9288
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11900 8294 11928 8910
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11900 7274 11928 8230
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11624 6118 11652 6802
rect 11808 6458 11836 6802
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11900 6458 11928 6734
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11808 6225 11836 6394
rect 11794 6216 11850 6225
rect 11794 6151 11850 6160
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11624 5914 11652 6054
rect 12268 5914 12296 7346
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12162 5400 12218 5409
rect 12162 5335 12164 5344
rect 12216 5335 12218 5344
rect 12164 5306 12216 5312
rect 12176 4593 12204 5306
rect 12268 5234 12296 5850
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12162 4584 12218 4593
rect 12162 4519 12218 4528
rect 12268 4321 12296 5170
rect 12254 4312 12310 4321
rect 12254 4247 12310 4256
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 12360 2530 12388 8774
rect 12544 8090 12572 10764
rect 12636 9625 12664 13903
rect 13082 13560 13138 13569
rect 13280 13530 13308 14447
rect 13082 13495 13138 13504
rect 13268 13524 13320 13530
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12820 12442 12848 12854
rect 13096 12617 13124 13495
rect 13268 13466 13320 13472
rect 13372 13274 13400 14606
rect 13910 14583 13966 14592
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13832 13705 13860 13942
rect 13818 13696 13874 13705
rect 13818 13631 13874 13640
rect 13280 13246 13400 13274
rect 13082 12608 13138 12617
rect 13082 12543 13138 12552
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12820 11762 12848 12378
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11218 12940 11494
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12912 10810 12940 11154
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12622 9616 12678 9625
rect 12622 9551 12678 9560
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12544 7993 12572 8026
rect 12530 7984 12586 7993
rect 12452 7942 12530 7970
rect 12452 7410 12480 7942
rect 12530 7919 12586 7928
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12636 6866 12664 9551
rect 12728 9110 12756 10066
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9518 12940 9862
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12808 9376 12860 9382
rect 12806 9344 12808 9353
rect 12860 9344 12862 9353
rect 12806 9279 12862 9288
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12728 8090 12756 9046
rect 12820 8906 12848 9279
rect 12912 9178 12940 9454
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13004 9042 13032 9318
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 13096 6746 13124 12543
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13188 9722 13216 9998
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13174 9072 13230 9081
rect 13174 9007 13176 9016
rect 13228 9007 13230 9016
rect 13176 8978 13228 8984
rect 13188 8566 13216 8978
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 13096 6718 13216 6746
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12806 6488 12862 6497
rect 12806 6423 12862 6432
rect 12820 6186 12848 6423
rect 13096 6254 13124 6598
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12530 5536 12586 5545
rect 12530 5471 12586 5480
rect 12544 4826 12572 5471
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12716 4616 12768 4622
rect 12820 4593 12848 5714
rect 12912 4826 12940 6054
rect 13096 5710 13124 6190
rect 13188 5914 13216 6718
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12716 4558 12768 4564
rect 12806 4584 12862 4593
rect 12728 4282 12756 4558
rect 12806 4519 12862 4528
rect 12912 4282 12940 4762
rect 13004 4758 13032 5510
rect 13096 5098 13124 5646
rect 13188 5545 13216 5850
rect 13174 5536 13230 5545
rect 13174 5471 13230 5480
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 13004 4146 13032 4694
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13280 3194 13308 13246
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 12986 13400 13126
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13740 12850 13768 12922
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13740 11626 13768 12786
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13372 8634 13400 9114
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13464 7721 13492 10406
rect 13832 10146 13860 11018
rect 13924 10198 13952 14583
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14016 13705 14044 14418
rect 14108 14278 14136 14980
rect 14188 14962 14240 14968
rect 14188 14816 14240 14822
rect 14186 14784 14188 14793
rect 14240 14784 14242 14793
rect 14186 14719 14242 14728
rect 14292 14634 14320 18090
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15028 17882 15056 18022
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 15016 17876 15068 17882
rect 15212 17864 15240 18022
rect 15016 17818 15068 17824
rect 15120 17836 15240 17864
rect 14660 17134 14688 17818
rect 15120 17542 15148 17836
rect 15304 17762 15332 18294
rect 15474 18184 15530 18193
rect 15474 18119 15476 18128
rect 15528 18119 15530 18128
rect 15476 18090 15528 18096
rect 15212 17746 15332 17762
rect 15200 17740 15332 17746
rect 15252 17734 15332 17740
rect 15200 17682 15252 17688
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 14922 17232 14978 17241
rect 15120 17202 15148 17478
rect 14922 17167 14924 17176
rect 14976 17167 14978 17176
rect 15108 17196 15160 17202
rect 14924 17138 14976 17144
rect 15108 17138 15160 17144
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 15212 16998 15240 17682
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15304 17082 15332 17614
rect 15566 17096 15622 17105
rect 15304 17054 15424 17082
rect 15396 16998 15424 17054
rect 15566 17031 15622 17040
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 14752 16794 14780 16934
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15028 16250 15056 16526
rect 15212 16522 15240 16934
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14200 14606 14320 14634
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14108 14074 14136 14214
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14002 13696 14058 13705
rect 14002 13631 14058 13640
rect 14200 11642 14228 14606
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 12782 14320 13126
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14384 12442 14412 12718
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14016 11614 14228 11642
rect 14016 10441 14044 11614
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14002 10432 14058 10441
rect 14002 10367 14058 10376
rect 13740 10118 13860 10146
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 13740 10062 13768 10118
rect 14108 10062 14136 11494
rect 14372 10736 14424 10742
rect 14370 10704 14372 10713
rect 14424 10704 14426 10713
rect 14370 10639 14426 10648
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14016 9722 14044 9998
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14108 9586 14136 9998
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 9178 14044 9318
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14108 8634 14136 9522
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14200 8945 14228 9318
rect 14186 8936 14242 8945
rect 14186 8871 14242 8880
rect 14200 8838 14228 8871
rect 14292 8838 14320 10134
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13450 7712 13506 7721
rect 13450 7647 13506 7656
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13372 6322 13400 6666
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13360 6112 13412 6118
rect 13358 6080 13360 6089
rect 13412 6080 13414 6089
rect 13358 6015 13414 6024
rect 13464 5574 13492 6802
rect 13924 6798 13952 7142
rect 13820 6792 13872 6798
rect 13818 6760 13820 6769
rect 13912 6792 13964 6798
rect 13872 6760 13874 6769
rect 13912 6734 13964 6740
rect 13818 6695 13874 6704
rect 13832 6322 13860 6695
rect 13924 6458 13952 6734
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13464 4049 13492 5510
rect 14200 5137 14228 8774
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14186 5128 14242 5137
rect 14186 5063 14242 5072
rect 14384 4622 14412 5238
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14384 4282 14412 4558
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 13450 4040 13506 4049
rect 13450 3975 13506 3984
rect 14476 3194 14504 12650
rect 14568 12345 14596 14894
rect 14554 12336 14610 12345
rect 14554 12271 14610 12280
rect 14646 10024 14702 10033
rect 14646 9959 14648 9968
rect 14700 9959 14702 9968
rect 14648 9930 14700 9936
rect 14660 9518 14688 9930
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14752 9178 14780 9522
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 4078 14596 5510
rect 14556 4072 14608 4078
rect 14660 4049 14688 8774
rect 15028 7449 15056 16186
rect 15212 15366 15240 16458
rect 15200 15360 15252 15366
rect 15120 15308 15200 15314
rect 15120 15302 15252 15308
rect 15120 15286 15240 15302
rect 15120 15026 15148 15286
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15212 12866 15240 13942
rect 15382 13696 15438 13705
rect 15382 13631 15438 13640
rect 15120 12838 15240 12866
rect 15120 12782 15148 12838
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15396 10266 15424 13631
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15488 12986 15516 13330
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15580 12918 15608 17031
rect 15672 16726 15700 22102
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 15750 18864 15806 18873
rect 15750 18799 15806 18808
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15672 15910 15700 16662
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15764 14618 15792 18799
rect 17682 18592 17738 18601
rect 15956 18524 16252 18544
rect 17682 18527 17738 18536
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 16394 17368 16450 17377
rect 16394 17303 16450 17312
rect 15842 17232 15898 17241
rect 15842 17167 15898 17176
rect 15856 16046 15884 17167
rect 15934 17096 15990 17105
rect 15934 17031 15990 17040
rect 15948 16794 15976 17031
rect 16304 16992 16356 16998
rect 16408 16969 16436 17303
rect 16304 16934 16356 16940
rect 16394 16960 16450 16969
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15856 15706 15884 15982
rect 16316 15978 16344 16934
rect 16394 16895 16450 16904
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15856 15502 15884 15642
rect 16316 15502 16344 15914
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 16394 14784 16450 14793
rect 16394 14719 16450 14728
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 13870 15700 14214
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 16316 14074 16344 14554
rect 16408 14113 16436 14719
rect 16394 14104 16450 14113
rect 16304 14068 16356 14074
rect 16394 14039 16450 14048
rect 16304 14010 16356 14016
rect 15750 13968 15806 13977
rect 16408 13954 16436 14039
rect 15750 13903 15752 13912
rect 15804 13903 15806 13912
rect 15844 13932 15896 13938
rect 15752 13874 15804 13880
rect 15844 13874 15896 13880
rect 16316 13926 16436 13954
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 15580 12442 15608 12650
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15764 12374 15792 13330
rect 15856 13326 15884 13874
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15856 12442 15884 13262
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 16316 12186 16344 13926
rect 15672 12158 16344 12186
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15396 9654 15424 10202
rect 15672 10130 15700 12158
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 16394 11928 16450 11937
rect 16394 11863 16450 11872
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15856 11286 15884 11698
rect 16408 11694 16436 11863
rect 16500 11801 16528 12038
rect 16486 11792 16542 11801
rect 16486 11727 16542 11736
rect 16500 11694 16528 11727
rect 16396 11688 16448 11694
rect 16302 11656 16358 11665
rect 16396 11630 16448 11636
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16302 11591 16304 11600
rect 16356 11591 16358 11600
rect 16304 11562 16356 11568
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15856 10810 15884 11222
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 16408 10674 16436 11494
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15014 7440 15070 7449
rect 15014 7375 15070 7384
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15212 7206 15240 7346
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15028 5574 15056 6734
rect 15212 6322 15240 7142
rect 15304 6798 15332 8298
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15212 5896 15240 6258
rect 15396 5930 15424 9590
rect 15672 9382 15700 10066
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15488 7585 15516 8298
rect 15672 8106 15700 9318
rect 15764 9178 15792 10066
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15856 9586 15884 9998
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 16408 9178 16436 10406
rect 16500 10169 16528 11630
rect 16592 10606 16620 18022
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 17241 16712 17478
rect 16670 17232 16726 17241
rect 16670 17167 16726 17176
rect 17604 16794 17632 17614
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17130 16008 17186 16017
rect 17130 15943 17186 15952
rect 17500 15972 17552 15978
rect 17144 15910 17172 15943
rect 17500 15914 17552 15920
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17144 15638 17172 15846
rect 17132 15632 17184 15638
rect 17132 15574 17184 15580
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16776 15162 16804 15438
rect 17144 15162 17172 15574
rect 17222 15464 17278 15473
rect 17222 15399 17278 15408
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16486 10160 16542 10169
rect 16486 10095 16542 10104
rect 15752 9172 15804 9178
rect 16396 9172 16448 9178
rect 15752 9114 15804 9120
rect 16316 9132 16396 9160
rect 15764 8401 15792 9114
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15750 8392 15806 8401
rect 15750 8327 15806 8336
rect 15672 8078 15792 8106
rect 15474 7576 15530 7585
rect 15474 7511 15530 7520
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15568 6248 15620 6254
rect 15566 6216 15568 6225
rect 15620 6216 15622 6225
rect 15566 6151 15622 6160
rect 15396 5902 15516 5930
rect 15672 5914 15700 7142
rect 15764 6458 15792 8078
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15856 6338 15884 8774
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 16316 8634 16344 9132
rect 16396 9114 16448 9120
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 15934 8392 15990 8401
rect 15934 8327 15936 8336
rect 15988 8327 15990 8336
rect 15936 8298 15988 8304
rect 16408 8090 16436 8910
rect 16500 8430 16528 8910
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16302 7984 16358 7993
rect 16302 7919 16358 7928
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 16316 7342 16344 7919
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16488 7744 16540 7750
rect 16684 7721 16712 14010
rect 16868 14006 16896 14350
rect 17144 14074 17172 14554
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16868 13802 16896 13942
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16868 13462 16896 13738
rect 17236 13530 17264 15399
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 14385 17448 14758
rect 17406 14376 17462 14385
rect 17406 14311 17462 14320
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16868 12986 16896 13398
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 17236 12850 17264 13466
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17328 12986 17356 13262
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16776 10713 16804 11494
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 16762 10704 16818 10713
rect 16762 10639 16818 10648
rect 16960 10470 16988 10950
rect 17052 10674 17080 10950
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 17052 10198 17080 10610
rect 17144 10606 17172 12038
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17144 10266 17172 10542
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17040 10192 17092 10198
rect 17328 10169 17356 12922
rect 17512 10985 17540 15914
rect 17696 12442 17724 18527
rect 17972 14498 18000 20742
rect 22480 20602 22508 23520
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 19062 19272 19118 19281
rect 19062 19207 19118 19216
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18616 18358 18644 18702
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18340 18086 18368 18158
rect 19076 18154 19104 19207
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 24492 18828 24544 18834
rect 24492 18770 24544 18776
rect 19168 18290 19196 18770
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 19996 18426 20024 18566
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18064 14618 18092 14758
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 17972 14470 18092 14498
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17696 11898 17724 12378
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17788 11898 17816 12242
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17880 11762 17908 12174
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 11014 17908 11698
rect 17868 11008 17920 11014
rect 17498 10976 17554 10985
rect 17868 10950 17920 10956
rect 17498 10911 17554 10920
rect 17512 10742 17540 10911
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17040 10134 17092 10140
rect 17314 10160 17370 10169
rect 17314 10095 17370 10104
rect 17130 9344 17186 9353
rect 17130 9279 17186 9288
rect 17144 7954 17172 9279
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17040 7880 17092 7886
rect 17038 7848 17040 7857
rect 17092 7848 17094 7857
rect 17038 7783 17094 7792
rect 16488 7686 16540 7692
rect 16670 7712 16726 7721
rect 16408 7585 16436 7686
rect 16394 7576 16450 7585
rect 16394 7511 16450 7520
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16408 7274 16436 7511
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 16408 6361 16436 7210
rect 16500 6662 16528 7686
rect 16670 7647 16726 7656
rect 17144 7002 17172 7890
rect 17236 7886 17264 8298
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17236 7478 17264 7822
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17328 7313 17356 10095
rect 17420 7750 17448 10406
rect 17880 9654 17908 10950
rect 17972 10010 18000 12582
rect 18064 10130 18092 14470
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17972 9982 18092 10010
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17880 8974 17908 9590
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17512 8090 17540 8774
rect 17880 8634 17908 8910
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17972 8106 18000 9862
rect 18064 9625 18092 9982
rect 18050 9616 18106 9625
rect 18050 9551 18106 9560
rect 18064 9058 18092 9551
rect 18156 9489 18184 17138
rect 18340 16561 18368 18022
rect 18892 17814 18920 18022
rect 18880 17808 18932 17814
rect 18880 17750 18932 17756
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18432 17338 18460 17682
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 18800 16794 18828 16934
rect 18892 16794 18920 17750
rect 19168 17610 19196 18226
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 18970 17504 19026 17513
rect 18970 17439 19026 17448
rect 18984 17202 19012 17439
rect 19168 17202 19196 17546
rect 19260 17338 19288 17614
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18326 16552 18382 16561
rect 18326 16487 18382 16496
rect 18340 14770 18368 16487
rect 19352 16046 19380 18294
rect 20364 17338 20392 18362
rect 21100 18290 21128 18566
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 22112 18086 22140 18770
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22100 18080 22152 18086
rect 20810 18048 20866 18057
rect 22020 18040 22100 18068
rect 20810 17983 20866 17992
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19444 16250 19472 17138
rect 20824 16658 20852 17983
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 22020 17678 22048 18040
rect 22100 18022 22152 18028
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 21376 17338 21404 17614
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 21284 16794 21312 17002
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 19522 16552 19578 16561
rect 19578 16510 19748 16538
rect 19522 16487 19578 16496
rect 19720 16454 19748 16510
rect 19708 16448 19760 16454
rect 19708 16390 19760 16396
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19614 16144 19670 16153
rect 19614 16079 19670 16088
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19352 15706 19380 15982
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19352 15570 19380 15642
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18418 15056 18474 15065
rect 18524 15026 18552 15302
rect 18418 14991 18474 15000
rect 18512 15020 18564 15026
rect 18432 14958 18460 14991
rect 18512 14962 18564 14968
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18510 14920 18566 14929
rect 18510 14855 18512 14864
rect 18564 14855 18566 14864
rect 18512 14826 18564 14832
rect 18340 14742 18552 14770
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18248 13938 18276 14418
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18340 13977 18368 14214
rect 18326 13968 18382 13977
rect 18236 13932 18288 13938
rect 18326 13903 18382 13912
rect 18236 13874 18288 13880
rect 18248 13841 18276 13874
rect 18234 13832 18290 13841
rect 18234 13767 18290 13776
rect 18248 12442 18276 13767
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18418 11928 18474 11937
rect 18418 11863 18474 11872
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18340 9654 18368 10066
rect 18328 9648 18380 9654
rect 18326 9616 18328 9625
rect 18380 9616 18382 9625
rect 18326 9551 18382 9560
rect 18142 9480 18198 9489
rect 18142 9415 18198 9424
rect 18064 9042 18184 9058
rect 18064 9036 18196 9042
rect 18064 9030 18144 9036
rect 18064 8634 18092 9030
rect 18144 8978 18196 8984
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17880 8078 18000 8106
rect 18340 8090 18368 8842
rect 18328 8084 18380 8090
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17512 7546 17540 8026
rect 17880 8022 17908 8078
rect 18328 8026 18380 8032
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17314 7304 17370 7313
rect 17314 7239 17370 7248
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17788 7002 17816 7210
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17880 6934 17908 7958
rect 18432 7546 18460 11863
rect 18524 9081 18552 14742
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18708 13870 18736 14418
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18708 13258 18736 13806
rect 18800 13530 18828 14350
rect 18892 14006 18920 14350
rect 19076 14074 19104 14962
rect 19352 14618 19380 15506
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19352 14346 19380 14554
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 19076 13802 19104 14010
rect 19168 13870 19196 14282
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18800 12986 18828 13466
rect 19248 13320 19300 13326
rect 18878 13288 18934 13297
rect 19248 13262 19300 13268
rect 18878 13223 18934 13232
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18892 12424 18920 13223
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 18800 12396 18920 12424
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18616 11218 18644 11698
rect 18696 11280 18748 11286
rect 18696 11222 18748 11228
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18616 10810 18644 11154
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18708 10742 18736 11222
rect 18696 10736 18748 10742
rect 18696 10678 18748 10684
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18616 9722 18644 10610
rect 18708 10146 18736 10678
rect 18800 10674 18828 12396
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18892 11558 18920 12242
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18892 10577 18920 11494
rect 18878 10568 18934 10577
rect 18878 10503 18934 10512
rect 18708 10118 18828 10146
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18510 9072 18566 9081
rect 18510 9007 18566 9016
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18616 7290 18644 9658
rect 18708 9178 18736 9998
rect 18800 9654 18828 10118
rect 18788 9648 18840 9654
rect 18788 9590 18840 9596
rect 18892 9518 18920 10503
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18788 9376 18840 9382
rect 18786 9344 18788 9353
rect 18840 9344 18842 9353
rect 18786 9279 18842 9288
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18708 8634 18736 9114
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18800 8430 18828 9279
rect 18892 9178 18920 9454
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18984 9058 19012 12650
rect 19260 12186 19288 13262
rect 19168 12158 19288 12186
rect 19168 12102 19196 12158
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 9450 19196 12038
rect 19352 11762 19380 14282
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19444 13326 19472 13738
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19444 12850 19472 13262
rect 19536 13025 19564 13330
rect 19522 13016 19578 13025
rect 19522 12951 19578 12960
rect 19536 12918 19564 12951
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19444 12442 19472 12786
rect 19536 12617 19564 12854
rect 19522 12608 19578 12617
rect 19522 12543 19578 12552
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19260 11014 19288 11290
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19260 10062 19288 10950
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19444 9489 19472 11834
rect 19536 10266 19564 12543
rect 19628 11898 19656 16079
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19720 11778 19748 16390
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20640 15706 20668 16186
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19628 11750 19748 11778
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19536 9518 19564 10202
rect 19524 9512 19576 9518
rect 19430 9480 19486 9489
rect 19156 9444 19208 9450
rect 19524 9454 19576 9460
rect 19430 9415 19486 9424
rect 19156 9386 19208 9392
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 9110 19104 9318
rect 18892 9030 19012 9058
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 18892 8974 18920 9030
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18892 8430 18920 8910
rect 19444 8498 19472 9415
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 18788 8424 18840 8430
rect 18880 8424 18932 8430
rect 18788 8366 18840 8372
rect 18878 8392 18880 8401
rect 18932 8392 18934 8401
rect 19444 8378 19472 8434
rect 18878 8327 18934 8336
rect 19260 8350 19472 8378
rect 18616 7262 18828 7290
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16394 6352 16450 6361
rect 15856 6310 16344 6338
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15120 5868 15240 5896
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 15120 5098 15148 5868
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15212 5370 15240 5714
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 15304 4826 15332 5510
rect 15396 5370 15424 5646
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 14556 4014 14608 4020
rect 14646 4040 14702 4049
rect 14568 3534 14596 4014
rect 14646 3975 14702 3984
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 13280 2990 13308 3130
rect 14476 2990 14504 3130
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 12360 2514 12480 2530
rect 12360 2508 12492 2514
rect 12360 2502 12440 2508
rect 12440 2450 12492 2456
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12084 480 12112 2382
rect 13464 480 13492 2858
rect 13726 2816 13782 2825
rect 13726 2751 13782 2760
rect 13740 2582 13768 2751
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 14936 480 14964 2858
rect 15304 2514 15332 4422
rect 15488 3913 15516 5902
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15672 5370 15700 5850
rect 15764 5778 15792 6054
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15856 5234 15884 6122
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 16316 5273 16344 6310
rect 16394 6287 16450 6296
rect 16302 5264 16358 5273
rect 15844 5228 15896 5234
rect 16302 5199 16358 5208
rect 15844 5170 15896 5176
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15764 4282 15792 4626
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15474 3904 15530 3913
rect 15474 3839 15530 3848
rect 15856 3738 15884 4762
rect 16500 4729 16528 6394
rect 16684 6322 16712 6598
rect 18524 6322 18552 6598
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 17960 6112 18012 6118
rect 17880 6060 17960 6066
rect 17880 6054 18012 6060
rect 17880 6038 18000 6054
rect 17880 5370 17908 6038
rect 17972 5846 18000 6038
rect 18524 5914 18552 6258
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 18050 5264 18106 5273
rect 18616 5234 18644 6258
rect 18708 6254 18736 7142
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18050 5199 18106 5208
rect 18604 5228 18656 5234
rect 16486 4720 16542 4729
rect 16486 4655 16542 4664
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 16316 4214 16344 4558
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 16316 3602 16344 4150
rect 17958 4040 18014 4049
rect 17958 3975 18014 3984
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 16316 3194 16344 3538
rect 17788 3398 17816 3538
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16408 3126 16436 3334
rect 17788 3194 17816 3334
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 16396 3120 16448 3126
rect 16396 3062 16448 3068
rect 17972 2990 18000 3975
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 16302 2816 16358 2825
rect 16302 2751 16358 2760
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 16316 480 16344 2751
rect 18064 2650 18092 5199
rect 18604 5170 18656 5176
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18524 3126 18552 3470
rect 18800 3194 18828 7262
rect 18892 6769 18920 8327
rect 19260 8090 19288 8350
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19154 7848 19210 7857
rect 19154 7783 19210 7792
rect 19168 7002 19196 7783
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 18878 6760 18934 6769
rect 18878 6695 18934 6704
rect 19168 6458 19196 6938
rect 19246 6896 19302 6905
rect 19246 6831 19248 6840
rect 19300 6831 19302 6840
rect 19248 6802 19300 6808
rect 19260 6458 19288 6802
rect 19444 6798 19472 7346
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19444 6254 19472 6734
rect 19536 6361 19564 9318
rect 19628 8430 19656 11750
rect 19706 11656 19762 11665
rect 19706 11591 19708 11600
rect 19760 11591 19762 11600
rect 19708 11562 19760 11568
rect 19904 10441 19932 15098
rect 20732 15026 20760 15914
rect 21284 15892 21312 16594
rect 21376 16250 21404 17070
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21364 15904 21416 15910
rect 21284 15864 21364 15892
rect 21364 15846 21416 15852
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21192 15162 21220 15438
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20732 14657 20760 14758
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20718 14648 20774 14657
rect 20956 14640 21252 14660
rect 20718 14583 20774 14592
rect 21284 14074 21312 14962
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21376 13954 21404 15846
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 21284 13926 21404 13954
rect 20732 13705 20760 13874
rect 21180 13864 21232 13870
rect 21178 13832 21180 13841
rect 21232 13832 21234 13841
rect 21178 13767 21234 13776
rect 20718 13696 20774 13705
rect 20718 13631 20774 13640
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 21284 13410 21312 13926
rect 21362 13832 21418 13841
rect 21468 13818 21496 17478
rect 21560 17270 21588 17614
rect 22204 17610 22232 18566
rect 24504 18290 24532 18770
rect 24584 18624 24636 18630
rect 24964 18601 24992 23559
rect 27526 23080 27582 23089
rect 27526 23015 27582 23024
rect 25042 22400 25098 22409
rect 25042 22335 25098 22344
rect 24584 18566 24636 18572
rect 24950 18592 25006 18601
rect 24492 18284 24544 18290
rect 24492 18226 24544 18232
rect 24596 18086 24624 18566
rect 25056 18578 25084 22335
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25686 21584 25742 21593
rect 25686 21519 25742 21528
rect 25502 21312 25558 21321
rect 25502 21247 25558 21256
rect 25410 18864 25466 18873
rect 25410 18799 25466 18808
rect 25056 18550 25268 18578
rect 24950 18527 25006 18536
rect 24858 18320 24914 18329
rect 24858 18255 24914 18264
rect 25044 18284 25096 18290
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22664 17338 22692 17682
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 21548 17264 21600 17270
rect 21548 17206 21600 17212
rect 23480 16720 23532 16726
rect 23480 16662 23532 16668
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21548 16516 21600 16522
rect 21548 16458 21600 16464
rect 21560 16114 21588 16458
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 21560 15706 21588 16050
rect 21652 15706 21680 16526
rect 21836 15978 21864 16526
rect 23492 16250 23520 16662
rect 23584 16658 23612 17546
rect 24228 17338 24256 17818
rect 24596 17610 24624 18022
rect 24872 17626 24900 18255
rect 25044 18226 25096 18232
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 24584 17604 24636 17610
rect 24584 17546 24636 17552
rect 24780 17598 24900 17626
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24780 17105 24808 17598
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24766 17096 24822 17105
rect 24766 17031 24822 17040
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21744 13841 21772 14894
rect 21836 14618 21864 15914
rect 21916 15904 21968 15910
rect 22836 15904 22888 15910
rect 21916 15846 21968 15852
rect 22742 15872 22798 15881
rect 21928 15162 21956 15846
rect 22836 15846 22888 15852
rect 22742 15807 22798 15816
rect 22756 15586 22784 15807
rect 22848 15706 22876 15846
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 22664 15570 22784 15586
rect 22652 15564 22784 15570
rect 22704 15558 22784 15564
rect 22652 15506 22704 15512
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 22296 15026 22324 15438
rect 22756 15162 22784 15558
rect 23584 15366 23612 16594
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24688 16114 24716 16390
rect 24872 16130 24900 17478
rect 24964 17270 24992 17682
rect 24952 17264 25004 17270
rect 24952 17206 25004 17212
rect 24964 16726 24992 17206
rect 24952 16720 25004 16726
rect 24952 16662 25004 16668
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24780 16102 24900 16130
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 22744 15156 22796 15162
rect 22664 15116 22744 15144
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21836 14113 21864 14418
rect 21822 14104 21878 14113
rect 21822 14039 21824 14048
rect 21876 14039 21878 14048
rect 21824 14010 21876 14016
rect 21836 13979 21864 14010
rect 21730 13832 21786 13841
rect 21468 13790 21680 13818
rect 21362 13767 21418 13776
rect 21376 13530 21404 13767
rect 21548 13728 21600 13734
rect 21548 13670 21600 13676
rect 21652 13682 21680 13790
rect 21730 13767 21786 13776
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21284 13382 21404 13410
rect 21560 13394 21588 13670
rect 21652 13654 21772 13682
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 21376 12424 21404 13382
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21560 12918 21588 13330
rect 21548 12912 21600 12918
rect 21548 12854 21600 12860
rect 21376 12396 21496 12424
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20824 11286 20852 11494
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 19890 10432 19946 10441
rect 19890 10367 19946 10376
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19720 8974 19748 9590
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19720 8634 19748 8910
rect 19812 8809 19840 8978
rect 19798 8800 19854 8809
rect 19798 8735 19854 8744
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19628 8090 19656 8366
rect 19720 8090 19748 8570
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 19522 6352 19578 6361
rect 19628 6322 19656 6938
rect 19522 6287 19578 6296
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19444 5914 19472 6190
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 18892 5370 18920 5646
rect 19076 5409 19104 5646
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19062 5400 19118 5409
rect 18880 5364 18932 5370
rect 19062 5335 19118 5344
rect 18880 5306 18932 5312
rect 18892 4826 18920 5306
rect 19076 5302 19104 5335
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 19076 4282 19104 5102
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 18880 3936 18932 3942
rect 18878 3904 18880 3913
rect 18932 3904 18934 3913
rect 18878 3839 18934 3848
rect 18984 3194 19012 3946
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18512 3120 18564 3126
rect 18512 3062 18564 3068
rect 18602 3088 18658 3097
rect 18602 3023 18658 3032
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18616 2582 18644 3023
rect 18800 2922 18828 3130
rect 19076 3058 19104 3538
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 19076 2650 19104 2994
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 19168 2530 19196 5510
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19260 4826 19288 5034
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19444 4758 19472 5850
rect 19904 4826 19932 10367
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20548 8634 20576 9590
rect 21468 9586 21496 12396
rect 21560 12306 21588 12854
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21560 11830 21588 12242
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 21560 11218 21588 11766
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21652 9722 21680 9998
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 21376 8945 21404 9522
rect 21362 8936 21418 8945
rect 21362 8871 21418 8880
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20548 7002 20576 8570
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 21376 7954 21404 8871
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20824 5234 20852 6054
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 21376 5166 21404 5714
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 21376 4826 21404 5102
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 19432 4752 19484 4758
rect 19246 4720 19302 4729
rect 19432 4694 19484 4700
rect 19246 4655 19302 4664
rect 19260 4622 19288 4655
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19260 4146 19288 4558
rect 19444 4146 19472 4694
rect 19904 4282 19932 4762
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19444 3738 19472 4082
rect 19904 4049 19932 4218
rect 19890 4040 19946 4049
rect 19890 3975 19946 3984
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19628 3641 19656 3878
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 19614 3632 19670 3641
rect 19614 3567 19670 3576
rect 21560 3194 21588 8774
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 19432 2984 19484 2990
rect 19430 2952 19432 2961
rect 19484 2952 19486 2961
rect 19430 2887 19486 2896
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 19168 2514 19380 2530
rect 19168 2508 19392 2514
rect 19168 2502 19340 2508
rect 19340 2450 19392 2456
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 17788 480 17816 2382
rect 19168 480 19196 2382
rect 20640 480 20668 2858
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 21744 2650 21772 13654
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21836 12986 21864 13330
rect 21928 13297 21956 14826
rect 22296 14414 22324 14962
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 22020 13938 22048 14282
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21914 13288 21970 13297
rect 21914 13223 21970 13232
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21836 10266 21864 12922
rect 22020 12889 22048 13874
rect 22006 12880 22062 12889
rect 22006 12815 22062 12824
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 21928 11898 21956 12242
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22192 11280 22244 11286
rect 22020 11240 22192 11268
rect 22020 10810 22048 11240
rect 22192 11222 22244 11228
rect 22296 10810 22324 11290
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21836 8906 21864 10202
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21928 9722 21956 10066
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21928 9450 21956 9658
rect 21916 9444 21968 9450
rect 21916 9386 21968 9392
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21836 8634 21864 8842
rect 22020 8634 22048 8910
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21836 7546 21864 8366
rect 21928 8022 21956 8434
rect 22020 8090 22048 8570
rect 22112 8498 22140 9386
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22388 8090 22416 8230
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 22376 8084 22428 8090
rect 22376 8026 22428 8032
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22296 6934 22324 7346
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22480 7002 22508 7142
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22284 6928 22336 6934
rect 22664 6905 22692 15116
rect 22744 15098 22796 15104
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23124 14414 23152 14758
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23124 13530 23152 14350
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23400 13682 23428 13806
rect 23400 13654 23520 13682
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23492 12442 23520 13654
rect 23938 12880 23994 12889
rect 23938 12815 23940 12824
rect 23992 12815 23994 12824
rect 23940 12786 23992 12792
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23032 11830 23060 12038
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 23032 11286 23060 11766
rect 23294 11656 23350 11665
rect 23294 11591 23350 11600
rect 23308 11354 23336 11591
rect 23848 11552 23900 11558
rect 23848 11494 23900 11500
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23020 11280 23072 11286
rect 23020 11222 23072 11228
rect 23308 11098 23336 11290
rect 23308 11070 23520 11098
rect 23492 10810 23520 11070
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23860 10674 23888 11494
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23204 9716 23256 9722
rect 23204 9658 23256 9664
rect 23216 8401 23244 9658
rect 23492 9058 23520 9862
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23400 9042 23520 9058
rect 23388 9036 23520 9042
rect 23440 9030 23520 9036
rect 23388 8978 23440 8984
rect 23294 8800 23350 8809
rect 23294 8735 23350 8744
rect 23202 8392 23258 8401
rect 23202 8327 23258 8336
rect 23112 7948 23164 7954
rect 23112 7890 23164 7896
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22848 7478 22876 7822
rect 22836 7472 22888 7478
rect 22836 7414 22888 7420
rect 22848 6934 22876 7414
rect 22940 7410 22968 7822
rect 23124 7721 23152 7890
rect 23110 7712 23166 7721
rect 23110 7647 23166 7656
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 23124 7206 23152 7647
rect 23112 7200 23164 7206
rect 23110 7168 23112 7177
rect 23164 7168 23166 7177
rect 23110 7103 23166 7112
rect 22836 6928 22888 6934
rect 22284 6870 22336 6876
rect 22650 6896 22706 6905
rect 22836 6870 22888 6876
rect 23216 6866 23244 8327
rect 23308 7002 23336 8735
rect 23388 8628 23440 8634
rect 23492 8616 23520 9030
rect 23440 8588 23520 8616
rect 23388 8570 23440 8576
rect 23584 8004 23612 9386
rect 23400 7976 23612 8004
rect 23400 7886 23428 7976
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23400 7154 23428 7210
rect 23400 7126 23520 7154
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 22650 6831 22706 6840
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23216 6322 23244 6802
rect 23308 6458 23336 6938
rect 23492 6458 23520 7126
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23584 6390 23612 6734
rect 23572 6384 23624 6390
rect 23478 6352 23534 6361
rect 23204 6316 23256 6322
rect 23572 6326 23624 6332
rect 23478 6287 23534 6296
rect 23204 6258 23256 6264
rect 23216 6225 23244 6258
rect 23492 6254 23520 6287
rect 23480 6248 23532 6254
rect 23202 6216 23258 6225
rect 23480 6190 23532 6196
rect 23202 6151 23258 6160
rect 22744 5840 22796 5846
rect 22744 5782 22796 5788
rect 22756 5409 22784 5782
rect 23388 5772 23440 5778
rect 23388 5714 23440 5720
rect 22742 5400 22798 5409
rect 23400 5370 23428 5714
rect 22742 5335 22744 5344
rect 22796 5335 22798 5344
rect 23388 5364 23440 5370
rect 22744 5306 22796 5312
rect 23388 5306 23440 5312
rect 23676 2990 23704 10406
rect 23860 10266 23888 10610
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 23768 8838 23796 9454
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23860 8430 23888 8910
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23952 7585 23980 8026
rect 23938 7576 23994 7585
rect 23938 7511 23994 7520
rect 23952 7342 23980 7511
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 24044 2650 24072 15846
rect 24228 14074 24256 16050
rect 24780 16046 24808 16102
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24492 15904 24544 15910
rect 24492 15846 24544 15852
rect 24504 15706 24532 15846
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24676 15632 24728 15638
rect 24676 15574 24728 15580
rect 24308 15360 24360 15366
rect 24308 15302 24360 15308
rect 24320 14278 24348 15302
rect 24688 15162 24716 15574
rect 24780 15570 24808 15982
rect 24964 15688 24992 16118
rect 24872 15660 24992 15688
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 24320 13870 24348 14214
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24214 13696 24270 13705
rect 24214 13631 24270 13640
rect 24228 13025 24256 13631
rect 24214 13016 24270 13025
rect 24214 12951 24270 12960
rect 24124 12164 24176 12170
rect 24124 12106 24176 12112
rect 24136 11694 24164 12106
rect 24124 11688 24176 11694
rect 24124 11630 24176 11636
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 7410 24164 7686
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24136 6390 24164 7346
rect 24228 6866 24256 12951
rect 24320 12918 24348 13806
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24308 12912 24360 12918
rect 24308 12854 24360 12860
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 24320 11762 24348 12582
rect 24412 12306 24440 12786
rect 24688 12782 24716 13126
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24766 12336 24822 12345
rect 24400 12300 24452 12306
rect 24766 12271 24768 12280
rect 24400 12242 24452 12248
rect 24820 12271 24822 12280
rect 24768 12242 24820 12248
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 24320 11354 24348 11698
rect 24412 11354 24440 12242
rect 24780 11898 24808 12242
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24490 11792 24546 11801
rect 24490 11727 24546 11736
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24504 8634 24532 11727
rect 24872 11286 24900 15660
rect 24950 15464 25006 15473
rect 24950 15399 25006 15408
rect 24964 12102 24992 15399
rect 25056 15366 25084 18226
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 25148 17134 25176 18022
rect 25240 17377 25268 18550
rect 25424 18057 25452 18799
rect 25410 18048 25466 18057
rect 25410 17983 25466 17992
rect 25320 17672 25372 17678
rect 25320 17614 25372 17620
rect 25226 17368 25282 17377
rect 25332 17338 25360 17614
rect 25226 17303 25282 17312
rect 25320 17332 25372 17338
rect 25320 17274 25372 17280
rect 25516 17218 25544 21247
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 18154 25636 18566
rect 25596 18148 25648 18154
rect 25596 18090 25648 18096
rect 25594 18048 25650 18057
rect 25594 17983 25650 17992
rect 25332 17190 25544 17218
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 25226 17096 25282 17105
rect 25226 17031 25282 17040
rect 25136 15904 25188 15910
rect 25136 15846 25188 15852
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 25042 13560 25098 13569
rect 25042 13495 25098 13504
rect 25056 12442 25084 13495
rect 25148 12481 25176 15846
rect 25240 13920 25268 17031
rect 25332 14940 25360 17190
rect 25502 17096 25558 17105
rect 25502 17031 25558 17040
rect 25412 16720 25464 16726
rect 25412 16662 25464 16668
rect 25424 15502 25452 16662
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25424 15094 25452 15438
rect 25412 15088 25464 15094
rect 25412 15030 25464 15036
rect 25332 14912 25452 14940
rect 25240 13892 25360 13920
rect 25226 13832 25282 13841
rect 25226 13767 25282 13776
rect 25240 13530 25268 13767
rect 25228 13524 25280 13530
rect 25228 13466 25280 13472
rect 25240 12918 25268 13466
rect 25332 13462 25360 13892
rect 25320 13456 25372 13462
rect 25320 13398 25372 13404
rect 25320 13320 25372 13326
rect 25318 13288 25320 13297
rect 25372 13288 25374 13297
rect 25318 13223 25374 13232
rect 25332 12986 25360 13223
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25228 12912 25280 12918
rect 25228 12854 25280 12860
rect 25134 12472 25190 12481
rect 25044 12436 25096 12442
rect 25134 12407 25190 12416
rect 25044 12378 25096 12384
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 25056 11898 25084 12378
rect 25240 12345 25268 12854
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 25226 12336 25282 12345
rect 25226 12271 25282 12280
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24860 11280 24912 11286
rect 24860 11222 24912 11228
rect 24964 11150 24992 11698
rect 25044 11280 25096 11286
rect 25044 11222 25096 11228
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24872 10690 24900 11018
rect 24964 10810 24992 11086
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 24780 10662 24900 10690
rect 24780 10606 24808 10662
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24952 10192 25004 10198
rect 25056 10169 25084 11222
rect 24952 10134 25004 10140
rect 25042 10160 25098 10169
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24872 9654 24900 9998
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24872 9178 24900 9590
rect 24964 9586 24992 10134
rect 25042 10095 25098 10104
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 25056 9382 25084 9998
rect 25044 9376 25096 9382
rect 24950 9344 25006 9353
rect 25044 9318 25096 9324
rect 24950 9279 25006 9288
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24504 8362 24532 8570
rect 24492 8356 24544 8362
rect 24492 8298 24544 8304
rect 24688 7206 24716 8774
rect 24308 7200 24360 7206
rect 24308 7142 24360 7148
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24136 5914 24164 6326
rect 24228 6186 24256 6802
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24320 5273 24348 7142
rect 24688 5778 24716 7142
rect 24964 6338 24992 9279
rect 25056 9110 25084 9318
rect 25044 9104 25096 9110
rect 25044 9046 25096 9052
rect 25148 8090 25176 12038
rect 25332 11506 25360 12786
rect 25424 11801 25452 14912
rect 25516 12850 25544 17031
rect 25608 16182 25636 17983
rect 25700 17513 25728 21519
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 25870 20496 25926 20505
rect 25870 20431 25926 20440
rect 25778 20088 25834 20097
rect 25778 20023 25834 20032
rect 25792 18737 25820 20023
rect 25778 18728 25834 18737
rect 25778 18663 25834 18672
rect 25884 17762 25912 20431
rect 25962 20360 26018 20369
rect 25962 20295 26018 20304
rect 25976 20262 26004 20295
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 26240 18080 26292 18086
rect 27540 18057 27568 23015
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 26240 18022 26292 18028
rect 26974 18048 27030 18057
rect 25792 17734 25912 17762
rect 25686 17504 25742 17513
rect 25686 17439 25742 17448
rect 25792 16266 25820 17734
rect 26148 17672 26200 17678
rect 26252 17660 26280 18022
rect 26974 17983 27030 17992
rect 27526 18048 27582 18057
rect 27526 17983 27582 17992
rect 26200 17632 26280 17660
rect 26792 17672 26844 17678
rect 26148 17614 26200 17620
rect 26792 17614 26844 17620
rect 26332 17604 26384 17610
rect 26332 17546 26384 17552
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 26344 17202 26372 17546
rect 26804 17270 26832 17614
rect 26792 17264 26844 17270
rect 26790 17232 26792 17241
rect 26844 17232 26846 17241
rect 26332 17196 26384 17202
rect 26790 17167 26846 17176
rect 26332 17138 26384 17144
rect 26240 17060 26292 17066
rect 26240 17002 26292 17008
rect 26252 16522 26280 17002
rect 26240 16516 26292 16522
rect 26240 16458 26292 16464
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 25700 16238 25820 16266
rect 25596 16176 25648 16182
rect 25596 16118 25648 16124
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 25608 15706 25636 15846
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25608 15162 25636 15642
rect 25596 15156 25648 15162
rect 25596 15098 25648 15104
rect 25700 15042 25728 16238
rect 25778 16144 25834 16153
rect 26344 16114 26372 17138
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 25778 16079 25834 16088
rect 26332 16108 26384 16114
rect 25792 15065 25820 16079
rect 26332 16050 26384 16056
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 25884 15162 25912 15914
rect 26436 15609 26464 16934
rect 26422 15600 26478 15609
rect 26422 15535 26478 15544
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 25872 15156 25924 15162
rect 25872 15098 25924 15104
rect 25608 15014 25728 15042
rect 25778 15056 25834 15065
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 25504 12708 25556 12714
rect 25504 12650 25556 12656
rect 25516 12442 25544 12650
rect 25608 12442 25636 15014
rect 26344 15026 26372 15302
rect 25778 14991 25834 15000
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25504 12436 25556 12442
rect 25504 12378 25556 12384
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25700 12322 25728 14758
rect 25778 14648 25834 14657
rect 25778 14583 25834 14592
rect 25792 13433 25820 14583
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 25872 13728 25924 13734
rect 25872 13670 25924 13676
rect 25778 13424 25834 13433
rect 25778 13359 25834 13368
rect 25780 13252 25832 13258
rect 25780 13194 25832 13200
rect 25516 12294 25728 12322
rect 25410 11792 25466 11801
rect 25410 11727 25466 11736
rect 25240 11478 25360 11506
rect 25240 10033 25268 11478
rect 25516 11370 25544 12294
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 25792 12186 25820 13194
rect 25884 13190 25912 13670
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 25884 12714 25912 13126
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 25872 12708 25924 12714
rect 25872 12650 25924 12656
rect 26148 12708 26200 12714
rect 26148 12650 26200 12656
rect 26160 12594 26188 12650
rect 26160 12566 26280 12594
rect 26252 12442 26280 12566
rect 26240 12436 26292 12442
rect 26240 12378 26292 12384
rect 25608 11937 25636 12174
rect 25688 12164 25740 12170
rect 25792 12158 25912 12186
rect 25688 12106 25740 12112
rect 25594 11928 25650 11937
rect 25594 11863 25650 11872
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25424 11342 25544 11370
rect 25332 10810 25360 11290
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25318 10160 25374 10169
rect 25318 10095 25374 10104
rect 25226 10024 25282 10033
rect 25226 9959 25282 9968
rect 25226 9616 25282 9625
rect 25226 9551 25282 9560
rect 25240 9178 25268 9551
rect 25332 9178 25360 10095
rect 25424 9722 25452 11342
rect 25504 11280 25556 11286
rect 25504 11222 25556 11228
rect 25516 10266 25544 11222
rect 25608 10985 25636 11494
rect 25594 10976 25650 10985
rect 25594 10911 25650 10920
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25608 10130 25636 10911
rect 25596 10124 25648 10130
rect 25596 10066 25648 10072
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25240 8634 25268 9114
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25332 8498 25360 9114
rect 25424 8634 25452 9522
rect 25504 9444 25556 9450
rect 25504 9386 25556 9392
rect 25516 8974 25544 9386
rect 25504 8968 25556 8974
rect 25504 8910 25556 8916
rect 25700 8809 25728 12106
rect 25884 12102 25912 12158
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25884 11762 25912 12038
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 25872 11756 25924 11762
rect 25872 11698 25924 11704
rect 25964 11688 26016 11694
rect 25884 11636 25964 11642
rect 25884 11630 26016 11636
rect 25884 11614 26004 11630
rect 25780 11552 25832 11558
rect 25780 11494 25832 11500
rect 25792 11354 25820 11494
rect 25780 11348 25832 11354
rect 25780 11290 25832 11296
rect 25884 11218 25912 11614
rect 25872 11212 25924 11218
rect 25872 11154 25924 11160
rect 25884 10810 25912 11154
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 25872 10804 25924 10810
rect 26436 10792 26464 15535
rect 26514 14920 26570 14929
rect 26514 14855 26570 14864
rect 26528 13870 26556 14855
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26620 14278 26648 14758
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 26620 12889 26648 14214
rect 26884 14000 26936 14006
rect 26884 13942 26936 13948
rect 26606 12880 26662 12889
rect 26606 12815 26662 12824
rect 26620 12170 26648 12815
rect 26896 12322 26924 13942
rect 26804 12294 26924 12322
rect 26608 12164 26660 12170
rect 26608 12106 26660 12112
rect 26516 11824 26568 11830
rect 26516 11766 26568 11772
rect 25872 10746 25924 10752
rect 26344 10764 26464 10792
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26344 9518 26372 10764
rect 26422 10704 26478 10713
rect 26422 10639 26478 10648
rect 26436 10606 26464 10639
rect 26424 10600 26476 10606
rect 26424 10542 26476 10548
rect 26528 9704 26556 11766
rect 26606 11656 26662 11665
rect 26606 11591 26662 11600
rect 26620 10742 26648 11591
rect 26698 11112 26754 11121
rect 26698 11047 26754 11056
rect 26608 10736 26660 10742
rect 26608 10678 26660 10684
rect 26606 10432 26662 10441
rect 26606 10367 26662 10376
rect 26436 9676 26556 9704
rect 26332 9512 26384 9518
rect 26332 9454 26384 9460
rect 25872 8832 25924 8838
rect 25686 8800 25742 8809
rect 25872 8774 25924 8780
rect 25686 8735 25742 8744
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25884 8514 25912 8774
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 25884 8498 26004 8514
rect 25320 8492 25372 8498
rect 25884 8492 26016 8498
rect 25884 8486 25964 8492
rect 25320 8434 25372 8440
rect 25964 8434 26016 8440
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 25872 8424 25924 8430
rect 25778 8392 25834 8401
rect 25872 8366 25924 8372
rect 25778 8327 25834 8336
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 25044 7948 25096 7954
rect 25044 7890 25096 7896
rect 25056 7546 25084 7890
rect 25504 7744 25556 7750
rect 25504 7686 25556 7692
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 25516 7449 25544 7686
rect 25502 7440 25558 7449
rect 25502 7375 25558 7384
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25240 6662 25268 7142
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25240 6390 25268 6598
rect 24780 6310 24992 6338
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 24780 6254 24808 6310
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24964 5817 24992 6310
rect 25686 6216 25742 6225
rect 25686 6151 25742 6160
rect 24950 5808 25006 5817
rect 24676 5772 24728 5778
rect 24950 5743 25006 5752
rect 24676 5714 24728 5720
rect 24306 5264 24362 5273
rect 24306 5199 24362 5208
rect 24320 4593 24348 5199
rect 24306 4584 24362 4593
rect 24306 4519 24362 4528
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 22020 480 22048 2382
rect 23492 480 23520 2382
rect 24872 480 24900 2858
rect 25700 2514 25728 6151
rect 25792 4593 25820 8327
rect 25884 8090 25912 8366
rect 26160 8242 26188 8434
rect 26160 8214 26372 8242
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 26344 8022 26372 8214
rect 26332 8016 26384 8022
rect 26332 7958 26384 7964
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 26344 7478 26372 7958
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 26436 6254 26464 9676
rect 26620 9654 26648 10367
rect 26712 10266 26740 11047
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26698 9888 26754 9897
rect 26698 9823 26754 9832
rect 26608 9648 26660 9654
rect 26608 9590 26660 9596
rect 26712 9178 26740 9823
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26514 9072 26570 9081
rect 26514 9007 26516 9016
rect 26568 9007 26570 9016
rect 26516 8978 26568 8984
rect 26528 8634 26556 8978
rect 26698 8664 26754 8673
rect 26516 8628 26568 8634
rect 26698 8599 26754 8608
rect 26516 8570 26568 8576
rect 26712 8090 26740 8599
rect 26804 8401 26832 12294
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26896 11286 26924 12174
rect 26988 11354 27016 17983
rect 27160 17740 27212 17746
rect 27160 17682 27212 17688
rect 27172 16998 27200 17682
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 27172 16794 27200 16934
rect 27160 16788 27212 16794
rect 27160 16730 27212 16736
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27172 16114 27200 16390
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27068 15632 27120 15638
rect 27068 15574 27120 15580
rect 27080 14822 27108 15574
rect 27172 15502 27200 16050
rect 27252 15564 27304 15570
rect 27252 15506 27304 15512
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 27068 14816 27120 14822
rect 27068 14758 27120 14764
rect 26976 11348 27028 11354
rect 26976 11290 27028 11296
rect 26884 11280 26936 11286
rect 26884 11222 26936 11228
rect 26896 10810 26924 11222
rect 26988 10810 27016 11290
rect 26884 10804 26936 10810
rect 26884 10746 26936 10752
rect 26976 10804 27028 10810
rect 26976 10746 27028 10752
rect 27080 9489 27108 14758
rect 27172 14618 27200 15438
rect 27264 14822 27292 15506
rect 27252 14816 27304 14822
rect 27252 14758 27304 14764
rect 27160 14612 27212 14618
rect 27160 14554 27212 14560
rect 27264 14113 27292 14758
rect 27250 14104 27306 14113
rect 27250 14039 27306 14048
rect 27264 13841 27292 14039
rect 27250 13832 27306 13841
rect 27250 13767 27306 13776
rect 27160 12640 27212 12646
rect 27160 12582 27212 12588
rect 27172 11218 27200 12582
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 27344 10124 27396 10130
rect 27344 10066 27396 10072
rect 27356 9722 27384 10066
rect 27344 9716 27396 9722
rect 27344 9658 27396 9664
rect 27066 9480 27122 9489
rect 27066 9415 27122 9424
rect 26790 8392 26846 8401
rect 26790 8327 26846 8336
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 26528 7857 26556 7890
rect 26514 7848 26570 7857
rect 26514 7783 26570 7792
rect 26528 7546 26556 7783
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 26514 7168 26570 7177
rect 26514 7103 26570 7112
rect 26528 6866 26556 7103
rect 26698 6896 26754 6905
rect 26516 6860 26568 6866
rect 26698 6831 26754 6840
rect 26516 6802 26568 6808
rect 26712 6730 26740 6831
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26608 6384 26660 6390
rect 26606 6352 26608 6361
rect 26660 6352 26662 6361
rect 26606 6287 26662 6296
rect 26424 6248 26476 6254
rect 26424 6190 26476 6196
rect 27080 5778 27108 9415
rect 27158 9344 27214 9353
rect 27158 9279 27214 9288
rect 27172 8634 27200 9279
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 27434 8120 27490 8129
rect 27434 8055 27490 8064
rect 27618 8120 27674 8129
rect 27618 8055 27674 8064
rect 27448 7342 27476 8055
rect 27632 7546 27660 8055
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27356 6458 27384 6802
rect 27344 6452 27396 6458
rect 27344 6394 27396 6400
rect 27434 5808 27490 5817
rect 27068 5772 27120 5778
rect 27434 5743 27490 5752
rect 27068 5714 27120 5720
rect 26698 5672 26754 5681
rect 26698 5607 26700 5616
rect 26752 5607 26754 5616
rect 26700 5578 26752 5584
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 27080 5370 27108 5714
rect 27068 5364 27120 5370
rect 27068 5306 27120 5312
rect 26514 5264 26570 5273
rect 26514 5199 26570 5208
rect 26424 5160 26476 5166
rect 26422 5128 26424 5137
rect 26476 5128 26478 5137
rect 26422 5063 26478 5072
rect 26528 4690 26556 5199
rect 26606 5128 26662 5137
rect 26606 5063 26662 5072
rect 26620 5030 26648 5063
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26516 4684 26568 4690
rect 26516 4626 26568 4632
rect 27344 4684 27396 4690
rect 27344 4626 27396 4632
rect 25778 4584 25834 4593
rect 25778 4519 25834 4528
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 26424 4072 26476 4078
rect 26424 4014 26476 4020
rect 26436 3505 26464 4014
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26514 3632 26570 3641
rect 26514 3567 26516 3576
rect 26568 3567 26570 3576
rect 26516 3538 26568 3544
rect 26422 3496 26478 3505
rect 26422 3431 26478 3440
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 26528 3194 26556 3538
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26238 3088 26294 3097
rect 26238 3023 26294 3032
rect 26252 2802 26280 3023
rect 26332 2984 26384 2990
rect 26330 2952 26332 2961
rect 26384 2952 26386 2961
rect 26330 2887 26386 2896
rect 26516 2848 26568 2854
rect 26252 2774 26372 2802
rect 26620 2825 26648 3878
rect 26712 3369 26740 4422
rect 27356 4282 27384 4626
rect 27344 4276 27396 4282
rect 27344 4218 27396 4224
rect 26792 3392 26844 3398
rect 26698 3360 26754 3369
rect 26792 3334 26844 3340
rect 26698 3295 26754 3304
rect 26516 2790 26568 2796
rect 26606 2816 26662 2825
rect 25688 2508 25740 2514
rect 25688 2450 25740 2456
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25884 921 25912 2246
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 25870 912 25926 921
rect 25870 847 25926 856
rect 26344 480 26372 2774
rect 2778 368 2834 377
rect 2778 303 2834 312
rect 3514 0 3570 480
rect 4894 0 4950 480
rect 6366 0 6422 480
rect 7746 0 7802 480
rect 9218 0 9274 480
rect 10598 0 10654 480
rect 12070 0 12126 480
rect 13450 0 13506 480
rect 14922 0 14978 480
rect 16302 0 16358 480
rect 17774 0 17830 480
rect 19154 0 19210 480
rect 20626 0 20682 480
rect 22006 0 22062 480
rect 23478 0 23534 480
rect 24858 0 24914 480
rect 26330 0 26386 480
rect 26528 377 26556 2790
rect 26606 2751 26662 2760
rect 26804 1465 26832 3334
rect 27448 2990 27476 5743
rect 27528 4072 27580 4078
rect 27526 4040 27528 4049
rect 27580 4040 27582 4049
rect 27526 3975 27582 3984
rect 27712 3936 27764 3942
rect 27710 3904 27712 3913
rect 27764 3904 27766 3913
rect 27710 3839 27766 3848
rect 27436 2984 27488 2990
rect 27436 2926 27488 2932
rect 27620 2848 27672 2854
rect 27816 2802 27844 20198
rect 29182 17640 29238 17649
rect 29182 17575 29238 17584
rect 29196 17066 29224 17575
rect 29184 17060 29236 17066
rect 29184 17002 29236 17008
rect 27620 2790 27672 2796
rect 27632 2145 27660 2790
rect 27724 2774 27844 2802
rect 27618 2136 27674 2145
rect 27618 2071 27674 2080
rect 26790 1456 26846 1465
rect 26790 1391 26846 1400
rect 27724 480 27752 2774
rect 29184 2304 29236 2310
rect 29184 2246 29236 2252
rect 29196 480 29224 2246
rect 26514 368 26570 377
rect 26514 303 26570 312
rect 27710 0 27766 480
rect 29182 0 29238 480
<< via2 >>
rect 2778 23568 2834 23624
rect 1122 16360 1178 16416
rect 2042 14048 2098 14104
rect 24950 23568 25006 23624
rect 3054 23024 3110 23080
rect 3422 22344 3478 22400
rect 4342 21800 4398 21856
rect 2962 21256 3018 21312
rect 3330 20576 3386 20632
rect 2870 20032 2926 20088
rect 1582 11600 1638 11656
rect 1582 10376 1638 10432
rect 1674 9968 1730 10024
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 2042 9016 2098 9072
rect 1582 8608 1638 8664
rect 662 7792 718 7848
rect 1582 7384 1638 7440
rect 1582 6840 1638 6896
rect 1398 6704 1454 6760
rect 2042 7268 2098 7304
rect 2042 7248 2044 7268
rect 2044 7248 2096 7268
rect 2096 7248 2098 7268
rect 2134 7112 2190 7168
rect 1582 6296 1638 6352
rect 1582 5616 1638 5672
rect 1582 5072 1638 5128
rect 2042 5092 2098 5128
rect 2042 5072 2044 5092
rect 2044 5072 2096 5092
rect 2096 5072 2098 5092
rect 3146 18264 3202 18320
rect 3054 18028 3056 18048
rect 3056 18028 3108 18048
rect 3108 18028 3110 18048
rect 3054 17992 3110 18028
rect 2778 13812 2780 13832
rect 2780 13812 2832 13832
rect 2832 13812 2834 13832
rect 2778 13776 2834 13812
rect 2870 13640 2926 13696
rect 2870 12824 2926 12880
rect 2594 11600 2650 11656
rect 4066 19352 4122 19408
rect 3514 18300 3516 18320
rect 3516 18300 3568 18320
rect 3568 18300 3570 18320
rect 3514 18264 3570 18300
rect 4066 17720 4122 17776
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 7470 20304 7526 20360
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 8206 18692 8262 18728
rect 8206 18672 8208 18692
rect 8208 18672 8260 18692
rect 8260 18672 8262 18692
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 4802 17040 4858 17096
rect 4342 16496 4398 16552
rect 3238 11464 3294 11520
rect 2686 9832 2742 9888
rect 2594 8064 2650 8120
rect 2502 6160 2558 6216
rect 1398 3304 1454 3360
rect 2502 3848 2558 3904
rect 2410 3576 2466 3632
rect 1582 2624 1638 2680
rect 2870 6840 2926 6896
rect 2870 5616 2926 5672
rect 2778 4392 2834 4448
rect 1766 1400 1822 1456
rect 2870 2080 2926 2136
rect 3238 9580 3294 9616
rect 3238 9560 3240 9580
rect 3240 9560 3292 9580
rect 3292 9560 3294 9580
rect 3790 15272 3846 15328
rect 3698 14356 3700 14376
rect 3700 14356 3752 14376
rect 3752 14356 3754 14376
rect 3698 14320 3754 14356
rect 3606 13948 3608 13968
rect 3608 13948 3660 13968
rect 3660 13948 3662 13968
rect 3606 13912 3662 13948
rect 3606 12280 3662 12336
rect 3698 8336 3754 8392
rect 3514 7928 3570 7984
rect 3238 6196 3240 6216
rect 3240 6196 3292 6216
rect 3292 6196 3294 6216
rect 3238 6160 3294 6196
rect 3146 4936 3202 4992
rect 3238 4020 3240 4040
rect 3240 4020 3292 4040
rect 3292 4020 3294 4040
rect 3238 3984 3294 4020
rect 4158 11056 4214 11112
rect 3882 9424 3938 9480
rect 3790 5888 3846 5944
rect 4434 15816 4490 15872
rect 4618 13368 4674 13424
rect 4618 10548 4620 10568
rect 4620 10548 4672 10568
rect 4672 10548 4674 10568
rect 4618 10512 4674 10548
rect 4618 7404 4674 7440
rect 4618 7384 4620 7404
rect 4620 7384 4672 7404
rect 4672 7384 4674 7404
rect 4618 7112 4674 7168
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5722 14592 5778 14648
rect 5630 13388 5686 13424
rect 5630 13368 5632 13388
rect 5632 13368 5684 13388
rect 5684 13368 5686 13388
rect 5170 12144 5226 12200
rect 5078 3440 5134 3496
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 6458 14048 6514 14104
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 5538 9968 5594 10024
rect 5354 8880 5410 8936
rect 5354 5208 5410 5264
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 7194 14764 7196 14784
rect 7196 14764 7248 14784
rect 7248 14764 7250 14784
rect 7194 14728 7250 14764
rect 7286 12180 7288 12200
rect 7288 12180 7340 12200
rect 7340 12180 7342 12200
rect 7286 12144 7342 12180
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 9770 18708 9772 18728
rect 9772 18708 9824 18728
rect 9824 18708 9826 18728
rect 9770 18672 9826 18708
rect 11794 18672 11850 18728
rect 9310 17584 9366 17640
rect 9310 17176 9366 17232
rect 9494 17040 9550 17096
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 11794 18128 11850 18184
rect 8666 16652 8722 16688
rect 8666 16632 8668 16652
rect 8668 16632 8720 16652
rect 8720 16632 8722 16652
rect 8114 15408 8170 15464
rect 8206 13776 8262 13832
rect 5630 3596 5686 3632
rect 5630 3576 5632 3596
rect 5632 3576 5684 3596
rect 5684 3576 5686 3596
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 6826 9152 6882 9208
rect 6366 8336 6422 8392
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 7286 7520 7342 7576
rect 6826 6704 6882 6760
rect 6366 3440 6422 3496
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 5814 2760 5870 2816
rect 2962 856 3018 912
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 7102 5208 7158 5264
rect 7010 4972 7012 4992
rect 7012 4972 7064 4992
rect 7064 4972 7066 4992
rect 7010 4936 7066 4972
rect 8022 5908 8078 5944
rect 8022 5888 8024 5908
rect 8024 5888 8076 5908
rect 8076 5888 8078 5908
rect 7930 5480 7986 5536
rect 8390 9560 8446 9616
rect 11610 17176 11666 17232
rect 9586 14864 9642 14920
rect 8850 13912 8906 13968
rect 9862 14864 9918 14920
rect 10046 13912 10102 13968
rect 10598 14456 10654 14512
rect 10138 13640 10194 13696
rect 10598 11500 10600 11520
rect 10600 11500 10652 11520
rect 10652 11500 10654 11520
rect 10598 11464 10654 11500
rect 9218 10648 9274 10704
rect 9954 9832 10010 9888
rect 9494 9016 9550 9072
rect 9862 7928 9918 7984
rect 8666 6568 8722 6624
rect 8206 6432 8262 6488
rect 9770 6724 9826 6760
rect 9770 6704 9772 6724
rect 9772 6704 9824 6724
rect 9824 6704 9826 6724
rect 9770 6568 9826 6624
rect 8574 5364 8630 5400
rect 8574 5344 8576 5364
rect 8576 5344 8628 5364
rect 8628 5344 8630 5364
rect 10322 7964 10324 7984
rect 10324 7964 10376 7984
rect 10376 7964 10378 7984
rect 10322 7928 10378 7964
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 11610 16088 11666 16144
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 11334 14612 11390 14648
rect 11334 14592 11336 14612
rect 11336 14592 11388 14612
rect 11388 14592 11390 14612
rect 10782 14456 10838 14512
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 11702 13504 11758 13560
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 10690 9152 10746 9208
rect 11334 10512 11390 10568
rect 11518 10512 11574 10568
rect 11334 10412 11336 10432
rect 11336 10412 11388 10432
rect 11388 10412 11390 10432
rect 11334 10376 11390 10412
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 11518 9968 11574 10024
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 10874 6704 10930 6760
rect 10506 6296 10562 6352
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 10046 5652 10048 5672
rect 10048 5652 10100 5672
rect 10100 5652 10102 5672
rect 10046 5616 10102 5652
rect 9954 5072 10010 5128
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 10138 4276 10194 4312
rect 10138 4256 10140 4276
rect 10140 4256 10192 4276
rect 10192 4256 10194 4276
rect 8390 4004 8446 4040
rect 8390 3984 8392 4004
rect 8392 3984 8444 4004
rect 8444 3984 8446 4004
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 9218 2760 9274 2816
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 13542 15988 13544 16008
rect 13544 15988 13596 16008
rect 13596 15988 13598 16008
rect 13542 15952 13598 15988
rect 13266 14492 13268 14512
rect 13268 14492 13320 14512
rect 13320 14492 13322 14512
rect 13266 14456 13322 14492
rect 13174 14048 13230 14104
rect 12622 13912 12678 13968
rect 12254 13640 12310 13696
rect 12346 9288 12402 9344
rect 11794 6160 11850 6216
rect 12162 5364 12218 5400
rect 12162 5344 12164 5364
rect 12164 5344 12216 5364
rect 12216 5344 12218 5364
rect 12162 4528 12218 4584
rect 12254 4256 12310 4312
rect 13082 13504 13138 13560
rect 13910 14592 13966 14648
rect 13818 13640 13874 13696
rect 13082 12552 13138 12608
rect 12622 9560 12678 9616
rect 12530 7928 12586 7984
rect 12806 9324 12808 9344
rect 12808 9324 12860 9344
rect 12860 9324 12862 9344
rect 12806 9288 12862 9324
rect 13174 9036 13230 9072
rect 13174 9016 13176 9036
rect 13176 9016 13228 9036
rect 13228 9016 13230 9036
rect 12806 6432 12862 6488
rect 12530 5480 12586 5536
rect 12806 4528 12862 4584
rect 13174 5480 13230 5536
rect 14186 14764 14188 14784
rect 14188 14764 14240 14784
rect 14240 14764 14242 14784
rect 14186 14728 14242 14764
rect 15474 18148 15530 18184
rect 15474 18128 15476 18148
rect 15476 18128 15528 18148
rect 15528 18128 15530 18148
rect 14922 17196 14978 17232
rect 14922 17176 14924 17196
rect 14924 17176 14976 17196
rect 14976 17176 14978 17196
rect 15566 17040 15622 17096
rect 14002 13640 14058 13696
rect 14002 10376 14058 10432
rect 14370 10684 14372 10704
rect 14372 10684 14424 10704
rect 14424 10684 14426 10704
rect 14370 10648 14426 10684
rect 14186 8880 14242 8936
rect 13450 7656 13506 7712
rect 13358 6060 13360 6080
rect 13360 6060 13412 6080
rect 13412 6060 13414 6080
rect 13358 6024 13414 6060
rect 13818 6740 13820 6760
rect 13820 6740 13872 6760
rect 13872 6740 13874 6760
rect 13818 6704 13874 6740
rect 14186 5072 14242 5128
rect 13450 3984 13506 4040
rect 14554 12280 14610 12336
rect 14646 9988 14702 10024
rect 14646 9968 14648 9988
rect 14648 9968 14700 9988
rect 14700 9968 14702 9988
rect 15382 13640 15438 13696
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 15750 18808 15806 18864
rect 17682 18536 17738 18592
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 16394 17312 16450 17368
rect 15842 17176 15898 17232
rect 15934 17040 15990 17096
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 16394 16904 16450 16960
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 16394 14728 16450 14784
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 16394 14048 16450 14104
rect 15750 13932 15806 13968
rect 15750 13912 15752 13932
rect 15752 13912 15804 13932
rect 15804 13912 15806 13932
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 16394 11872 16450 11928
rect 16486 11736 16542 11792
rect 16302 11620 16358 11656
rect 16302 11600 16304 11620
rect 16304 11600 16356 11620
rect 16356 11600 16358 11620
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15014 7384 15070 7440
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 16670 17176 16726 17232
rect 17130 15952 17186 16008
rect 17222 15408 17278 15464
rect 16486 10104 16542 10160
rect 15750 8336 15806 8392
rect 15474 7520 15530 7576
rect 15566 6196 15568 6216
rect 15568 6196 15620 6216
rect 15620 6196 15622 6216
rect 15566 6160 15622 6196
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 15934 8356 15990 8392
rect 15934 8336 15936 8356
rect 15936 8336 15988 8356
rect 15988 8336 15990 8356
rect 16302 7928 16358 7984
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 17406 14320 17462 14376
rect 16762 10648 16818 10704
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 19062 19216 19118 19272
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 17498 10920 17554 10976
rect 17314 10104 17370 10160
rect 17130 9288 17186 9344
rect 17038 7828 17040 7848
rect 17040 7828 17092 7848
rect 17092 7828 17094 7848
rect 17038 7792 17094 7828
rect 16394 7520 16450 7576
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 16670 7656 16726 7712
rect 18050 9560 18106 9616
rect 18970 17448 19026 17504
rect 18326 16496 18382 16552
rect 20810 17992 20866 18048
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 19522 16496 19578 16552
rect 19614 16088 19670 16144
rect 18418 15000 18474 15056
rect 18510 14884 18566 14920
rect 18510 14864 18512 14884
rect 18512 14864 18564 14884
rect 18564 14864 18566 14884
rect 18326 13912 18382 13968
rect 18234 13776 18290 13832
rect 18418 11872 18474 11928
rect 18326 9596 18328 9616
rect 18328 9596 18380 9616
rect 18380 9596 18382 9616
rect 18326 9560 18382 9596
rect 18142 9424 18198 9480
rect 17314 7248 17370 7304
rect 18878 13232 18934 13288
rect 18878 10512 18934 10568
rect 18510 9016 18566 9072
rect 18786 9324 18788 9344
rect 18788 9324 18840 9344
rect 18840 9324 18842 9344
rect 18786 9288 18842 9324
rect 19522 12960 19578 13016
rect 19522 12552 19578 12608
rect 19430 9424 19486 9480
rect 18878 8372 18880 8392
rect 18880 8372 18932 8392
rect 18932 8372 18934 8392
rect 18878 8336 18934 8372
rect 14646 3984 14702 4040
rect 13726 2760 13782 2816
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 16394 6296 16450 6352
rect 16302 5208 16358 5264
rect 15474 3848 15530 3904
rect 18050 5208 18106 5264
rect 16486 4664 16542 4720
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 17958 3984 18014 4040
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 16302 2760 16358 2816
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 19154 7792 19210 7848
rect 18878 6704 18934 6760
rect 19246 6860 19302 6896
rect 19246 6840 19248 6860
rect 19248 6840 19300 6860
rect 19300 6840 19302 6860
rect 19706 11620 19762 11656
rect 19706 11600 19708 11620
rect 19708 11600 19760 11620
rect 19760 11600 19762 11620
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 20718 14592 20774 14648
rect 21178 13812 21180 13832
rect 21180 13812 21232 13832
rect 21232 13812 21234 13832
rect 21178 13776 21234 13812
rect 20718 13640 20774 13696
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 21362 13776 21418 13832
rect 27526 23024 27582 23080
rect 25042 22344 25098 22400
rect 24950 18536 25006 18592
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25686 21528 25742 21584
rect 25502 21256 25558 21312
rect 25410 18808 25466 18864
rect 24858 18264 24914 18320
rect 24766 17040 24822 17096
rect 22742 15816 22798 15872
rect 21822 14068 21878 14104
rect 21822 14048 21824 14068
rect 21824 14048 21876 14068
rect 21876 14048 21878 14068
rect 21730 13776 21786 13832
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 19890 10376 19946 10432
rect 19798 8744 19854 8800
rect 19522 6296 19578 6352
rect 19062 5344 19118 5400
rect 18878 3884 18880 3904
rect 18880 3884 18932 3904
rect 18932 3884 18934 3904
rect 18878 3848 18934 3884
rect 18602 3032 18658 3088
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 21362 8880 21418 8936
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 19246 4664 19302 4720
rect 19890 3984 19946 4040
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 19614 3576 19670 3632
rect 19430 2932 19432 2952
rect 19432 2932 19484 2952
rect 19484 2932 19486 2952
rect 19430 2896 19486 2932
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 21914 13232 21970 13288
rect 22006 12824 22062 12880
rect 23938 12844 23994 12880
rect 23938 12824 23940 12844
rect 23940 12824 23992 12844
rect 23992 12824 23994 12844
rect 23294 11600 23350 11656
rect 23294 8744 23350 8800
rect 23202 8336 23258 8392
rect 23110 7656 23166 7712
rect 23110 7148 23112 7168
rect 23112 7148 23164 7168
rect 23164 7148 23166 7168
rect 23110 7112 23166 7148
rect 22650 6840 22706 6896
rect 23478 6296 23534 6352
rect 23202 6160 23258 6216
rect 22742 5364 22798 5400
rect 22742 5344 22744 5364
rect 22744 5344 22796 5364
rect 22796 5344 22798 5364
rect 23938 7520 23994 7576
rect 24214 13640 24270 13696
rect 24214 12960 24270 13016
rect 24766 12300 24822 12336
rect 24766 12280 24768 12300
rect 24768 12280 24820 12300
rect 24820 12280 24822 12300
rect 24490 11736 24546 11792
rect 24950 15408 25006 15464
rect 25410 17992 25466 18048
rect 25226 17312 25282 17368
rect 25594 17992 25650 18048
rect 25226 17040 25282 17096
rect 25042 13504 25098 13560
rect 25502 17040 25558 17096
rect 25226 13776 25282 13832
rect 25318 13268 25320 13288
rect 25320 13268 25372 13288
rect 25372 13268 25374 13288
rect 25318 13232 25374 13268
rect 25134 12416 25190 12472
rect 25226 12280 25282 12336
rect 25042 10104 25098 10160
rect 24950 9288 25006 9344
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 25870 20440 25926 20496
rect 25778 20032 25834 20088
rect 25778 18672 25834 18728
rect 25962 20304 26018 20360
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25686 17448 25742 17504
rect 26974 17992 27030 18048
rect 27526 17992 27582 18048
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 26790 17212 26792 17232
rect 26792 17212 26844 17232
rect 26844 17212 26846 17232
rect 26790 17176 26846 17212
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25778 16088 25834 16144
rect 26422 15544 26478 15600
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25778 15000 25834 15056
rect 25778 14592 25834 14648
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 25778 13368 25834 13424
rect 25410 11736 25466 11792
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25594 11872 25650 11928
rect 25318 10104 25374 10160
rect 25226 9968 25282 10024
rect 25226 9560 25282 9616
rect 25594 10920 25650 10976
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 26514 14864 26570 14920
rect 26606 12824 26662 12880
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 26422 10648 26478 10704
rect 26606 11600 26662 11656
rect 26698 11056 26754 11112
rect 26606 10376 26662 10432
rect 25686 8744 25742 8800
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 25778 8336 25834 8392
rect 25502 7384 25558 7440
rect 25686 6160 25742 6216
rect 24950 5752 25006 5808
rect 24306 5208 24362 5264
rect 24306 4528 24362 4584
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 26698 9832 26754 9888
rect 26514 9036 26570 9072
rect 26514 9016 26516 9036
rect 26516 9016 26568 9036
rect 26568 9016 26570 9036
rect 26698 8608 26754 8664
rect 27250 14048 27306 14104
rect 27250 13776 27306 13832
rect 27066 9424 27122 9480
rect 26790 8336 26846 8392
rect 26514 7792 26570 7848
rect 26514 7112 26570 7168
rect 26698 6840 26754 6896
rect 26606 6332 26608 6352
rect 26608 6332 26660 6352
rect 26660 6332 26662 6352
rect 26606 6296 26662 6332
rect 27158 9288 27214 9344
rect 27434 8064 27490 8120
rect 27618 8064 27674 8120
rect 27434 5752 27490 5808
rect 26698 5636 26754 5672
rect 26698 5616 26700 5636
rect 26700 5616 26752 5636
rect 26752 5616 26754 5636
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 26514 5208 26570 5264
rect 26422 5108 26424 5128
rect 26424 5108 26476 5128
rect 26476 5108 26478 5128
rect 26422 5072 26478 5108
rect 26606 5072 26662 5128
rect 25778 4528 25834 4584
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 26514 3596 26570 3632
rect 26514 3576 26516 3596
rect 26516 3576 26568 3596
rect 26568 3576 26570 3596
rect 26422 3440 26478 3496
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 26238 3032 26294 3088
rect 26330 2932 26332 2952
rect 26332 2932 26384 2952
rect 26384 2932 26386 2952
rect 26330 2896 26386 2932
rect 26698 3304 26754 3360
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 25870 856 25926 912
rect 2778 312 2834 368
rect 26606 2760 26662 2816
rect 27526 4020 27528 4040
rect 27528 4020 27580 4040
rect 27580 4020 27582 4040
rect 27526 3984 27582 4020
rect 27710 3884 27712 3904
rect 27712 3884 27764 3904
rect 27764 3884 27766 3904
rect 27710 3848 27766 3884
rect 29182 17584 29238 17640
rect 27618 2080 27674 2136
rect 26790 1400 26846 1456
rect 26514 312 26570 368
<< metal3 >>
rect 0 23626 480 23656
rect 2773 23626 2839 23629
rect 0 23624 2839 23626
rect 0 23568 2778 23624
rect 2834 23568 2839 23624
rect 0 23566 2839 23568
rect 0 23536 480 23566
rect 2773 23563 2839 23566
rect 24945 23626 25011 23629
rect 29520 23626 30000 23656
rect 24945 23624 30000 23626
rect 24945 23568 24950 23624
rect 25006 23568 30000 23624
rect 24945 23566 30000 23568
rect 24945 23563 25011 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 3049 23082 3115 23085
rect 0 23080 3115 23082
rect 0 23024 3054 23080
rect 3110 23024 3115 23080
rect 0 23022 3115 23024
rect 0 22992 480 23022
rect 3049 23019 3115 23022
rect 27521 23082 27587 23085
rect 29520 23082 30000 23112
rect 27521 23080 30000 23082
rect 27521 23024 27526 23080
rect 27582 23024 30000 23080
rect 27521 23022 30000 23024
rect 27521 23019 27587 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 3417 22402 3483 22405
rect 0 22400 3483 22402
rect 0 22344 3422 22400
rect 3478 22344 3483 22400
rect 0 22342 3483 22344
rect 0 22312 480 22342
rect 3417 22339 3483 22342
rect 25037 22402 25103 22405
rect 29520 22402 30000 22432
rect 25037 22400 30000 22402
rect 25037 22344 25042 22400
rect 25098 22344 30000 22400
rect 25037 22342 30000 22344
rect 25037 22339 25103 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 4337 21858 4403 21861
rect 29520 21858 30000 21888
rect 0 21856 4403 21858
rect 0 21800 4342 21856
rect 4398 21800 4403 21856
rect 0 21798 4403 21800
rect 0 21768 480 21798
rect 4337 21795 4403 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 25681 21586 25747 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 25681 21584 26434 21586
rect 25681 21528 25686 21584
rect 25742 21528 26434 21584
rect 25681 21526 26434 21528
rect 25681 21523 25747 21526
rect 0 21314 480 21344
rect 2957 21314 3023 21317
rect 0 21312 3023 21314
rect 0 21256 2962 21312
rect 3018 21256 3023 21312
rect 0 21254 3023 21256
rect 0 21224 480 21254
rect 2957 21251 3023 21254
rect 25497 21314 25563 21317
rect 29520 21314 30000 21344
rect 25497 21312 30000 21314
rect 25497 21256 25502 21312
rect 25558 21256 30000 21312
rect 25497 21254 30000 21256
rect 25497 21251 25563 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 3325 20634 3391 20637
rect 29520 20634 30000 20664
rect 0 20632 3391 20634
rect 0 20576 3330 20632
rect 3386 20576 3391 20632
rect 0 20574 3391 20576
rect 0 20544 480 20574
rect 3325 20571 3391 20574
rect 26374 20574 30000 20634
rect 25865 20498 25931 20501
rect 26374 20498 26434 20574
rect 29520 20544 30000 20574
rect 25865 20496 26434 20498
rect 25865 20440 25870 20496
rect 25926 20440 26434 20496
rect 25865 20438 26434 20440
rect 25865 20435 25931 20438
rect 7465 20362 7531 20365
rect 25957 20362 26023 20365
rect 7465 20360 26023 20362
rect 7465 20304 7470 20360
rect 7526 20304 25962 20360
rect 26018 20304 26023 20360
rect 7465 20302 26023 20304
rect 7465 20299 7531 20302
rect 25957 20299 26023 20302
rect 10944 20160 11264 20161
rect 0 20090 480 20120
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 2865 20090 2931 20093
rect 0 20088 2931 20090
rect 0 20032 2870 20088
rect 2926 20032 2931 20088
rect 0 20030 2931 20032
rect 0 20000 480 20030
rect 2865 20027 2931 20030
rect 25773 20090 25839 20093
rect 29520 20090 30000 20120
rect 25773 20088 30000 20090
rect 25773 20032 25778 20088
rect 25834 20032 30000 20088
rect 25773 20030 30000 20032
rect 25773 20027 25839 20030
rect 29520 20000 30000 20030
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 0 19410 480 19440
rect 4061 19410 4127 19413
rect 29520 19410 30000 19440
rect 0 19408 4127 19410
rect 0 19352 4066 19408
rect 4122 19352 4127 19408
rect 0 19350 4127 19352
rect 0 19320 480 19350
rect 4061 19347 4127 19350
rect 25040 19350 30000 19410
rect 19057 19274 19123 19277
rect 25040 19274 25100 19350
rect 29520 19320 30000 19350
rect 19057 19272 25100 19274
rect 19057 19216 19062 19272
rect 19118 19216 25100 19272
rect 19057 19214 25100 19216
rect 19057 19211 19123 19214
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 0 18866 480 18896
rect 15745 18866 15811 18869
rect 0 18864 15811 18866
rect 0 18808 15750 18864
rect 15806 18808 15811 18864
rect 0 18806 15811 18808
rect 0 18776 480 18806
rect 15745 18803 15811 18806
rect 25405 18866 25471 18869
rect 29520 18866 30000 18896
rect 25405 18864 30000 18866
rect 25405 18808 25410 18864
rect 25466 18808 30000 18864
rect 25405 18806 30000 18808
rect 25405 18803 25471 18806
rect 29520 18776 30000 18806
rect 8201 18730 8267 18733
rect 9765 18730 9831 18733
rect 8201 18728 9831 18730
rect 8201 18672 8206 18728
rect 8262 18672 9770 18728
rect 9826 18672 9831 18728
rect 8201 18670 9831 18672
rect 8201 18667 8267 18670
rect 9765 18667 9831 18670
rect 11789 18730 11855 18733
rect 25773 18730 25839 18733
rect 11789 18728 25839 18730
rect 11789 18672 11794 18728
rect 11850 18672 25778 18728
rect 25834 18672 25839 18728
rect 11789 18670 25839 18672
rect 11789 18667 11855 18670
rect 25773 18667 25839 18670
rect 17677 18594 17743 18597
rect 24945 18594 25011 18597
rect 17358 18592 25011 18594
rect 17358 18536 17682 18592
rect 17738 18536 24950 18592
rect 25006 18536 25011 18592
rect 17358 18534 25011 18536
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 0 18322 480 18352
rect 3141 18322 3207 18325
rect 0 18320 3207 18322
rect 0 18264 3146 18320
rect 3202 18264 3207 18320
rect 0 18262 3207 18264
rect 0 18232 480 18262
rect 3141 18259 3207 18262
rect 3509 18322 3575 18325
rect 17358 18322 17418 18534
rect 17677 18531 17743 18534
rect 24945 18531 25011 18534
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 3509 18320 17418 18322
rect 3509 18264 3514 18320
rect 3570 18264 17418 18320
rect 3509 18262 17418 18264
rect 24853 18322 24919 18325
rect 29520 18322 30000 18352
rect 24853 18320 30000 18322
rect 24853 18264 24858 18320
rect 24914 18264 30000 18320
rect 24853 18262 30000 18264
rect 3509 18259 3575 18262
rect 24853 18259 24919 18262
rect 29520 18232 30000 18262
rect 11789 18186 11855 18189
rect 5168 18184 11855 18186
rect 5168 18128 11794 18184
rect 11850 18128 11855 18184
rect 5168 18126 11855 18128
rect 3049 18050 3115 18053
rect 5168 18050 5228 18126
rect 11789 18123 11855 18126
rect 15469 18186 15535 18189
rect 15469 18184 25882 18186
rect 15469 18128 15474 18184
rect 15530 18128 25882 18184
rect 15469 18126 25882 18128
rect 15469 18123 15535 18126
rect 20805 18050 20871 18053
rect 3049 18048 5228 18050
rect 3049 17992 3054 18048
rect 3110 17992 5228 18048
rect 3049 17990 5228 17992
rect 19382 18048 20871 18050
rect 19382 17992 20810 18048
rect 20866 17992 20871 18048
rect 19382 17990 20871 17992
rect 3049 17987 3115 17990
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 19382 17914 19442 17990
rect 20805 17987 20871 17990
rect 25405 18050 25471 18053
rect 25589 18050 25655 18053
rect 25405 18048 25655 18050
rect 25405 17992 25410 18048
rect 25466 17992 25594 18048
rect 25650 17992 25655 18048
rect 25405 17990 25655 17992
rect 25822 18050 25882 18126
rect 26969 18050 27035 18053
rect 27521 18050 27587 18053
rect 25822 18048 27587 18050
rect 25822 17992 26974 18048
rect 27030 17992 27526 18048
rect 27582 17992 27587 18048
rect 25822 17990 27587 17992
rect 25405 17987 25471 17990
rect 25589 17987 25655 17990
rect 26969 17987 27035 17990
rect 27521 17987 27587 17990
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 14414 17854 19442 17914
rect 4061 17778 4127 17781
rect 14414 17778 14474 17854
rect 4061 17776 14474 17778
rect 4061 17720 4066 17776
rect 4122 17720 14474 17776
rect 4061 17718 14474 17720
rect 4061 17715 4127 17718
rect 0 17642 480 17672
rect 9305 17642 9371 17645
rect 0 17640 9371 17642
rect 0 17584 9310 17640
rect 9366 17584 9371 17640
rect 0 17582 9371 17584
rect 0 17552 480 17582
rect 9305 17579 9371 17582
rect 29177 17642 29243 17645
rect 29520 17642 30000 17672
rect 29177 17640 30000 17642
rect 29177 17584 29182 17640
rect 29238 17584 30000 17640
rect 29177 17582 30000 17584
rect 29177 17579 29243 17582
rect 29520 17552 30000 17582
rect 18965 17506 19031 17509
rect 25681 17506 25747 17509
rect 18965 17504 25747 17506
rect 18965 17448 18970 17504
rect 19026 17448 25686 17504
rect 25742 17448 25747 17504
rect 18965 17446 25747 17448
rect 18965 17443 19031 17446
rect 25681 17443 25747 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 16389 17370 16455 17373
rect 25221 17370 25287 17373
rect 16389 17368 25287 17370
rect 16389 17312 16394 17368
rect 16450 17312 25226 17368
rect 25282 17312 25287 17368
rect 16389 17310 25287 17312
rect 16389 17307 16455 17310
rect 25221 17307 25287 17310
rect 9305 17234 9371 17237
rect 11605 17234 11671 17237
rect 9305 17232 11671 17234
rect 9305 17176 9310 17232
rect 9366 17176 11610 17232
rect 11666 17176 11671 17232
rect 9305 17174 11671 17176
rect 9305 17171 9371 17174
rect 11605 17171 11671 17174
rect 14917 17234 14983 17237
rect 15837 17234 15903 17237
rect 16665 17234 16731 17237
rect 14917 17232 16731 17234
rect 14917 17176 14922 17232
rect 14978 17176 15842 17232
rect 15898 17176 16670 17232
rect 16726 17176 16731 17232
rect 14917 17174 16731 17176
rect 25224 17234 25284 17307
rect 26785 17234 26851 17237
rect 25224 17232 26851 17234
rect 25224 17176 26790 17232
rect 26846 17176 26851 17232
rect 25224 17174 26851 17176
rect 14917 17171 14983 17174
rect 15837 17171 15903 17174
rect 16665 17171 16731 17174
rect 26785 17171 26851 17174
rect 0 17098 480 17128
rect 4797 17098 4863 17101
rect 0 17096 4863 17098
rect 0 17040 4802 17096
rect 4858 17040 4863 17096
rect 0 17038 4863 17040
rect 0 17008 480 17038
rect 4797 17035 4863 17038
rect 9489 17098 9555 17101
rect 15561 17098 15627 17101
rect 15929 17098 15995 17101
rect 24761 17098 24827 17101
rect 25221 17098 25287 17101
rect 9489 17096 15808 17098
rect 9489 17040 9494 17096
rect 9550 17040 15566 17096
rect 15622 17040 15808 17096
rect 9489 17038 15808 17040
rect 9489 17035 9555 17038
rect 15561 17035 15627 17038
rect 15748 16962 15808 17038
rect 15929 17096 25287 17098
rect 15929 17040 15934 17096
rect 15990 17040 24766 17096
rect 24822 17040 25226 17096
rect 25282 17040 25287 17096
rect 15929 17038 25287 17040
rect 15929 17035 15995 17038
rect 24761 17035 24827 17038
rect 25221 17035 25287 17038
rect 25497 17098 25563 17101
rect 29520 17098 30000 17128
rect 25497 17096 30000 17098
rect 25497 17040 25502 17096
rect 25558 17040 30000 17096
rect 25497 17038 30000 17040
rect 25497 17035 25563 17038
rect 29520 17008 30000 17038
rect 16389 16962 16455 16965
rect 15748 16960 16455 16962
rect 15748 16904 16394 16960
rect 16450 16904 16455 16960
rect 15748 16902 16455 16904
rect 16389 16899 16455 16902
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 8661 16690 8727 16693
rect 8661 16688 19580 16690
rect 8661 16632 8666 16688
rect 8722 16632 19580 16688
rect 8661 16630 19580 16632
rect 8661 16627 8727 16630
rect 19520 16557 19580 16630
rect 4337 16554 4403 16557
rect 18321 16554 18387 16557
rect 4337 16552 18387 16554
rect 4337 16496 4342 16552
rect 4398 16496 18326 16552
rect 18382 16496 18387 16552
rect 4337 16494 18387 16496
rect 4337 16491 4403 16494
rect 18321 16491 18387 16494
rect 19517 16552 19583 16557
rect 19517 16496 19522 16552
rect 19578 16496 19583 16552
rect 19517 16491 19583 16496
rect 0 16418 480 16448
rect 1117 16418 1183 16421
rect 29520 16418 30000 16448
rect 0 16416 1183 16418
rect 0 16360 1122 16416
rect 1178 16360 1183 16416
rect 0 16358 1183 16360
rect 0 16328 480 16358
rect 1117 16355 1183 16358
rect 26374 16358 30000 16418
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 11605 16146 11671 16149
rect 19609 16146 19675 16149
rect 11605 16144 19675 16146
rect 11605 16088 11610 16144
rect 11666 16088 19614 16144
rect 19670 16088 19675 16144
rect 11605 16086 19675 16088
rect 11605 16083 11671 16086
rect 19609 16083 19675 16086
rect 25773 16146 25839 16149
rect 26374 16146 26434 16358
rect 29520 16328 30000 16358
rect 25773 16144 26434 16146
rect 25773 16088 25778 16144
rect 25834 16088 26434 16144
rect 25773 16086 26434 16088
rect 25773 16083 25839 16086
rect 13537 16010 13603 16013
rect 17125 16010 17191 16013
rect 13537 16008 17191 16010
rect 13537 15952 13542 16008
rect 13598 15952 17130 16008
rect 17186 15952 17191 16008
rect 13537 15950 17191 15952
rect 13537 15947 13603 15950
rect 17125 15947 17191 15950
rect 0 15874 480 15904
rect 4429 15874 4495 15877
rect 0 15872 4495 15874
rect 0 15816 4434 15872
rect 4490 15816 4495 15872
rect 0 15814 4495 15816
rect 0 15784 480 15814
rect 4429 15811 4495 15814
rect 22737 15874 22803 15877
rect 29520 15874 30000 15904
rect 22737 15872 30000 15874
rect 22737 15816 22742 15872
rect 22798 15816 30000 15872
rect 22737 15814 30000 15816
rect 22737 15811 22803 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 26417 15602 26483 15605
rect 24718 15600 26483 15602
rect 24718 15544 26422 15600
rect 26478 15544 26483 15600
rect 24718 15542 26483 15544
rect 8109 15466 8175 15469
rect 17217 15466 17283 15469
rect 24718 15466 24778 15542
rect 26417 15539 26483 15542
rect 8109 15464 24778 15466
rect 8109 15408 8114 15464
rect 8170 15408 17222 15464
rect 17278 15408 24778 15464
rect 8109 15406 24778 15408
rect 24945 15466 25011 15469
rect 24945 15464 26434 15466
rect 24945 15408 24950 15464
rect 25006 15408 26434 15464
rect 24945 15406 26434 15408
rect 8109 15403 8175 15406
rect 17217 15403 17283 15406
rect 24945 15403 25011 15406
rect 0 15330 480 15360
rect 3785 15330 3851 15333
rect 0 15328 3851 15330
rect 0 15272 3790 15328
rect 3846 15272 3851 15328
rect 0 15270 3851 15272
rect 26374 15330 26434 15406
rect 29520 15330 30000 15360
rect 26374 15270 30000 15330
rect 0 15240 480 15270
rect 3785 15267 3851 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 18413 15058 18479 15061
rect 25773 15058 25839 15061
rect 18413 15056 25839 15058
rect 18413 15000 18418 15056
rect 18474 15000 25778 15056
rect 25834 15000 25839 15056
rect 18413 14998 25839 15000
rect 18413 14995 18479 14998
rect 25773 14995 25839 14998
rect 9581 14922 9647 14925
rect 9857 14922 9923 14925
rect 9581 14920 9923 14922
rect 9581 14864 9586 14920
rect 9642 14864 9862 14920
rect 9918 14864 9923 14920
rect 9581 14862 9923 14864
rect 9581 14859 9647 14862
rect 9857 14859 9923 14862
rect 18505 14922 18571 14925
rect 26509 14922 26575 14925
rect 18505 14920 26575 14922
rect 18505 14864 18510 14920
rect 18566 14864 26514 14920
rect 26570 14864 26575 14920
rect 18505 14862 26575 14864
rect 18505 14859 18571 14862
rect 26509 14859 26575 14862
rect 7189 14786 7255 14789
rect 9622 14786 9628 14788
rect 7189 14784 9628 14786
rect 7189 14728 7194 14784
rect 7250 14728 9628 14784
rect 7189 14726 9628 14728
rect 7189 14723 7255 14726
rect 9622 14724 9628 14726
rect 9692 14724 9698 14788
rect 14181 14786 14247 14789
rect 16389 14786 16455 14789
rect 14181 14784 16455 14786
rect 14181 14728 14186 14784
rect 14242 14728 16394 14784
rect 16450 14728 16455 14784
rect 14181 14726 16455 14728
rect 14181 14723 14247 14726
rect 16389 14723 16455 14726
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 5717 14650 5783 14653
rect 0 14648 5783 14650
rect 0 14592 5722 14648
rect 5778 14592 5783 14648
rect 0 14590 5783 14592
rect 0 14560 480 14590
rect 5717 14587 5783 14590
rect 11329 14650 11395 14653
rect 13905 14650 13971 14653
rect 20713 14650 20779 14653
rect 11329 14648 20779 14650
rect 11329 14592 11334 14648
rect 11390 14592 13910 14648
rect 13966 14592 20718 14648
rect 20774 14592 20779 14648
rect 11329 14590 20779 14592
rect 11329 14587 11395 14590
rect 13905 14587 13971 14590
rect 20713 14587 20779 14590
rect 25773 14650 25839 14653
rect 29520 14650 30000 14680
rect 25773 14648 30000 14650
rect 25773 14592 25778 14648
rect 25834 14592 30000 14648
rect 25773 14590 30000 14592
rect 25773 14587 25839 14590
rect 29520 14560 30000 14590
rect 9622 14452 9628 14516
rect 9692 14514 9698 14516
rect 10593 14514 10659 14517
rect 9692 14512 10659 14514
rect 9692 14456 10598 14512
rect 10654 14456 10659 14512
rect 9692 14454 10659 14456
rect 9692 14452 9698 14454
rect 10593 14451 10659 14454
rect 10777 14514 10843 14517
rect 13261 14514 13327 14517
rect 10777 14512 13327 14514
rect 10777 14456 10782 14512
rect 10838 14456 13266 14512
rect 13322 14456 13327 14512
rect 10777 14454 13327 14456
rect 10777 14451 10843 14454
rect 13261 14451 13327 14454
rect 3693 14378 3759 14381
rect 17401 14378 17467 14381
rect 3693 14376 17467 14378
rect 3693 14320 3698 14376
rect 3754 14320 17406 14376
rect 17462 14320 17467 14376
rect 3693 14318 17467 14320
rect 3693 14315 3759 14318
rect 17401 14315 17467 14318
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 2037 14106 2103 14109
rect 0 14104 2103 14106
rect 0 14048 2042 14104
rect 2098 14048 2103 14104
rect 0 14046 2103 14048
rect 0 14016 480 14046
rect 2037 14043 2103 14046
rect 6453 14106 6519 14109
rect 13169 14106 13235 14109
rect 6453 14104 13235 14106
rect 6453 14048 6458 14104
rect 6514 14048 13174 14104
rect 13230 14048 13235 14104
rect 6453 14046 13235 14048
rect 6453 14043 6519 14046
rect 13169 14043 13235 14046
rect 16389 14106 16455 14109
rect 21817 14106 21883 14109
rect 16389 14104 21883 14106
rect 16389 14048 16394 14104
rect 16450 14048 21822 14104
rect 21878 14048 21883 14104
rect 16389 14046 21883 14048
rect 16389 14043 16455 14046
rect 21817 14043 21883 14046
rect 27245 14106 27311 14109
rect 29520 14106 30000 14136
rect 27245 14104 30000 14106
rect 27245 14048 27250 14104
rect 27306 14048 30000 14104
rect 27245 14046 30000 14048
rect 27245 14043 27311 14046
rect 29520 14016 30000 14046
rect 3601 13970 3667 13973
rect 8845 13970 8911 13973
rect 3601 13968 8911 13970
rect 3601 13912 3606 13968
rect 3662 13912 8850 13968
rect 8906 13912 8911 13968
rect 3601 13910 8911 13912
rect 3601 13907 3667 13910
rect 8845 13907 8911 13910
rect 10041 13970 10107 13973
rect 12617 13970 12683 13973
rect 10041 13968 12683 13970
rect 10041 13912 10046 13968
rect 10102 13912 12622 13968
rect 12678 13912 12683 13968
rect 10041 13910 12683 13912
rect 10041 13907 10107 13910
rect 12617 13907 12683 13910
rect 15745 13970 15811 13973
rect 18321 13970 18387 13973
rect 15745 13968 18387 13970
rect 15745 13912 15750 13968
rect 15806 13912 18326 13968
rect 18382 13912 18387 13968
rect 15745 13910 18387 13912
rect 15745 13907 15811 13910
rect 18321 13907 18387 13910
rect 2773 13834 2839 13837
rect 8201 13834 8267 13837
rect 2773 13832 8267 13834
rect 2773 13776 2778 13832
rect 2834 13776 8206 13832
rect 8262 13776 8267 13832
rect 2773 13774 8267 13776
rect 2773 13771 2839 13774
rect 8201 13771 8267 13774
rect 18229 13834 18295 13837
rect 21173 13834 21239 13837
rect 21357 13834 21423 13837
rect 18229 13832 21423 13834
rect 18229 13776 18234 13832
rect 18290 13776 21178 13832
rect 21234 13776 21362 13832
rect 21418 13776 21423 13832
rect 18229 13774 21423 13776
rect 18229 13771 18295 13774
rect 21173 13771 21239 13774
rect 21357 13771 21423 13774
rect 21725 13834 21791 13837
rect 25221 13834 25287 13837
rect 27245 13834 27311 13837
rect 21725 13832 25287 13834
rect 21725 13776 21730 13832
rect 21786 13776 25226 13832
rect 25282 13776 25287 13832
rect 21725 13774 25287 13776
rect 21725 13771 21791 13774
rect 25221 13771 25287 13774
rect 26006 13832 27311 13834
rect 26006 13776 27250 13832
rect 27306 13776 27311 13832
rect 26006 13774 27311 13776
rect 2865 13698 2931 13701
rect 10133 13698 10199 13701
rect 2865 13696 10199 13698
rect 2865 13640 2870 13696
rect 2926 13640 10138 13696
rect 10194 13640 10199 13696
rect 2865 13638 10199 13640
rect 2865 13635 2931 13638
rect 10133 13635 10199 13638
rect 12249 13698 12315 13701
rect 13813 13698 13879 13701
rect 12249 13696 13879 13698
rect 12249 13640 12254 13696
rect 12310 13640 13818 13696
rect 13874 13640 13879 13696
rect 12249 13638 13879 13640
rect 12249 13635 12315 13638
rect 13813 13635 13879 13638
rect 13997 13698 14063 13701
rect 15377 13698 15443 13701
rect 20713 13698 20779 13701
rect 13997 13696 20779 13698
rect 13997 13640 14002 13696
rect 14058 13640 15382 13696
rect 15438 13640 20718 13696
rect 20774 13640 20779 13696
rect 13997 13638 20779 13640
rect 13997 13635 14063 13638
rect 15377 13635 15443 13638
rect 20713 13635 20779 13638
rect 24209 13698 24275 13701
rect 26006 13698 26066 13774
rect 27245 13771 27311 13774
rect 24209 13696 26066 13698
rect 24209 13640 24214 13696
rect 24270 13640 26066 13696
rect 24209 13638 26066 13640
rect 24209 13635 24275 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 11697 13562 11763 13565
rect 13077 13562 13143 13565
rect 11697 13560 13143 13562
rect 11697 13504 11702 13560
rect 11758 13504 13082 13560
rect 13138 13504 13143 13560
rect 11697 13502 13143 13504
rect 11697 13499 11763 13502
rect 13077 13499 13143 13502
rect 25037 13562 25103 13565
rect 25037 13560 26066 13562
rect 25037 13504 25042 13560
rect 25098 13504 26066 13560
rect 25037 13502 26066 13504
rect 25037 13499 25103 13502
rect 0 13426 480 13456
rect 4613 13426 4679 13429
rect 0 13424 4679 13426
rect 0 13368 4618 13424
rect 4674 13368 4679 13424
rect 0 13366 4679 13368
rect 0 13336 480 13366
rect 4613 13363 4679 13366
rect 5625 13426 5691 13429
rect 25773 13426 25839 13429
rect 5625 13424 25839 13426
rect 5625 13368 5630 13424
rect 5686 13368 25778 13424
rect 25834 13368 25839 13424
rect 5625 13366 25839 13368
rect 26006 13426 26066 13502
rect 29520 13426 30000 13456
rect 26006 13366 30000 13426
rect 5625 13363 5691 13366
rect 25773 13363 25839 13366
rect 29520 13336 30000 13366
rect 18873 13290 18939 13293
rect 21909 13290 21975 13293
rect 25313 13290 25379 13293
rect 18873 13288 25379 13290
rect 18873 13232 18878 13288
rect 18934 13232 21914 13288
rect 21970 13232 25318 13288
rect 25374 13232 25379 13288
rect 18873 13230 25379 13232
rect 18873 13227 18939 13230
rect 21909 13227 21975 13230
rect 25313 13227 25379 13230
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 19517 13018 19583 13021
rect 24209 13018 24275 13021
rect 19517 13016 24275 13018
rect 19517 12960 19522 13016
rect 19578 12960 24214 13016
rect 24270 12960 24275 13016
rect 19517 12958 24275 12960
rect 19517 12955 19583 12958
rect 24209 12955 24275 12958
rect 0 12882 480 12912
rect 2865 12882 2931 12885
rect 0 12880 2931 12882
rect 0 12824 2870 12880
rect 2926 12824 2931 12880
rect 0 12822 2931 12824
rect 0 12792 480 12822
rect 2865 12819 2931 12822
rect 22001 12882 22067 12885
rect 23933 12882 23999 12885
rect 22001 12880 23999 12882
rect 22001 12824 22006 12880
rect 22062 12824 23938 12880
rect 23994 12824 23999 12880
rect 22001 12822 23999 12824
rect 22001 12819 22067 12822
rect 23933 12819 23999 12822
rect 26601 12882 26667 12885
rect 29520 12882 30000 12912
rect 26601 12880 30000 12882
rect 26601 12824 26606 12880
rect 26662 12824 30000 12880
rect 26601 12822 30000 12824
rect 26601 12819 26667 12822
rect 29520 12792 30000 12822
rect 13077 12610 13143 12613
rect 19517 12610 19583 12613
rect 13077 12608 19583 12610
rect 13077 12552 13082 12608
rect 13138 12552 19522 12608
rect 19578 12552 19583 12608
rect 13077 12550 19583 12552
rect 13077 12547 13143 12550
rect 19517 12547 19583 12550
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 25129 12476 25195 12477
rect 25078 12412 25084 12476
rect 25148 12474 25195 12476
rect 25148 12472 25240 12474
rect 25190 12416 25240 12472
rect 25148 12414 25240 12416
rect 25148 12412 25195 12414
rect 25129 12411 25195 12412
rect 0 12338 480 12368
rect 3601 12338 3667 12341
rect 0 12336 3667 12338
rect 0 12280 3606 12336
rect 3662 12280 3667 12336
rect 0 12278 3667 12280
rect 0 12248 480 12278
rect 3601 12275 3667 12278
rect 14549 12338 14615 12341
rect 24761 12338 24827 12341
rect 14549 12336 24827 12338
rect 14549 12280 14554 12336
rect 14610 12280 24766 12336
rect 24822 12280 24827 12336
rect 14549 12278 24827 12280
rect 14549 12275 14615 12278
rect 24761 12275 24827 12278
rect 25221 12338 25287 12341
rect 29520 12338 30000 12368
rect 25221 12336 30000 12338
rect 25221 12280 25226 12336
rect 25282 12280 30000 12336
rect 25221 12278 30000 12280
rect 25221 12275 25287 12278
rect 29520 12248 30000 12278
rect 5165 12202 5231 12205
rect 7281 12202 7347 12205
rect 5165 12200 7347 12202
rect 5165 12144 5170 12200
rect 5226 12144 7286 12200
rect 7342 12144 7347 12200
rect 5165 12142 7347 12144
rect 5165 12139 5231 12142
rect 7281 12139 7347 12142
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 16389 11930 16455 11933
rect 18413 11930 18479 11933
rect 25589 11930 25655 11933
rect 16389 11928 25655 11930
rect 16389 11872 16394 11928
rect 16450 11872 18418 11928
rect 18474 11872 25594 11928
rect 25650 11872 25655 11928
rect 16389 11870 25655 11872
rect 16389 11867 16455 11870
rect 18413 11867 18479 11870
rect 25589 11867 25655 11870
rect 16481 11794 16547 11797
rect 24485 11794 24551 11797
rect 25405 11794 25471 11797
rect 16481 11792 25471 11794
rect 16481 11736 16486 11792
rect 16542 11736 24490 11792
rect 24546 11736 25410 11792
rect 25466 11736 25471 11792
rect 16481 11734 25471 11736
rect 16481 11731 16547 11734
rect 24485 11731 24551 11734
rect 25405 11731 25471 11734
rect 0 11658 480 11688
rect 1577 11658 1643 11661
rect 0 11656 1643 11658
rect 0 11600 1582 11656
rect 1638 11600 1643 11656
rect 0 11598 1643 11600
rect 0 11568 480 11598
rect 1577 11595 1643 11598
rect 2589 11658 2655 11661
rect 16297 11658 16363 11661
rect 2589 11656 16363 11658
rect 2589 11600 2594 11656
rect 2650 11600 16302 11656
rect 16358 11600 16363 11656
rect 2589 11598 16363 11600
rect 2589 11595 2655 11598
rect 16297 11595 16363 11598
rect 19701 11658 19767 11661
rect 23289 11658 23355 11661
rect 19701 11656 23355 11658
rect 19701 11600 19706 11656
rect 19762 11600 23294 11656
rect 23350 11600 23355 11656
rect 19701 11598 23355 11600
rect 19701 11595 19767 11598
rect 23289 11595 23355 11598
rect 26601 11658 26667 11661
rect 29520 11658 30000 11688
rect 26601 11656 30000 11658
rect 26601 11600 26606 11656
rect 26662 11600 30000 11656
rect 26601 11598 30000 11600
rect 26601 11595 26667 11598
rect 29520 11568 30000 11598
rect 3233 11522 3299 11525
rect 10593 11522 10659 11525
rect 3233 11520 10659 11522
rect 3233 11464 3238 11520
rect 3294 11464 10598 11520
rect 10654 11464 10659 11520
rect 3233 11462 10659 11464
rect 3233 11459 3299 11462
rect 10593 11459 10659 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 0 11114 480 11144
rect 4153 11114 4219 11117
rect 0 11112 4219 11114
rect 0 11056 4158 11112
rect 4214 11056 4219 11112
rect 0 11054 4219 11056
rect 0 11024 480 11054
rect 4153 11051 4219 11054
rect 26693 11114 26759 11117
rect 29520 11114 30000 11144
rect 26693 11112 30000 11114
rect 26693 11056 26698 11112
rect 26754 11056 30000 11112
rect 26693 11054 30000 11056
rect 26693 11051 26759 11054
rect 29520 11024 30000 11054
rect 17493 10978 17559 10981
rect 25589 10978 25655 10981
rect 17493 10976 25655 10978
rect 17493 10920 17498 10976
rect 17554 10920 25594 10976
rect 25650 10920 25655 10976
rect 17493 10918 25655 10920
rect 17493 10915 17559 10918
rect 25589 10915 25655 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 9213 10706 9279 10709
rect 14365 10706 14431 10709
rect 16757 10706 16823 10709
rect 26417 10706 26483 10709
rect 9213 10704 14474 10706
rect 9213 10648 9218 10704
rect 9274 10648 14370 10704
rect 14426 10648 14474 10704
rect 9213 10646 14474 10648
rect 9213 10643 9279 10646
rect 14365 10643 14474 10646
rect 16757 10704 26483 10706
rect 16757 10648 16762 10704
rect 16818 10648 26422 10704
rect 26478 10648 26483 10704
rect 16757 10646 26483 10648
rect 16757 10643 16823 10646
rect 26417 10643 26483 10646
rect 4613 10570 4679 10573
rect 11329 10570 11395 10573
rect 4613 10568 11395 10570
rect 4613 10512 4618 10568
rect 4674 10512 11334 10568
rect 11390 10512 11395 10568
rect 4613 10510 11395 10512
rect 4613 10507 4679 10510
rect 11329 10507 11395 10510
rect 11513 10570 11579 10573
rect 14414 10570 14474 10643
rect 18873 10570 18939 10573
rect 11513 10568 14290 10570
rect 11513 10512 11518 10568
rect 11574 10512 14290 10568
rect 11513 10510 14290 10512
rect 14414 10568 18939 10570
rect 14414 10512 18878 10568
rect 18934 10512 18939 10568
rect 14414 10510 18939 10512
rect 11513 10507 11579 10510
rect 0 10434 480 10464
rect 1577 10434 1643 10437
rect 0 10432 1643 10434
rect 0 10376 1582 10432
rect 1638 10376 1643 10432
rect 0 10374 1643 10376
rect 0 10344 480 10374
rect 1577 10371 1643 10374
rect 11329 10434 11395 10437
rect 13997 10434 14063 10437
rect 11329 10432 14063 10434
rect 11329 10376 11334 10432
rect 11390 10376 14002 10432
rect 14058 10376 14063 10432
rect 11329 10374 14063 10376
rect 14230 10434 14290 10510
rect 18873 10507 18939 10510
rect 19885 10434 19951 10437
rect 14230 10432 19951 10434
rect 14230 10376 19890 10432
rect 19946 10376 19951 10432
rect 14230 10374 19951 10376
rect 11329 10371 11395 10374
rect 13997 10371 14063 10374
rect 19885 10371 19951 10374
rect 26601 10434 26667 10437
rect 29520 10434 30000 10464
rect 26601 10432 30000 10434
rect 26601 10376 26606 10432
rect 26662 10376 30000 10432
rect 26601 10374 30000 10376
rect 26601 10371 26667 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 16481 10162 16547 10165
rect 2868 10160 16547 10162
rect 2868 10104 16486 10160
rect 16542 10104 16547 10160
rect 2868 10102 16547 10104
rect 1669 10026 1735 10029
rect 2868 10026 2928 10102
rect 16481 10099 16547 10102
rect 17309 10162 17375 10165
rect 25037 10162 25103 10165
rect 25313 10162 25379 10165
rect 17309 10160 25379 10162
rect 17309 10104 17314 10160
rect 17370 10104 25042 10160
rect 25098 10104 25318 10160
rect 25374 10104 25379 10160
rect 17309 10102 25379 10104
rect 17309 10099 17375 10102
rect 25037 10099 25103 10102
rect 25313 10099 25379 10102
rect 1669 10024 2928 10026
rect 1669 9968 1674 10024
rect 1730 9968 2928 10024
rect 1669 9966 2928 9968
rect 5533 10026 5599 10029
rect 11513 10026 11579 10029
rect 14641 10026 14707 10029
rect 25221 10026 25287 10029
rect 5533 10024 11579 10026
rect 5533 9968 5538 10024
rect 5594 9968 11518 10024
rect 11574 9968 11579 10024
rect 5533 9966 11579 9968
rect 1669 9963 1735 9966
rect 5533 9963 5599 9966
rect 11513 9963 11579 9966
rect 14598 10024 25287 10026
rect 14598 9968 14646 10024
rect 14702 9968 25226 10024
rect 25282 9968 25287 10024
rect 14598 9966 25287 9968
rect 14598 9963 14707 9966
rect 25221 9963 25287 9966
rect 0 9890 480 9920
rect 2681 9890 2747 9893
rect 0 9888 2747 9890
rect 0 9832 2686 9888
rect 2742 9832 2747 9888
rect 0 9830 2747 9832
rect 0 9800 480 9830
rect 2681 9827 2747 9830
rect 9949 9890 10015 9893
rect 14598 9890 14658 9963
rect 9949 9888 14658 9890
rect 9949 9832 9954 9888
rect 10010 9832 14658 9888
rect 9949 9830 14658 9832
rect 26693 9890 26759 9893
rect 29520 9890 30000 9920
rect 26693 9888 30000 9890
rect 26693 9832 26698 9888
rect 26754 9832 30000 9888
rect 26693 9830 30000 9832
rect 9949 9827 10015 9830
rect 26693 9827 26759 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 3233 9618 3299 9621
rect 8385 9618 8451 9621
rect 3233 9616 8451 9618
rect 3233 9560 3238 9616
rect 3294 9560 8390 9616
rect 8446 9560 8451 9616
rect 3233 9558 8451 9560
rect 3233 9555 3299 9558
rect 8385 9555 8451 9558
rect 12617 9618 12683 9621
rect 18045 9618 18111 9621
rect 12617 9616 18111 9618
rect 12617 9560 12622 9616
rect 12678 9560 18050 9616
rect 18106 9560 18111 9616
rect 12617 9558 18111 9560
rect 12617 9555 12683 9558
rect 18045 9555 18111 9558
rect 18321 9618 18387 9621
rect 25221 9618 25287 9621
rect 18321 9616 25287 9618
rect 18321 9560 18326 9616
rect 18382 9560 25226 9616
rect 25282 9560 25287 9616
rect 18321 9558 25287 9560
rect 18321 9555 18387 9558
rect 25221 9555 25287 9558
rect 3877 9482 3943 9485
rect 18137 9482 18203 9485
rect 3877 9480 18203 9482
rect 3877 9424 3882 9480
rect 3938 9424 18142 9480
rect 18198 9424 18203 9480
rect 3877 9422 18203 9424
rect 3877 9419 3943 9422
rect 18137 9419 18203 9422
rect 19425 9482 19491 9485
rect 27061 9482 27127 9485
rect 19425 9480 27127 9482
rect 19425 9424 19430 9480
rect 19486 9424 27066 9480
rect 27122 9424 27127 9480
rect 19425 9422 27127 9424
rect 19425 9419 19491 9422
rect 27061 9419 27127 9422
rect 0 9346 480 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 480 9286
rect 1577 9283 1643 9286
rect 12341 9346 12407 9349
rect 12801 9346 12867 9349
rect 12341 9344 12867 9346
rect 12341 9288 12346 9344
rect 12402 9288 12806 9344
rect 12862 9288 12867 9344
rect 12341 9286 12867 9288
rect 12341 9283 12407 9286
rect 12801 9283 12867 9286
rect 17125 9346 17191 9349
rect 18781 9346 18847 9349
rect 17125 9344 18847 9346
rect 17125 9288 17130 9344
rect 17186 9288 18786 9344
rect 18842 9288 18847 9344
rect 17125 9286 18847 9288
rect 17125 9283 17191 9286
rect 18781 9283 18847 9286
rect 24945 9346 25011 9349
rect 25078 9346 25084 9348
rect 24945 9344 25084 9346
rect 24945 9288 24950 9344
rect 25006 9288 25084 9344
rect 24945 9286 25084 9288
rect 24945 9283 25011 9286
rect 25078 9284 25084 9286
rect 25148 9284 25154 9348
rect 27153 9346 27219 9349
rect 29520 9346 30000 9376
rect 27153 9344 30000 9346
rect 27153 9288 27158 9344
rect 27214 9288 30000 9344
rect 27153 9286 30000 9288
rect 27153 9283 27219 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 6821 9210 6887 9213
rect 10685 9210 10751 9213
rect 6821 9208 10751 9210
rect 6821 9152 6826 9208
rect 6882 9152 10690 9208
rect 10746 9152 10751 9208
rect 6821 9150 10751 9152
rect 6821 9147 6887 9150
rect 10685 9147 10751 9150
rect 2037 9074 2103 9077
rect 9489 9074 9555 9077
rect 2037 9072 9555 9074
rect 2037 9016 2042 9072
rect 2098 9016 9494 9072
rect 9550 9016 9555 9072
rect 2037 9014 9555 9016
rect 2037 9011 2103 9014
rect 9489 9011 9555 9014
rect 13169 9074 13235 9077
rect 18505 9074 18571 9077
rect 26509 9074 26575 9077
rect 13169 9072 17418 9074
rect 13169 9016 13174 9072
rect 13230 9016 17418 9072
rect 13169 9014 17418 9016
rect 13169 9011 13235 9014
rect 5349 8938 5415 8941
rect 14181 8938 14247 8941
rect 5349 8936 14247 8938
rect 5349 8880 5354 8936
rect 5410 8880 14186 8936
rect 14242 8880 14247 8936
rect 5349 8878 14247 8880
rect 17358 8938 17418 9014
rect 18505 9072 26575 9074
rect 18505 9016 18510 9072
rect 18566 9016 26514 9072
rect 26570 9016 26575 9072
rect 18505 9014 26575 9016
rect 18505 9011 18571 9014
rect 26509 9011 26575 9014
rect 21357 8938 21423 8941
rect 17358 8936 21423 8938
rect 17358 8880 21362 8936
rect 21418 8880 21423 8936
rect 17358 8878 21423 8880
rect 5349 8875 5415 8878
rect 14181 8875 14247 8878
rect 21357 8875 21423 8878
rect 19793 8802 19859 8805
rect 23289 8802 23355 8805
rect 25681 8802 25747 8805
rect 19793 8800 25747 8802
rect 19793 8744 19798 8800
rect 19854 8744 23294 8800
rect 23350 8744 25686 8800
rect 25742 8744 25747 8800
rect 19793 8742 25747 8744
rect 19793 8739 19859 8742
rect 23289 8739 23355 8742
rect 25681 8739 25747 8742
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 1577 8666 1643 8669
rect 0 8664 1643 8666
rect 0 8608 1582 8664
rect 1638 8608 1643 8664
rect 0 8606 1643 8608
rect 0 8576 480 8606
rect 1577 8603 1643 8606
rect 26693 8666 26759 8669
rect 29520 8666 30000 8696
rect 26693 8664 30000 8666
rect 26693 8608 26698 8664
rect 26754 8608 30000 8664
rect 26693 8606 30000 8608
rect 26693 8603 26759 8606
rect 29520 8576 30000 8606
rect 3693 8394 3759 8397
rect 6361 8394 6427 8397
rect 3693 8392 6427 8394
rect 3693 8336 3698 8392
rect 3754 8336 6366 8392
rect 6422 8336 6427 8392
rect 3693 8334 6427 8336
rect 3693 8331 3759 8334
rect 6361 8331 6427 8334
rect 15745 8394 15811 8397
rect 15929 8394 15995 8397
rect 15745 8392 15995 8394
rect 15745 8336 15750 8392
rect 15806 8336 15934 8392
rect 15990 8336 15995 8392
rect 15745 8334 15995 8336
rect 15745 8331 15811 8334
rect 15929 8331 15995 8334
rect 18873 8394 18939 8397
rect 23197 8394 23263 8397
rect 18873 8392 23263 8394
rect 18873 8336 18878 8392
rect 18934 8336 23202 8392
rect 23258 8336 23263 8392
rect 18873 8334 23263 8336
rect 18873 8331 18939 8334
rect 23197 8331 23263 8334
rect 25773 8394 25839 8397
rect 26785 8394 26851 8397
rect 25773 8392 26851 8394
rect 25773 8336 25778 8392
rect 25834 8336 26790 8392
rect 26846 8336 26851 8392
rect 25773 8334 26851 8336
rect 25773 8331 25839 8334
rect 26785 8331 26851 8334
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 2589 8122 2655 8125
rect 27429 8122 27495 8125
rect 0 8120 2655 8122
rect 0 8064 2594 8120
rect 2650 8064 2655 8120
rect 0 8062 2655 8064
rect 0 8032 480 8062
rect 2589 8059 2655 8062
rect 21406 8120 27495 8122
rect 21406 8064 27434 8120
rect 27490 8064 27495 8120
rect 21406 8062 27495 8064
rect 3509 7986 3575 7989
rect 9857 7986 9923 7989
rect 10317 7986 10383 7989
rect 12525 7986 12591 7989
rect 16297 7986 16363 7989
rect 21406 7986 21466 8062
rect 27429 8059 27495 8062
rect 27613 8122 27679 8125
rect 29520 8122 30000 8152
rect 27613 8120 30000 8122
rect 27613 8064 27618 8120
rect 27674 8064 30000 8120
rect 27613 8062 30000 8064
rect 27613 8059 27679 8062
rect 29520 8032 30000 8062
rect 3509 7984 10058 7986
rect 3509 7928 3514 7984
rect 3570 7928 9862 7984
rect 9918 7928 10058 7984
rect 3509 7926 10058 7928
rect 3509 7923 3575 7926
rect 9857 7923 9923 7926
rect 657 7850 723 7853
rect 9998 7850 10058 7926
rect 10317 7984 12591 7986
rect 10317 7928 10322 7984
rect 10378 7928 12530 7984
rect 12586 7928 12591 7984
rect 10317 7926 12591 7928
rect 10317 7923 10383 7926
rect 12525 7923 12591 7926
rect 16254 7984 21466 7986
rect 16254 7928 16302 7984
rect 16358 7928 21466 7984
rect 16254 7926 21466 7928
rect 16254 7923 16363 7926
rect 16254 7850 16314 7923
rect 657 7848 7666 7850
rect 657 7792 662 7848
rect 718 7792 7666 7848
rect 657 7790 7666 7792
rect 9998 7790 16314 7850
rect 17033 7850 17099 7853
rect 19149 7850 19215 7853
rect 26509 7850 26575 7853
rect 17033 7848 26575 7850
rect 17033 7792 17038 7848
rect 17094 7792 19154 7848
rect 19210 7792 26514 7848
rect 26570 7792 26575 7848
rect 17033 7790 26575 7792
rect 657 7787 723 7790
rect 7606 7714 7666 7790
rect 17033 7787 17099 7790
rect 19149 7787 19215 7790
rect 26509 7787 26575 7790
rect 13445 7714 13511 7717
rect 7606 7712 13511 7714
rect 7606 7656 13450 7712
rect 13506 7656 13511 7712
rect 7606 7654 13511 7656
rect 13445 7651 13511 7654
rect 16665 7714 16731 7717
rect 23105 7714 23171 7717
rect 16665 7712 23171 7714
rect 16665 7656 16670 7712
rect 16726 7656 23110 7712
rect 23166 7656 23171 7712
rect 16665 7654 23171 7656
rect 16665 7651 16731 7654
rect 23105 7651 23171 7654
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 7281 7578 7347 7581
rect 15469 7578 15535 7581
rect 7281 7576 15535 7578
rect 7281 7520 7286 7576
rect 7342 7520 15474 7576
rect 15530 7520 15535 7576
rect 7281 7518 15535 7520
rect 7281 7515 7347 7518
rect 15469 7515 15535 7518
rect 16389 7578 16455 7581
rect 23933 7578 23999 7581
rect 16389 7576 23999 7578
rect 16389 7520 16394 7576
rect 16450 7520 23938 7576
rect 23994 7520 23999 7576
rect 16389 7518 23999 7520
rect 16389 7515 16455 7518
rect 23933 7515 23999 7518
rect 0 7442 480 7472
rect 1577 7442 1643 7445
rect 0 7440 1643 7442
rect 0 7384 1582 7440
rect 1638 7384 1643 7440
rect 0 7382 1643 7384
rect 0 7352 480 7382
rect 1577 7379 1643 7382
rect 4613 7442 4679 7445
rect 15009 7442 15075 7445
rect 4613 7440 15075 7442
rect 4613 7384 4618 7440
rect 4674 7384 15014 7440
rect 15070 7384 15075 7440
rect 4613 7382 15075 7384
rect 4613 7379 4679 7382
rect 15009 7379 15075 7382
rect 25497 7442 25563 7445
rect 29520 7442 30000 7472
rect 25497 7440 30000 7442
rect 25497 7384 25502 7440
rect 25558 7384 30000 7440
rect 25497 7382 30000 7384
rect 25497 7379 25563 7382
rect 29520 7352 30000 7382
rect 2037 7306 2103 7309
rect 17309 7306 17375 7309
rect 2037 7304 17375 7306
rect 2037 7248 2042 7304
rect 2098 7248 17314 7304
rect 17370 7248 17375 7304
rect 2037 7246 17375 7248
rect 2037 7243 2103 7246
rect 17309 7243 17375 7246
rect 2129 7170 2195 7173
rect 4613 7170 4679 7173
rect 2129 7168 4679 7170
rect 2129 7112 2134 7168
rect 2190 7112 4618 7168
rect 4674 7112 4679 7168
rect 2129 7110 4679 7112
rect 2129 7107 2195 7110
rect 4613 7107 4679 7110
rect 23105 7170 23171 7173
rect 26509 7170 26575 7173
rect 23105 7168 26575 7170
rect 23105 7112 23110 7168
rect 23166 7112 26514 7168
rect 26570 7112 26575 7168
rect 23105 7110 26575 7112
rect 23105 7107 23171 7110
rect 26509 7107 26575 7110
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 0 6898 480 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 480 6838
rect 1577 6835 1643 6838
rect 2865 6898 2931 6901
rect 19241 6898 19307 6901
rect 22645 6898 22711 6901
rect 2865 6896 22711 6898
rect 2865 6840 2870 6896
rect 2926 6840 19246 6896
rect 19302 6840 22650 6896
rect 22706 6840 22711 6896
rect 2865 6838 22711 6840
rect 2865 6835 2931 6838
rect 19241 6835 19307 6838
rect 22645 6835 22711 6838
rect 26693 6898 26759 6901
rect 29520 6898 30000 6928
rect 26693 6896 30000 6898
rect 26693 6840 26698 6896
rect 26754 6840 30000 6896
rect 26693 6838 30000 6840
rect 26693 6835 26759 6838
rect 29520 6808 30000 6838
rect 1393 6762 1459 6765
rect 6821 6762 6887 6765
rect 9765 6762 9831 6765
rect 10869 6762 10935 6765
rect 13813 6762 13879 6765
rect 18873 6762 18939 6765
rect 1393 6760 6562 6762
rect 1393 6704 1398 6760
rect 1454 6704 6562 6760
rect 1393 6702 6562 6704
rect 1393 6699 1459 6702
rect 6502 6626 6562 6702
rect 6821 6760 9831 6762
rect 6821 6704 6826 6760
rect 6882 6704 9770 6760
rect 9826 6704 9831 6760
rect 6821 6702 9831 6704
rect 6821 6699 6887 6702
rect 9765 6699 9831 6702
rect 9998 6760 18939 6762
rect 9998 6704 10874 6760
rect 10930 6704 13818 6760
rect 13874 6704 18878 6760
rect 18934 6704 18939 6760
rect 9998 6702 18939 6704
rect 8661 6626 8727 6629
rect 6502 6624 8727 6626
rect 6502 6568 8666 6624
rect 8722 6568 8727 6624
rect 6502 6566 8727 6568
rect 8661 6563 8727 6566
rect 9765 6626 9831 6629
rect 9998 6626 10058 6702
rect 10869 6699 10935 6702
rect 13813 6699 13879 6702
rect 18873 6699 18939 6702
rect 9765 6624 10058 6626
rect 9765 6568 9770 6624
rect 9826 6568 10058 6624
rect 9765 6566 10058 6568
rect 9765 6563 9831 6566
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 8201 6490 8267 6493
rect 12801 6490 12867 6493
rect 8201 6488 12867 6490
rect 8201 6432 8206 6488
rect 8262 6432 12806 6488
rect 12862 6432 12867 6488
rect 8201 6430 12867 6432
rect 8201 6427 8267 6430
rect 12801 6427 12867 6430
rect 0 6354 480 6384
rect 1577 6354 1643 6357
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 480 6294
rect 1577 6291 1643 6294
rect 10501 6354 10567 6357
rect 16389 6354 16455 6357
rect 10501 6352 16455 6354
rect 10501 6296 10506 6352
rect 10562 6296 16394 6352
rect 16450 6296 16455 6352
rect 10501 6294 16455 6296
rect 10501 6291 10567 6294
rect 16389 6291 16455 6294
rect 19517 6354 19583 6357
rect 23473 6354 23539 6357
rect 19517 6352 23539 6354
rect 19517 6296 19522 6352
rect 19578 6296 23478 6352
rect 23534 6296 23539 6352
rect 19517 6294 23539 6296
rect 19517 6291 19583 6294
rect 23473 6291 23539 6294
rect 26601 6354 26667 6357
rect 29520 6354 30000 6384
rect 26601 6352 30000 6354
rect 26601 6296 26606 6352
rect 26662 6296 30000 6352
rect 26601 6294 30000 6296
rect 26601 6291 26667 6294
rect 2497 6218 2563 6221
rect 3233 6218 3299 6221
rect 11789 6218 11855 6221
rect 15561 6218 15627 6221
rect 2497 6216 15627 6218
rect 2497 6160 2502 6216
rect 2558 6160 3238 6216
rect 3294 6160 11794 6216
rect 11850 6160 15566 6216
rect 15622 6160 15627 6216
rect 2497 6158 15627 6160
rect 2497 6155 2563 6158
rect 3233 6155 3299 6158
rect 11789 6155 11855 6158
rect 15561 6155 15627 6158
rect 13353 6082 13419 6085
rect 19520 6082 19580 6291
rect 29520 6264 30000 6294
rect 23197 6218 23263 6221
rect 25681 6218 25747 6221
rect 23197 6216 25747 6218
rect 23197 6160 23202 6216
rect 23258 6160 25686 6216
rect 25742 6160 25747 6216
rect 23197 6158 25747 6160
rect 23197 6155 23263 6158
rect 25681 6155 25747 6158
rect 13353 6080 19580 6082
rect 13353 6024 13358 6080
rect 13414 6024 19580 6080
rect 13353 6022 19580 6024
rect 13353 6019 13419 6022
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 3785 5946 3851 5949
rect 8017 5946 8083 5949
rect 3785 5944 8083 5946
rect 3785 5888 3790 5944
rect 3846 5888 8022 5944
rect 8078 5888 8083 5944
rect 3785 5886 8083 5888
rect 3785 5883 3851 5886
rect 8017 5883 8083 5886
rect 24945 5810 25011 5813
rect 27429 5810 27495 5813
rect 24945 5808 27495 5810
rect 24945 5752 24950 5808
rect 25006 5752 27434 5808
rect 27490 5752 27495 5808
rect 24945 5750 27495 5752
rect 24945 5747 25011 5750
rect 27429 5747 27495 5750
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 2865 5674 2931 5677
rect 10041 5674 10107 5677
rect 2865 5672 10107 5674
rect 2865 5616 2870 5672
rect 2926 5616 10046 5672
rect 10102 5616 10107 5672
rect 2865 5614 10107 5616
rect 2865 5611 2931 5614
rect 10041 5611 10107 5614
rect 26693 5674 26759 5677
rect 29520 5674 30000 5704
rect 26693 5672 30000 5674
rect 26693 5616 26698 5672
rect 26754 5616 30000 5672
rect 26693 5614 30000 5616
rect 26693 5611 26759 5614
rect 29520 5584 30000 5614
rect 7925 5538 7991 5541
rect 12525 5538 12591 5541
rect 13169 5538 13235 5541
rect 7925 5536 13235 5538
rect 7925 5480 7930 5536
rect 7986 5480 12530 5536
rect 12586 5480 13174 5536
rect 13230 5480 13235 5536
rect 7925 5478 13235 5480
rect 7925 5475 7991 5478
rect 12525 5475 12591 5478
rect 13169 5475 13235 5478
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 8569 5402 8635 5405
rect 12157 5402 12223 5405
rect 8569 5400 12223 5402
rect 8569 5344 8574 5400
rect 8630 5344 12162 5400
rect 12218 5344 12223 5400
rect 8569 5342 12223 5344
rect 8569 5339 8635 5342
rect 12157 5339 12223 5342
rect 19057 5402 19123 5405
rect 22737 5402 22803 5405
rect 19057 5400 22803 5402
rect 19057 5344 19062 5400
rect 19118 5344 22742 5400
rect 22798 5344 22803 5400
rect 19057 5342 22803 5344
rect 19057 5339 19123 5342
rect 22737 5339 22803 5342
rect 5349 5266 5415 5269
rect 7097 5266 7163 5269
rect 5349 5264 7163 5266
rect 5349 5208 5354 5264
rect 5410 5208 7102 5264
rect 7158 5208 7163 5264
rect 5349 5206 7163 5208
rect 5349 5203 5415 5206
rect 7097 5203 7163 5206
rect 16297 5266 16363 5269
rect 18045 5266 18111 5269
rect 16297 5264 18111 5266
rect 16297 5208 16302 5264
rect 16358 5208 18050 5264
rect 18106 5208 18111 5264
rect 16297 5206 18111 5208
rect 16297 5203 16363 5206
rect 18045 5203 18111 5206
rect 24301 5266 24367 5269
rect 26509 5266 26575 5269
rect 24301 5264 26575 5266
rect 24301 5208 24306 5264
rect 24362 5208 26514 5264
rect 26570 5208 26575 5264
rect 24301 5206 26575 5208
rect 24301 5203 24367 5206
rect 26509 5203 26575 5206
rect 0 5130 480 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 480 5070
rect 1577 5067 1643 5070
rect 2037 5130 2103 5133
rect 9949 5130 10015 5133
rect 2037 5128 10015 5130
rect 2037 5072 2042 5128
rect 2098 5072 9954 5128
rect 10010 5072 10015 5128
rect 2037 5070 10015 5072
rect 2037 5067 2103 5070
rect 9949 5067 10015 5070
rect 14181 5130 14247 5133
rect 26417 5130 26483 5133
rect 14181 5128 26483 5130
rect 14181 5072 14186 5128
rect 14242 5072 26422 5128
rect 26478 5072 26483 5128
rect 14181 5070 26483 5072
rect 14181 5067 14247 5070
rect 26417 5067 26483 5070
rect 26601 5130 26667 5133
rect 29520 5130 30000 5160
rect 26601 5128 30000 5130
rect 26601 5072 26606 5128
rect 26662 5072 30000 5128
rect 26601 5070 30000 5072
rect 26601 5067 26667 5070
rect 29520 5040 30000 5070
rect 3141 4994 3207 4997
rect 7005 4994 7071 4997
rect 3141 4992 7071 4994
rect 3141 4936 3146 4992
rect 3202 4936 7010 4992
rect 7066 4936 7071 4992
rect 3141 4934 7071 4936
rect 3141 4931 3207 4934
rect 7005 4931 7071 4934
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 16481 4722 16547 4725
rect 19241 4722 19307 4725
rect 16481 4720 19307 4722
rect 16481 4664 16486 4720
rect 16542 4664 19246 4720
rect 19302 4664 19307 4720
rect 16481 4662 19307 4664
rect 16481 4659 16547 4662
rect 19241 4659 19307 4662
rect 12157 4586 12223 4589
rect 12801 4586 12867 4589
rect 24301 4586 24367 4589
rect 12157 4584 24367 4586
rect 12157 4528 12162 4584
rect 12218 4528 12806 4584
rect 12862 4528 24306 4584
rect 24362 4528 24367 4584
rect 12157 4526 24367 4528
rect 12157 4523 12223 4526
rect 12801 4523 12867 4526
rect 24301 4523 24367 4526
rect 25773 4586 25839 4589
rect 25773 4584 26434 4586
rect 25773 4528 25778 4584
rect 25834 4528 26434 4584
rect 25773 4526 26434 4528
rect 25773 4523 25839 4526
rect 0 4450 480 4480
rect 2773 4450 2839 4453
rect 0 4448 2839 4450
rect 0 4392 2778 4448
rect 2834 4392 2839 4448
rect 0 4390 2839 4392
rect 26374 4450 26434 4526
rect 29520 4450 30000 4480
rect 26374 4390 30000 4450
rect 0 4360 480 4390
rect 2773 4387 2839 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 10133 4314 10199 4317
rect 12249 4314 12315 4317
rect 10133 4312 12315 4314
rect 10133 4256 10138 4312
rect 10194 4256 12254 4312
rect 12310 4256 12315 4312
rect 10133 4254 12315 4256
rect 10133 4251 10199 4254
rect 12249 4251 12315 4254
rect 3233 4042 3299 4045
rect 8385 4042 8451 4045
rect 13445 4042 13511 4045
rect 3233 4040 13511 4042
rect 3233 3984 3238 4040
rect 3294 3984 8390 4040
rect 8446 3984 13450 4040
rect 13506 3984 13511 4040
rect 3233 3982 13511 3984
rect 3233 3979 3299 3982
rect 8385 3979 8451 3982
rect 13445 3979 13511 3982
rect 14641 4042 14707 4045
rect 17953 4042 18019 4045
rect 14641 4040 18019 4042
rect 14641 3984 14646 4040
rect 14702 3984 17958 4040
rect 18014 3984 18019 4040
rect 14641 3982 18019 3984
rect 14641 3979 14707 3982
rect 17953 3979 18019 3982
rect 19885 4042 19951 4045
rect 27521 4042 27587 4045
rect 19885 4040 27587 4042
rect 19885 3984 19890 4040
rect 19946 3984 27526 4040
rect 27582 3984 27587 4040
rect 19885 3982 27587 3984
rect 19885 3979 19951 3982
rect 27521 3979 27587 3982
rect 0 3906 480 3936
rect 2497 3906 2563 3909
rect 0 3904 2563 3906
rect 0 3848 2502 3904
rect 2558 3848 2563 3904
rect 0 3846 2563 3848
rect 0 3816 480 3846
rect 2497 3843 2563 3846
rect 15469 3906 15535 3909
rect 18873 3906 18939 3909
rect 15469 3904 18939 3906
rect 15469 3848 15474 3904
rect 15530 3848 18878 3904
rect 18934 3848 18939 3904
rect 15469 3846 18939 3848
rect 15469 3843 15535 3846
rect 18873 3843 18939 3846
rect 27705 3906 27771 3909
rect 29520 3906 30000 3936
rect 27705 3904 30000 3906
rect 27705 3848 27710 3904
rect 27766 3848 30000 3904
rect 27705 3846 30000 3848
rect 27705 3843 27771 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 2405 3634 2471 3637
rect 5625 3634 5691 3637
rect 2405 3632 5691 3634
rect 2405 3576 2410 3632
rect 2466 3576 5630 3632
rect 5686 3576 5691 3632
rect 2405 3574 5691 3576
rect 2405 3571 2471 3574
rect 5625 3571 5691 3574
rect 19609 3634 19675 3637
rect 26509 3634 26575 3637
rect 19609 3632 26575 3634
rect 19609 3576 19614 3632
rect 19670 3576 26514 3632
rect 26570 3576 26575 3632
rect 19609 3574 26575 3576
rect 19609 3571 19675 3574
rect 26509 3571 26575 3574
rect 5073 3498 5139 3501
rect 6361 3498 6427 3501
rect 26417 3498 26483 3501
rect 5073 3496 26483 3498
rect 5073 3440 5078 3496
rect 5134 3440 6366 3496
rect 6422 3440 26422 3496
rect 26478 3440 26483 3496
rect 5073 3438 26483 3440
rect 5073 3435 5139 3438
rect 6361 3435 6427 3438
rect 26417 3435 26483 3438
rect 0 3362 480 3392
rect 1393 3362 1459 3365
rect 0 3360 1459 3362
rect 0 3304 1398 3360
rect 1454 3304 1459 3360
rect 0 3302 1459 3304
rect 0 3272 480 3302
rect 1393 3299 1459 3302
rect 26693 3362 26759 3365
rect 29520 3362 30000 3392
rect 26693 3360 30000 3362
rect 26693 3304 26698 3360
rect 26754 3304 30000 3360
rect 26693 3302 30000 3304
rect 26693 3299 26759 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 18597 3090 18663 3093
rect 26233 3090 26299 3093
rect 18597 3088 26299 3090
rect 18597 3032 18602 3088
rect 18658 3032 26238 3088
rect 26294 3032 26299 3088
rect 18597 3030 26299 3032
rect 18597 3027 18663 3030
rect 26233 3027 26299 3030
rect 19425 2954 19491 2957
rect 26325 2954 26391 2957
rect 19425 2952 26391 2954
rect 19425 2896 19430 2952
rect 19486 2896 26330 2952
rect 26386 2896 26391 2952
rect 19425 2894 26391 2896
rect 19425 2891 19491 2894
rect 26325 2891 26391 2894
rect 5809 2818 5875 2821
rect 9213 2818 9279 2821
rect 5809 2816 9279 2818
rect 5809 2760 5814 2816
rect 5870 2760 9218 2816
rect 9274 2760 9279 2816
rect 5809 2758 9279 2760
rect 5809 2755 5875 2758
rect 9213 2755 9279 2758
rect 13721 2818 13787 2821
rect 16297 2818 16363 2821
rect 13721 2816 16363 2818
rect 13721 2760 13726 2816
rect 13782 2760 16302 2816
rect 16358 2760 16363 2816
rect 13721 2758 16363 2760
rect 13721 2755 13787 2758
rect 16297 2755 16363 2758
rect 26601 2818 26667 2821
rect 26601 2816 26802 2818
rect 26601 2760 26606 2816
rect 26662 2760 26802 2816
rect 26601 2758 26802 2760
rect 26601 2755 26667 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 1577 2682 1643 2685
rect 0 2680 1643 2682
rect 0 2624 1582 2680
rect 1638 2624 1643 2680
rect 0 2622 1643 2624
rect 26742 2682 26802 2758
rect 29520 2682 30000 2712
rect 26742 2622 30000 2682
rect 0 2592 480 2622
rect 1577 2619 1643 2622
rect 29520 2592 30000 2622
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 2865 2138 2931 2141
rect 0 2136 2931 2138
rect 0 2080 2870 2136
rect 2926 2080 2931 2136
rect 0 2078 2931 2080
rect 0 2048 480 2078
rect 2865 2075 2931 2078
rect 27613 2138 27679 2141
rect 29520 2138 30000 2168
rect 27613 2136 30000 2138
rect 27613 2080 27618 2136
rect 27674 2080 30000 2136
rect 27613 2078 30000 2080
rect 27613 2075 27679 2078
rect 29520 2048 30000 2078
rect 0 1458 480 1488
rect 1761 1458 1827 1461
rect 0 1456 1827 1458
rect 0 1400 1766 1456
rect 1822 1400 1827 1456
rect 0 1398 1827 1400
rect 0 1368 480 1398
rect 1761 1395 1827 1398
rect 26785 1458 26851 1461
rect 29520 1458 30000 1488
rect 26785 1456 30000 1458
rect 26785 1400 26790 1456
rect 26846 1400 30000 1456
rect 26785 1398 30000 1400
rect 26785 1395 26851 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 2957 914 3023 917
rect 0 912 3023 914
rect 0 856 2962 912
rect 3018 856 3023 912
rect 0 854 3023 856
rect 0 824 480 854
rect 2957 851 3023 854
rect 25865 914 25931 917
rect 29520 914 30000 944
rect 25865 912 30000 914
rect 25865 856 25870 912
rect 25926 856 30000 912
rect 25865 854 30000 856
rect 25865 851 25931 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 2773 370 2839 373
rect 0 368 2839 370
rect 0 312 2778 368
rect 2834 312 2839 368
rect 0 310 2839 312
rect 0 280 480 310
rect 2773 307 2839 310
rect 26509 370 26575 373
rect 29520 370 30000 400
rect 26509 368 30000 370
rect 26509 312 26514 368
rect 26570 312 30000 368
rect 26509 310 30000 312
rect 26509 307 26575 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 9628 14724 9692 14788
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 9628 14452 9692 14516
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 25084 12472 25148 12476
rect 25084 12416 25134 12472
rect 25134 12416 25148 12472
rect 25084 12412 25148 12416
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 25084 9284 25148 9348
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 9627 14788 9693 14789
rect 9627 14724 9628 14788
rect 9692 14724 9693 14788
rect 9627 14723 9693 14724
rect 9630 14517 9690 14723
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 9627 14516 9693 14517
rect 9627 14452 9628 14516
rect 9692 14452 9693 14516
rect 9627 14451 9693 14452
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25083 12476 25149 12477
rect 25083 12412 25084 12476
rect 25148 12412 25149 12476
rect 25083 12411 25149 12412
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 25086 9349 25146 12411
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25083 9348 25149 9349
rect 25083 9284 25084 9348
rect 25148 9284 25149 9348
rect 25083 9283 25149 9284
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_9 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1564 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1604681595
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20
timestamp 1604681595
transform 1 0 2944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 2668 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1472 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_28
timestamp 1604681595
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25
timestamp 1604681595
transform 1 0 3404 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3036 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1604681595
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1604681595
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3128 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38
timestamp 1604681595
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_41
timestamp 1604681595
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_49
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1604681595
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46
timestamp 1604681595
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42
timestamp 1604681595
transform 1 0 4968 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5520 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8648 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 1604681595
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_73
timestamp 1604681595
transform 1 0 7820 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_74 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_88
timestamp 1604681595
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_92
timestamp 1604681595
transform 1 0 9568 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_104
timestamp 1604681595
transform 1 0 10672 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_110
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_116
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1604681595
transform 1 0 13340 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1604681595
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13156 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1604681595
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13708 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1604681595
transform 1 0 14076 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_164
timestamp 1604681595
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15732 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_180
timestamp 1604681595
transform 1 0 17664 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 1604681595
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_168
timestamp 1604681595
transform 1 0 16560 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_190
timestamp 1604681595
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1604681595
transform 1 0 19228 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18952 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1604681595
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1604681595
transform 1 0 20148 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_217
timestamp 1604681595
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_228
timestamp 1604681595
transform 1 0 22080 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_224
timestamp 1604681595
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_221
timestamp 1604681595
transform 1 0 21436 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_233
timestamp 1604681595
transform 1 0 22540 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22632 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_241
timestamp 1604681595
transform 1 0 23276 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_261
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_251
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_255
timestamp 1604681595
transform 1 0 24564 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_267
timestamp 1604681595
transform 1 0 25668 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1604681595
transform 1 0 26680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_273
timestamp 1604681595
transform 1 0 26220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1604681595
transform 1 0 26404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 26864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 26312 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_290
timestamp 1604681595
transform 1 0 27784 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_282
timestamp 1604681595
transform 1 0 27048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 27232 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 27416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_284
timestamp 1604681595
transform 1 0 27232 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 27968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp 1604681595
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_294
timestamp 1604681595
transform 1 0 28152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_298
timestamp 1604681595
transform 1 0 28520 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 2300 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5612 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_55
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_67
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_77
timestamp 1604681595
transform 1 0 8188 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1604681595
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16008 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1604681595
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1604681595
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_186
timestamp 1604681595
transform 1 0 18216 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18492 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_205
timestamp 1604681595
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1604681595
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_280
timestamp 1604681595
transform 1 0 26864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 1604681595
transform 1 0 27968 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1604681595
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1472 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1604681595
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4600 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1604681595
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_30
timestamp 1604681595
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_34
timestamp 1604681595
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1604681595
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_66
timestamp 1604681595
transform 1 0 7176 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_84
timestamp 1604681595
transform 1 0 8832 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_92
timestamp 1604681595
transform 1 0 9568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_95
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_99
timestamp 1604681595
transform 1 0 10212 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_111
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1604681595
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1604681595
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1604681595
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_143
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 14536 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1604681595
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1604681595
transform 1 0 17480 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1604681595
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18492 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_188
timestamp 1604681595
transform 1 0 18400 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_191
timestamp 1604681595
transform 1 0 18676 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1604681595
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_212
timestamp 1604681595
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_216
timestamp 1604681595
transform 1 0 20976 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_228
timestamp 1604681595
transform 1 0 22080 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_240
timestamp 1604681595
transform 1 0 23184 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 27508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 26404 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 27324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_279
timestamp 1604681595
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_283
timestamp 1604681595
transform 1 0 27140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_291
timestamp 1604681595
transform 1 0 27876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_295
timestamp 1604681595
transform 1 0 28244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 2760 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_16
timestamp 1604681595
transform 1 0 2576 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1604681595
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_26
timestamp 1604681595
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1604681595
transform 1 0 4876 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_53
timestamp 1604681595
transform 1 0 5980 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_61
timestamp 1604681595
transform 1 0 6716 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_78
timestamp 1604681595
transform 1 0 8280 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1604681595
transform 1 0 11132 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1604681595
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_134
timestamp 1604681595
transform 1 0 13432 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_146
timestamp 1604681595
transform 1 0 14536 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1604681595
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_163
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_175
timestamp 1604681595
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_187
timestamp 1604681595
transform 1 0 18308 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_194
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 21344 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1604681595
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_222
timestamp 1604681595
transform 1 0 21528 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_234
timestamp 1604681595
transform 1 0 22632 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_246
timestamp 1604681595
transform 1 0 23736 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_258
timestamp 1604681595
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_270
timestamp 1604681595
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1604681595
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1604681595
transform 1 0 26864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_292
timestamp 1604681595
transform 1 0 27968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1604681595
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1604681595
transform 1 0 2576 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_20
timestamp 1604681595
transform 1 0 2944 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3956 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1604681595
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5704 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_48
timestamp 1604681595
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_52
timestamp 1604681595
transform 1 0 5888 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1604681595
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7544 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1604681595
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_79
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_83
timestamp 1604681595
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_87
timestamp 1604681595
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_91
timestamp 1604681595
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_103
timestamp 1604681595
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_115
timestamp 1604681595
transform 1 0 11684 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1604681595
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_143
timestamp 1604681595
transform 1 0 14260 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _18_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 15916 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_149
timestamp 1604681595
transform 1 0 14812 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_160
timestamp 1604681595
transform 1 0 15824 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_164
timestamp 1604681595
transform 1 0 16192 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_176
timestamp 1604681595
transform 1 0 17296 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_180
timestamp 1604681595
transform 1 0 17664 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_190
timestamp 1604681595
transform 1 0 18584 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_202
timestamp 1604681595
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_206
timestamp 1604681595
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1604681595
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_214
timestamp 1604681595
transform 1 0 20792 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604681595
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_279
timestamp 1604681595
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_283
timestamp 1604681595
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_287
timestamp 1604681595
transform 1 0 27508 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1604681595
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1604681595
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1604681595
transform 1 0 4876 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 3956 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_7_47
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_56
timestamp 1604681595
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_52
timestamp 1604681595
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_53
timestamp 1604681595
transform 1 0 5980 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1604681595
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_60
timestamp 1604681595
transform 1 0 6624 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_57
timestamp 1604681595
transform 1 0 6348 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7728 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1604681595
transform 1 0 7176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_81
timestamp 1604681595
transform 1 0 8556 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_73
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_81
timestamp 1604681595
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_93
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_89
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 1604681595
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1604681595
transform 1 0 9292 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10028 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 10212 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_102
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1604681595
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_106
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_114
timestamp 1604681595
transform 1 0 11592 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_116
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_120
timestamp 1604681595
transform 1 0 12144 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_132
timestamp 1604681595
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12880 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1604681595
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_141
timestamp 1604681595
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_137
timestamp 1604681595
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_136
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1604681595
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1604681595
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_148
timestamp 1604681595
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_163
timestamp 1604681595
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_176
timestamp 1604681595
transform 1 0 17296 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_172
timestamp 1604681595
transform 1 0 16928 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_168
timestamp 1604681595
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_175
timestamp 1604681595
transform 1 0 17204 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_186
timestamp 1604681595
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_183
timestamp 1604681595
transform 1 0 17940 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18400 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_205
timestamp 1604681595
transform 1 0 19964 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1604681595
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1604681595
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_217
timestamp 1604681595
transform 1 0 21068 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_229
timestamp 1604681595
transform 1 0 22172 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1604681595
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 22724 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_254
timestamp 1604681595
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_258
timestamp 1604681595
transform 1 0 24840 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_270
timestamp 1604681595
transform 1 0 25944 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_279
timestamp 1604681595
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_274
timestamp 1604681595
transform 1 0 26312 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_283
timestamp 1604681595
transform 1 0 27140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 27324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_287
timestamp 1604681595
transform 1 0 27508 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1604681595
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_292
timestamp 1604681595
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1604681595
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1604681595
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_71
timestamp 1604681595
transform 1 0 7636 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_83
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_119
timestamp 1604681595
transform 1 0 12052 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_123
timestamp 1604681595
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_126
timestamp 1604681595
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_130
timestamp 1604681595
transform 1 0 13064 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_142
timestamp 1604681595
transform 1 0 14168 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1604681595
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1604681595
transform 1 0 16744 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_174
timestamp 1604681595
transform 1 0 17112 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_177
timestamp 1604681595
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_184
timestamp 1604681595
transform 1 0 18032 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18768 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1604681595
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_205
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_229
timestamp 1604681595
transform 1 0 22172 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23000 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24012 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_233
timestamp 1604681595
transform 1 0 22540 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_237
timestamp 1604681595
transform 1 0 22908 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_247
timestamp 1604681595
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_259
timestamp 1604681595
transform 1 0 24932 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_264
timestamp 1604681595
transform 1 0 25392 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_272
timestamp 1604681595
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604681595
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604681595
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604681595
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1604681595
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1604681595
transform 1 0 5060 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_78
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_102
timestamp 1604681595
transform 1 0 10488 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1604681595
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15640 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_151
timestamp 1604681595
transform 1 0 14996 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_154
timestamp 1604681595
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_167
timestamp 1604681595
transform 1 0 16468 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_173
timestamp 1604681595
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_177
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18676 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_188
timestamp 1604681595
transform 1 0 18400 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1604681595
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_204
timestamp 1604681595
transform 1 0 19872 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_216
timestamp 1604681595
transform 1 0 20976 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604681595
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 25208 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_254
timestamp 1604681595
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_258
timestamp 1604681595
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 27416 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 26864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1604681595
transform 1 0 26680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_282
timestamp 1604681595
transform 1 0 27048 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_290
timestamp 1604681595
transform 1 0 27784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 27968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_294
timestamp 1604681595
transform 1 0 28152 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_298
timestamp 1604681595
transform 1 0 28520 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1604681595
transform 1 0 5980 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_61
timestamp 1604681595
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6900 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_70
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_82
timestamp 1604681595
transform 1 0 8648 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_101
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1604681595
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_125
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_130
timestamp 1604681595
transform 1 0 13064 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_142
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1604681595
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_160
timestamp 1604681595
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_164
timestamp 1604681595
transform 1 0 16192 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17204 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 16928 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19320 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_188
timestamp 1604681595
transform 1 0 18400 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_196
timestamp 1604681595
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_200
timestamp 1604681595
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1604681595
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1604681595
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_221
timestamp 1604681595
transform 1 0 21436 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_224
timestamp 1604681595
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_228
timestamp 1604681595
transform 1 0 22080 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 22356 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_240
timestamp 1604681595
transform 1 0 23184 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_244
timestamp 1604681595
transform 1 0 23552 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_247
timestamp 1604681595
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 24840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 1604681595
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_260
timestamp 1604681595
transform 1 0 25024 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_267
timestamp 1604681595
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1604681595
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604681595
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604681595
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604681595
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_17
timestamp 1604681595
transform 1 0 2668 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_36
timestamp 1604681595
transform 1 0 4416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_48
timestamp 1604681595
transform 1 0 5520 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_54
timestamp 1604681595
transform 1 0 6072 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_78
timestamp 1604681595
transform 1 0 8280 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 9844 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_90
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_127
timestamp 1604681595
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_130
timestamp 1604681595
transform 1 0 13064 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_134
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_137
timestamp 1604681595
transform 1 0 13708 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_145
timestamp 1604681595
transform 1 0 14444 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 15640 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1604681595
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1604681595
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_174
timestamp 1604681595
transform 1 0 17112 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp 1604681595
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18952 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_190
timestamp 1604681595
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1604681595
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_207
timestamp 1604681595
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21896 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_214
timestamp 1604681595
transform 1 0 20792 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_224
timestamp 1604681595
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23276 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_235
timestamp 1604681595
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_239
timestamp 1604681595
transform 1 0 23092 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1604681595
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1604681595
transform 1 0 25392 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_253
timestamp 1604681595
transform 1 0 24380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_256
timestamp 1604681595
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_260
timestamp 1604681595
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 26956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 27508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_273
timestamp 1604681595
transform 1 0 26220 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_278
timestamp 1604681595
transform 1 0 26680 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_285
timestamp 1604681595
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_289
timestamp 1604681595
transform 1 0 27692 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_297
timestamp 1604681595
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_35
timestamp 1604681595
transform 1 0 4324 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_47
timestamp 1604681595
transform 1 0 5428 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_61
timestamp 1604681595
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_65
timestamp 1604681595
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_69
timestamp 1604681595
transform 1 0 7452 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_81
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1604681595
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_98
timestamp 1604681595
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_102
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_110
timestamp 1604681595
transform 1 0 11224 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1604681595
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_124
timestamp 1604681595
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12880 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1604681595
transform 1 0 13708 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_142
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15916 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 15640 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_146
timestamp 1604681595
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_160
timestamp 1604681595
transform 1 0 15824 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_170
timestamp 1604681595
transform 1 0 16744 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_187
timestamp 1604681595
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19044 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_191
timestamp 1604681595
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_204
timestamp 1604681595
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21528 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1604681595
transform 1 0 21436 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 23828 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_231
timestamp 1604681595
transform 1 0 22356 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_243
timestamp 1604681595
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_250
timestamp 1604681595
transform 1 0 24104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1604681595
transform 1 0 24840 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_255
timestamp 1604681595
transform 1 0 24564 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_267
timestamp 1604681595
transform 1 0 25668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1604681595
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_280
timestamp 1604681595
transform 1 0 26864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_292
timestamp 1604681595
transform 1 0 27968 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1604681595
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_7
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1604681595
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1604681595
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 1604681595
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2760 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_31
timestamp 1604681595
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_38
timestamp 1604681595
transform 1 0 4600 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_38
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 4324 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1604681595
transform 1 0 5796 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_52
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1604681595
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_44
timestamp 1604681595
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4968 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1604681595
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_13_78
timestamp 1604681595
transform 1 0 8280 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9292 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9936 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_88
timestamp 1604681595
transform 1 0 9200 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604681595
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1604681595
transform 1 0 11132 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_109
timestamp 1604681595
transform 1 0 11132 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_122
timestamp 1604681595
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_115
timestamp 1604681595
transform 1 0 11684 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12696 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_132
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_137
timestamp 1604681595
transform 1 0 13708 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1604681595
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604681595
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1604681595
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_153
timestamp 1604681595
transform 1 0 15180 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_163
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1604681595
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_164
timestamp 1604681595
transform 1 0 16192 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1604681595
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_184
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_180
timestamp 1604681595
transform 1 0 17664 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18216 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_172
timestamp 1604681595
transform 1 0 16928 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_195
timestamp 1604681595
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1604681595
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 18768 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19044 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1604681595
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_199
timestamp 1604681595
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 21620 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1604681595
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_229
timestamp 1604681595
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1604681595
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_241
timestamp 1604681595
transform 1 0 23276 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_247
timestamp 1604681595
transform 1 0 23828 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24380 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_261
timestamp 1604681595
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_265
timestamp 1604681595
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_262
timestamp 1604681595
transform 1 0 25208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_266
timestamp 1604681595
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1604681595
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_279
timestamp 1604681595
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 26404 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_283
timestamp 1604681595
transform 1 0 27140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 27324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_280
timestamp 1604681595
transform 1 0 26864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_287
timestamp 1604681595
transform 1 0 27508 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_292
timestamp 1604681595
transform 1 0 27968 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1604681595
transform 1 0 28520 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_10
timestamp 1604681595
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 3956 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1604681595
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_35
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_39
timestamp 1604681595
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1604681595
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_133
timestamp 1604681595
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_156
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_160
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_164
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_192
timestamp 1604681595
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_228
timestamp 1604681595
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_254
timestamp 1604681595
transform 1 0 24472 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_260
timestamp 1604681595
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_264
timestamp 1604681595
transform 1 0 25392 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_268
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 26220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_271
timestamp 1604681595
transform 1 0 26036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_279
timestamp 1604681595
transform 1 0 26772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_283
timestamp 1604681595
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_287
timestamp 1604681595
transform 1 0 27508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4692 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1604681595
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1604681595
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_52
timestamp 1604681595
transform 1 0 5888 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 8280 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_64
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1604681595
transform 1 0 7728 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_75
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_81
timestamp 1604681595
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10120 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1604681595
transform 1 0 8924 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1604681595
transform 1 0 9292 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_97
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_107
timestamp 1604681595
transform 1 0 10948 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_119
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_143
timestamp 1604681595
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 16008 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_182
timestamp 1604681595
transform 1 0 17848 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 21896 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_223
timestamp 1604681595
transform 1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_242
timestamp 1604681595
transform 1 0 23368 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_246
timestamp 1604681595
transform 1 0 23736 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_249
timestamp 1604681595
transform 1 0 24012 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24840 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_255
timestamp 1604681595
transform 1 0 24564 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_267
timestamp 1604681595
transform 1 0 25668 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1604681595
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_285
timestamp 1604681595
transform 1 0 27324 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1604681595
transform 1 0 28428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_11
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1604681595
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_20
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 3404 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_41
timestamp 1604681595
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_45
timestamp 1604681595
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_49
timestamp 1604681595
transform 1 0 5612 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_66
timestamp 1604681595
transform 1 0 7176 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1604681595
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_103
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604681595
transform 1 0 10948 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12788 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_143
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_155
timestamp 1604681595
transform 1 0 15364 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1604681595
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_187
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19412 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_191
timestamp 1604681595
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_195
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1604681595
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1604681595
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23828 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_241
timestamp 1604681595
transform 1 0 23276 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1604681595
transform 1 0 25760 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_256
timestamp 1604681595
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_260
timestamp 1604681595
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1604681595
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_277
timestamp 1604681595
transform 1 0 26588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_289
timestamp 1604681595
transform 1 0 27692 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1604681595
transform 1 0 28428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_19
timestamp 1604681595
transform 1 0 2852 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_40
timestamp 1604681595
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4968 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_58
timestamp 1604681595
transform 1 0 6440 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_70
timestamp 1604681595
transform 1 0 7544 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_114
timestamp 1604681595
transform 1 0 11592 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_126
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_129
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_137
timestamp 1604681595
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1604681595
transform 1 0 15548 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16008 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_160
timestamp 1604681595
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_164
timestamp 1604681595
transform 1 0 16192 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1604681595
transform 1 0 17112 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_168
timestamp 1604681595
transform 1 0 16560 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_183
timestamp 1604681595
transform 1 0 17940 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 19044 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19504 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_191
timestamp 1604681595
transform 1 0 18676 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_194
timestamp 1604681595
transform 1 0 18952 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1604681595
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 21620 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_239
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_249
timestamp 1604681595
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24380 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25392 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_262
timestamp 1604681595
transform 1 0 25208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_266
timestamp 1604681595
transform 1 0 25576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_270
timestamp 1604681595
transform 1 0 25944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1604681595
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_279
timestamp 1604681595
transform 1 0 26772 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_291
timestamp 1604681595
transform 1 0 27876 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1604681595
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_20_25
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1604681595
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_38
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_34
timestamp 1604681595
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_31
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_40
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5244 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_54
timestamp 1604681595
transform 1 0 6072 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_55
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 8096 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8188 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1604681595
transform 1 0 7176 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_72
timestamp 1604681595
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1604681595
transform 1 0 7084 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1604681595
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_87
timestamp 1604681595
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1604681595
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1604681595
transform 1 0 10028 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_96
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_109
timestamp 1604681595
transform 1 0 11132 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_108
timestamp 1604681595
transform 1 0 11040 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_117
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 11960 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13892 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_127
timestamp 1604681595
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_138
timestamp 1604681595
transform 1 0 13800 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1604681595
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1604681595
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_165
timestamp 1604681595
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15456 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1604681595
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1604681595
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_186
timestamp 1604681595
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_180
timestamp 1604681595
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_189
timestamp 1604681595
transform 1 0 18492 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp 1604681595
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18768 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_205
timestamp 1604681595
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_201
timestamp 1604681595
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1604681595
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_222
timestamp 1604681595
transform 1 0 21528 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1604681595
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_226
timestamp 1604681595
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1604681595
transform 1 0 21436 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 21344 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_209
timestamp 1604681595
transform 1 0 20332 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21712 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24012 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_230
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_240
timestamp 1604681595
transform 1 0 23184 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_248
timestamp 1604681595
transform 1 0 23920 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1604681595
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1604681595
transform 1 0 24380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_260
timestamp 1604681595
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24196 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 1604681595
transform 1 0 25392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25208 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 25760 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_284
timestamp 1604681595
transform 1 0 27232 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1604681595
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_288
timestamp 1604681595
transform 1 0 27600 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_296
timestamp 1604681595
transform 1 0 28336 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 1604681595
transform 1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1604681595
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_28
timestamp 1604681595
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_32
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_36
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1604681595
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8924 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_105
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1604681595
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1604681595
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1604681595
transform 1 0 14260 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_147
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp 1604681595
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_163
timestamp 1604681595
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_167
timestamp 1604681595
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18952 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_189
timestamp 1604681595
transform 1 0 18492 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_193
timestamp 1604681595
transform 1 0 18860 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_212
timestamp 1604681595
transform 1 0 20608 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_223
timestamp 1604681595
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_227
timestamp 1604681595
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 24104 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_231
timestamp 1604681595
transform 1 0 22356 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_243
timestamp 1604681595
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_249
timestamp 1604681595
transform 1 0 24012 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 24288 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_268
timestamp 1604681595
transform 1 0 25760 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 26496 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 27048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_280
timestamp 1604681595
transform 1 0 26864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_284
timestamp 1604681595
transform 1 0 27232 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_296
timestamp 1604681595
transform 1 0 28336 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_7
timestamp 1604681595
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1604681595
transform 1 0 2116 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_36
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5428 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_42
timestamp 1604681595
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_46
timestamp 1604681595
transform 1 0 5336 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1604681595
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_64
timestamp 1604681595
transform 1 0 6992 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_76
timestamp 1604681595
transform 1 0 8096 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1604681595
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_102
timestamp 1604681595
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_107
timestamp 1604681595
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1604681595
transform 1 0 12052 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1604681595
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_142
timestamp 1604681595
transform 1 0 14168 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16284 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_150
timestamp 1604681595
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_158
timestamp 1604681595
transform 1 0 15640 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_164
timestamp 1604681595
transform 1 0 16192 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 18032 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_174
timestamp 1604681595
transform 1 0 17112 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_182
timestamp 1604681595
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_196
timestamp 1604681595
transform 1 0 19136 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_200
timestamp 1604681595
transform 1 0 19504 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21620 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_232
timestamp 1604681595
transform 1 0 22448 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1604681595
transform 1 0 23552 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 24288 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_254
timestamp 1604681595
transform 1 0 24472 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_266
timestamp 1604681595
transform 1 0 25576 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 26680 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1604681595
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_280
timestamp 1604681595
transform 1 0 26864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_292
timestamp 1604681595
transform 1 0 27968 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_298
timestamp 1604681595
transform 1 0 28520 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_19
timestamp 1604681595
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1604681595
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_36
timestamp 1604681595
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_40
timestamp 1604681595
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_75
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_87
timestamp 1604681595
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_91
timestamp 1604681595
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_95
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13708 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_129
timestamp 1604681595
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_133
timestamp 1604681595
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_146
timestamp 1604681595
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_150
timestamp 1604681595
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_166
timestamp 1604681595
transform 1 0 16376 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_197
timestamp 1604681595
transform 1 0 19228 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21620 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1604681595
transform 1 0 20332 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_215
timestamp 1604681595
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_219
timestamp 1604681595
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_253
timestamp 1604681595
transform 1 0 24380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_256
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_260
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_264
timestamp 1604681595
transform 1 0 25392 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 26864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 27232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1604681595
transform 1 0 26680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_282
timestamp 1604681595
transform 1 0 27048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_286
timestamp 1604681595
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_298
timestamp 1604681595
transform 1 0 28520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1604681595
transform 1 0 2116 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6164 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_46
timestamp 1604681595
transform 1 0 5336 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_54
timestamp 1604681595
transform 1 0 6072 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_71
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_83
timestamp 1604681595
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1604681595
transform 1 0 11132 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1604681595
transform 1 0 12236 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_142
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 16192 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1604681595
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1604681595
transform 1 0 15640 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_162
timestamp 1604681595
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17112 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_196
timestamp 1604681595
transform 1 0 19136 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_199
timestamp 1604681595
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1604681595
transform 1 0 21712 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21160 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21528 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 1604681595
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_220
timestamp 1604681595
transform 1 0 21344 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_233
timestamp 1604681595
transform 1 0 22540 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_241
timestamp 1604681595
transform 1 0 23276 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_245
timestamp 1604681595
transform 1 0 23644 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_255
timestamp 1604681595
transform 1 0 24564 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_267
timestamp 1604681595
transform 1 0 25668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1604681595
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_285
timestamp 1604681595
transform 1 0 27324 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1604681595
transform 1 0 28428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_26
timestamp 1604681595
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_30
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_34
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_46
timestamp 1604681595
transform 1 0 5336 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_49
timestamp 1604681595
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1604681595
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 1604681595
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9476 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_85
timestamp 1604681595
transform 1 0 8924 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1604681595
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1604681595
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_108
timestamp 1604681595
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1604681595
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_128
timestamp 1604681595
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_141
timestamp 1604681595
transform 1 0 14076 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_149
timestamp 1604681595
transform 1 0 14812 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_152
timestamp 1604681595
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_156
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_192
timestamp 1604681595
transform 1 0 18768 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_213
timestamp 1604681595
transform 1 0 20700 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_217
timestamp 1604681595
transform 1 0 21068 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_238
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_234
timestamp 1604681595
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_230
timestamp 1604681595
transform 1 0 22264 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 25576 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_262
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 26588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1604681595
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_279
timestamp 1604681595
transform 1 0 26772 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_291
timestamp 1604681595
transform 1 0 27876 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1604681595
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_8
timestamp 1604681595
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_19
timestamp 1604681595
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_12
timestamp 1604681595
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2024 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1604681595
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_37
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_31
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_40
timestamp 1604681595
transform 1 0 4784 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4876 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5428 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_43
timestamp 1604681595
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_50
timestamp 1604681595
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_54
timestamp 1604681595
transform 1 0 6072 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1604681595
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8188 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_63
timestamp 1604681595
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_66
timestamp 1604681595
transform 1 0 7176 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1604681595
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_90
timestamp 1604681595
transform 1 0 9384 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_102
timestamp 1604681595
transform 1 0 10488 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_105
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_119
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_131
timestamp 1604681595
transform 1 0 13156 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_134
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1604681595
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_152
timestamp 1604681595
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_156
timestamp 1604681595
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_163
timestamp 1604681595
transform 1 0 16100 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 18216 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_175
timestamp 1604681595
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_187
timestamp 1604681595
transform 1 0 18308 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_175
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18400 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1604681595
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_201
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_206
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_194
timestamp 1604681595
transform 1 0 18952 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1604681595
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21160 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_228
timestamp 1604681595
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_224
timestamp 1604681595
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22172 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_236
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_249
timestamp 1604681595
transform 1 0 24012 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 24104 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_231
timestamp 1604681595
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 23460 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_256
timestamp 1604681595
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_252
timestamp 1604681595
transform 1 0 24288 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_259
timestamp 1604681595
transform 1 0 24932 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1604681595
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_260
timestamp 1604681595
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_267
timestamp 1604681595
transform 1 0 25668 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25208 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1604681595
transform 1 0 25760 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_270
timestamp 1604681595
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1604681595
transform 1 0 26956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_277
timestamp 1604681595
transform 1 0 26588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_279
timestamp 1604681595
transform 1 0 26772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1604681595
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 26956 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 26772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 27140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_285
timestamp 1604681595
transform 1 0 27324 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_283
timestamp 1604681595
transform 1 0 27140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_295
timestamp 1604681595
transform 1 0 28244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1604681595
transform 1 0 28428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1656 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 4600 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_22
timestamp 1604681595
transform 1 0 3128 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604681595
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_54
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_62
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 6992 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_67
timestamp 1604681595
transform 1 0 7268 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_98
timestamp 1604681595
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11592 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_130
timestamp 1604681595
transform 1 0 13064 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_142
timestamp 1604681595
transform 1 0 14168 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604681595
transform 1 0 17572 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_170
timestamp 1604681595
transform 1 0 16744 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_182
timestamp 1604681595
transform 1 0 17848 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_199
timestamp 1604681595
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1604681595
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_224
timestamp 1604681595
transform 1 0 21712 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_229
timestamp 1604681595
transform 1 0 22172 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_241
timestamp 1604681595
transform 1 0 23276 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24840 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1604681595
transform 1 0 24380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_257
timestamp 1604681595
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_267
timestamp 1604681595
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_285
timestamp 1604681595
transform 1 0 27324 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1604681595
transform 1 0 28428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2024 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_19
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1604681595
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_30
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_54
timestamp 1604681595
transform 1 0 6072 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1604681595
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8096 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_92
timestamp 1604681595
transform 1 0 9568 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_97
timestamp 1604681595
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_101
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12604 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1604681595
transform 1 0 11500 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1604681595
transform 1 0 12052 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_141
timestamp 1604681595
transform 1 0 14076 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1604681595
transform 1 0 14996 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_160
timestamp 1604681595
transform 1 0 15824 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_172
timestamp 1604681595
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_180
timestamp 1604681595
transform 1 0 17664 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18584 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1604681595
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1604681595
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_207
timestamp 1604681595
transform 1 0 20148 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 21068 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_211
timestamp 1604681595
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_233
timestamp 1604681595
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_237
timestamp 1604681595
transform 1 0 22908 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1604681595
transform 1 0 23460 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 25208 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 24196 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_253
timestamp 1604681595
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_278
timestamp 1604681595
transform 1 0 26680 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_290
timestamp 1604681595
transform 1 0 27784 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp 1604681595
transform 1 0 28520 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_18
timestamp 1604681595
transform 1 0 2760 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1604681595
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8096 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_78
timestamp 1604681595
transform 1 0 8280 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 9844 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_111
timestamp 1604681595
transform 1 0 11316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_123
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_127
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_139
timestamp 1604681595
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 21068 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_219
timestamp 1604681595
transform 1 0 21252 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_243
timestamp 1604681595
transform 1 0 23460 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_267
timestamp 1604681595
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1604681595
transform 1 0 27600 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1604681595
transform 1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1604681595
transform 1 0 26956 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1604681595
transform 1 0 28060 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1604681595
transform 1 0 27600 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_296
timestamp 1604681595
transform 1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_216
timestamp 1604681595
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_234
timestamp 1604681595
transform 1 0 22632 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_242
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604681595
transform 1 0 25760 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_265
timestamp 1604681595
transform 1 0 25484 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604681595
transform 1 0 26312 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_272
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_288
timestamp 1604681595
transform 1 0 27600 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604681595
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_296
timestamp 1604681595
transform 1 0 28336 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604681595
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604681595
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604681595
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604681595
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604681595
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604681595
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 27710 0 27766 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 7470 23520 7526 24000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 29182 0 29238 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 22466 23520 22522 24000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 bottom_grid_pin_0_
port 4 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 bottom_grid_pin_10_
port 5 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 bottom_grid_pin_11_
port 6 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 bottom_grid_pin_12_
port 7 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 bottom_grid_pin_13_
port 8 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 bottom_grid_pin_14_
port 9 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 bottom_grid_pin_15_
port 10 nsew default tristate
rlabel metal2 s 6366 0 6422 480 6 bottom_grid_pin_1_
port 11 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 bottom_grid_pin_2_
port 12 nsew default tristate
rlabel metal2 s 9218 0 9274 480 6 bottom_grid_pin_3_
port 13 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 bottom_grid_pin_4_
port 14 nsew default tristate
rlabel metal2 s 12070 0 12126 480 6 bottom_grid_pin_5_
port 15 nsew default tristate
rlabel metal2 s 13450 0 13506 480 6 bottom_grid_pin_6_
port 16 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 bottom_grid_pin_7_
port 17 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 bottom_grid_pin_8_
port 18 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 bottom_grid_pin_9_
port 19 nsew default tristate
rlabel metal2 s 2042 0 2098 480 6 ccff_head
port 20 nsew default input
rlabel metal2 s 3514 0 3570 480 6 ccff_tail
port 21 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 22 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 23 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 24 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 25 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 26 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 27 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 28 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 29 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 30 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 31 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 32 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 33 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 34 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 35 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 36 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 37 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 38 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 39 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 40 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 41 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 42 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 43 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 44 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 45 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 46 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 47 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 48 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 49 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 50 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 51 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 52 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 53 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 54 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 55 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 56 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 57 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 58 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 59 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 60 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 61 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 62 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 63 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 64 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 65 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 66 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 67 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 68 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 69 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 70 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 71 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 72 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 73 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 74 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 75 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 76 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 77 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 78 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 79 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 80 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 81 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 82 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 83 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 84 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 85 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 86 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 87 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 88 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 89 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 90 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 91 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 92 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 93 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 94 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 95 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 96 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 97 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 98 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 99 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 100 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 101 nsew default tristate
rlabel metal2 s 662 0 718 480 6 prog_clk
port 102 nsew default input
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 103 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 104 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
